module h_adder (a,b,s);
parameter NBIT = 8;
input [NBIT-1:0] a,b;
output reg [NBIT:0] s;
//assign s = a + b;
always @(*)
begin
    casex({a,b})
	{8'd0,8'd0} : s = 0;
	{8'd0,8'd1} : s = 256;
	{8'd0,8'd2} : s = 128;
	{8'd0,8'd3} : s = 384;
	{8'd0,8'd4} : s = 64;
	{8'd0,8'd5} : s = 320;
	{8'd0,8'd6} : s = 288;
	{8'd0,8'd7} : s = 448;
	{8'd0,8'd8} : s = 32;
	{8'd0,8'd9} : s = 272;
	{8'd0,8'd10} : s = 264;
	{8'd0,8'd11} : s = 416;
	{8'd0,8'd12} : s = 260;
	{8'd0,8'd13} : s = 400;
	{8'd0,8'd14} : s = 392;
	{8'd0,8'd15} : s = 480;
	{8'd0,8'd16} : s = 8;
	{8'd0,8'd17} : s = 258;
	{8'd0,8'd18} : s = 257;
	{8'd0,8'd19} : s = 388;
	{8'd0,8'd20} : s = 192;
	{8'd0,8'd21} : s = 386;
	{8'd0,8'd22} : s = 385;
	{8'd0,8'd23} : s = 464;
	{8'd0,8'd24} : s = 160;
	{8'd0,8'd25} : s = 352;
	{8'd0,8'd26} : s = 336;
	{8'd0,8'd27} : s = 456;
	{8'd0,8'd28} : s = 328;
	{8'd0,8'd29} : s = 452;
	{8'd0,8'd30} : s = 450;
	{8'd0,8'd31} : s = 496;
	{8'd0,8'd32} : s = 16;
	{8'd0,8'd33} : s = 144;
	{8'd0,8'd34} : s = 136;
	{8'd0,8'd35} : s = 324;
	{8'd0,8'd36} : s = 132;
	{8'd0,8'd37} : s = 322;
	{8'd0,8'd38} : s = 321;
	{8'd0,8'd39} : s = 449;
	{8'd0,8'd40} : s = 130;
	{8'd0,8'd41} : s = 304;
	{8'd0,8'd42} : s = 296;
	{8'd0,8'd43} : s = 432;
	{8'd0,8'd44} : s = 292;
	{8'd0,8'd45} : s = 424;
	{8'd0,8'd46} : s = 420;
	{8'd0,8'd47} : s = 488;
	{8'd0,8'd48} : s = 129;
	{8'd0,8'd49} : s = 290;
	{8'd0,8'd50} : s = 289;
	{8'd0,8'd51} : s = 418;
	{8'd0,8'd52} : s = 280;
	{8'd0,8'd53} : s = 417;
	{8'd0,8'd54} : s = 408;
	{8'd0,8'd55} : s = 484;
	{8'd0,8'd56} : s = 276;
	{8'd0,8'd57} : s = 404;
	{8'd0,8'd58} : s = 402;
	{8'd0,8'd59} : s = 482;
	{8'd0,8'd60} : s = 401;
	{8'd0,8'd61} : s = 481;
	{8'd0,8'd62} : s = 472;
	{8'd0,8'd63} : s = 504;
	{8'd0,8'd64} : s = 4;
	{8'd0,8'd65} : s = 96;
	{8'd0,8'd66} : s = 80;
	{8'd0,8'd67} : s = 274;
	{8'd0,8'd68} : s = 72;
	{8'd0,8'd69} : s = 273;
	{8'd0,8'd70} : s = 268;
	{8'd0,8'd71} : s = 396;
	{8'd0,8'd72} : s = 68;
	{8'd0,8'd73} : s = 266;
	{8'd0,8'd74} : s = 265;
	{8'd0,8'd75} : s = 394;
	{8'd0,8'd76} : s = 262;
	{8'd0,8'd77} : s = 393;
	{8'd0,8'd78} : s = 390;
	{8'd0,8'd79} : s = 468;
	{8'd0,8'd80} : s = 66;
	{8'd0,8'd81} : s = 261;
	{8'd0,8'd82} : s = 259;
	{8'd0,8'd83} : s = 389;
	{8'd0,8'd84} : s = 224;
	{8'd0,8'd85} : s = 387;
	{8'd0,8'd86} : s = 368;
	{8'd0,8'd87} : s = 466;
	{8'd0,8'd88} : s = 208;
	{8'd0,8'd89} : s = 360;
	{8'd0,8'd90} : s = 356;
	{8'd0,8'd91} : s = 465;
	{8'd0,8'd92} : s = 354;
	{8'd0,8'd93} : s = 460;
	{8'd0,8'd94} : s = 458;
	{8'd0,8'd95} : s = 500;
	{8'd0,8'd96} : s = 65;
	{8'd0,8'd97} : s = 200;
	{8'd0,8'd98} : s = 196;
	{8'd0,8'd99} : s = 353;
	{8'd0,8'd100} : s = 194;
	{8'd0,8'd101} : s = 344;
	{8'd0,8'd102} : s = 340;
	{8'd0,8'd103} : s = 457;
	{8'd0,8'd104} : s = 193;
	{8'd0,8'd105} : s = 338;
	{8'd0,8'd106} : s = 337;
	{8'd0,8'd107} : s = 454;
	{8'd0,8'd108} : s = 332;
	{8'd0,8'd109} : s = 453;
	{8'd0,8'd110} : s = 451;
	{8'd0,8'd111} : s = 498;
	{8'd0,8'd112} : s = 176;
	{8'd0,8'd113} : s = 330;
	{8'd0,8'd114} : s = 329;
	{8'd0,8'd115} : s = 440;
	{8'd0,8'd116} : s = 326;
	{8'd0,8'd117} : s = 436;
	{8'd0,8'd118} : s = 434;
	{8'd0,8'd119} : s = 497;
	{8'd0,8'd120} : s = 325;
	{8'd0,8'd121} : s = 433;
	{8'd0,8'd122} : s = 428;
	{8'd0,8'd123} : s = 492;
	{8'd0,8'd124} : s = 426;
	{8'd0,8'd125} : s = 490;
	{8'd0,8'd126} : s = 489;
	{8'd0,8'd127} : s = 508;
	{8'd0,8'd128} : s = 2;
	{8'd0,8'd129} : s = 48;
	{8'd0,8'd130} : s = 40;
	{8'd0,8'd131} : s = 168;
	{8'd0,8'd132} : s = 36;
	{8'd0,8'd133} : s = 164;
	{8'd0,8'd134} : s = 162;
	{8'd0,8'd135} : s = 323;
	{8'd0,8'd136} : s = 34;
	{8'd0,8'd137} : s = 161;
	{8'd0,8'd138} : s = 152;
	{8'd0,8'd139} : s = 312;
	{8'd0,8'd140} : s = 148;
	{8'd0,8'd141} : s = 308;
	{8'd0,8'd142} : s = 306;
	{8'd0,8'd143} : s = 425;
	{8'd0,8'd144} : s = 33;
	{8'd0,8'd145} : s = 146;
	{8'd0,8'd146} : s = 145;
	{8'd0,8'd147} : s = 305;
	{8'd0,8'd148} : s = 140;
	{8'd0,8'd149} : s = 300;
	{8'd0,8'd150} : s = 298;
	{8'd0,8'd151} : s = 422;
	{8'd0,8'd152} : s = 138;
	{8'd0,8'd153} : s = 297;
	{8'd0,8'd154} : s = 294;
	{8'd0,8'd155} : s = 421;
	{8'd0,8'd156} : s = 293;
	{8'd0,8'd157} : s = 419;
	{8'd0,8'd158} : s = 412;
	{8'd0,8'd159} : s = 486;
	{8'd0,8'd160} : s = 24;
	{8'd0,8'd161} : s = 137;
	{8'd0,8'd162} : s = 134;
	{8'd0,8'd163} : s = 291;
	{8'd0,8'd164} : s = 133;
	{8'd0,8'd165} : s = 284;
	{8'd0,8'd166} : s = 282;
	{8'd0,8'd167} : s = 410;
	{8'd0,8'd168} : s = 131;
	{8'd0,8'd169} : s = 281;
	{8'd0,8'd170} : s = 278;
	{8'd0,8'd171} : s = 409;
	{8'd0,8'd172} : s = 277;
	{8'd0,8'd173} : s = 406;
	{8'd0,8'd174} : s = 405;
	{8'd0,8'd175} : s = 485;
	{8'd0,8'd176} : s = 112;
	{8'd0,8'd177} : s = 275;
	{8'd0,8'd178} : s = 270;
	{8'd0,8'd179} : s = 403;
	{8'd0,8'd180} : s = 269;
	{8'd0,8'd181} : s = 398;
	{8'd0,8'd182} : s = 397;
	{8'd0,8'd183} : s = 483;
	{8'd0,8'd184} : s = 267;
	{8'd0,8'd185} : s = 395;
	{8'd0,8'd186} : s = 391;
	{8'd0,8'd187} : s = 476;
	{8'd0,8'd188} : s = 376;
	{8'd0,8'd189} : s = 474;
	{8'd0,8'd190} : s = 473;
	{8'd0,8'd191} : s = 506;
	{8'd0,8'd192} : s = 20;
	{8'd0,8'd193} : s = 104;
	{8'd0,8'd194} : s = 100;
	{8'd0,8'd195} : s = 263;
	{8'd0,8'd196} : s = 98;
	{8'd0,8'd197} : s = 240;
	{8'd0,8'd198} : s = 232;
	{8'd0,8'd199} : s = 372;
	{8'd0,8'd200} : s = 97;
	{8'd0,8'd201} : s = 228;
	{8'd0,8'd202} : s = 226;
	{8'd0,8'd203} : s = 370;
	{8'd0,8'd204} : s = 225;
	{8'd0,8'd205} : s = 369;
	{8'd0,8'd206} : s = 364;
	{8'd0,8'd207} : s = 470;
	{8'd0,8'd208} : s = 88;
	{8'd0,8'd209} : s = 216;
	{8'd0,8'd210} : s = 212;
	{8'd0,8'd211} : s = 362;
	{8'd0,8'd212} : s = 210;
	{8'd0,8'd213} : s = 361;
	{8'd0,8'd214} : s = 358;
	{8'd0,8'd215} : s = 469;
	{8'd0,8'd216} : s = 209;
	{8'd0,8'd217} : s = 357;
	{8'd0,8'd218} : s = 355;
	{8'd0,8'd219} : s = 467;
	{8'd0,8'd220} : s = 348;
	{8'd0,8'd221} : s = 462;
	{8'd0,8'd222} : s = 461;
	{8'd0,8'd223} : s = 505;
	{8'd0,8'd224} : s = 84;
	{8'd0,8'd225} : s = 204;
	{8'd0,8'd226} : s = 202;
	{8'd0,8'd227} : s = 346;
	{8'd0,8'd228} : s = 201;
	{8'd0,8'd229} : s = 345;
	{8'd0,8'd230} : s = 342;
	{8'd0,8'd231} : s = 459;
	{8'd0,8'd232} : s = 198;
	{8'd0,8'd233} : s = 341;
	{8'd0,8'd234} : s = 339;
	{8'd0,8'd235} : s = 455;
	{8'd0,8'd236} : s = 334;
	{8'd0,8'd237} : s = 444;
	{8'd0,8'd238} : s = 442;
	{8'd0,8'd239} : s = 502;
	{8'd0,8'd240} : s = 197;
	{8'd0,8'd241} : s = 333;
	{8'd0,8'd242} : s = 331;
	{8'd0,8'd243} : s = 441;
	{8'd0,8'd244} : s = 327;
	{8'd0,8'd245} : s = 438;
	{8'd0,8'd246} : s = 437;
	{8'd0,8'd247} : s = 501;
	{8'd0,8'd248} : s = 316;
	{8'd0,8'd249} : s = 435;
	{8'd0,8'd250} : s = 430;
	{8'd0,8'd251} : s = 499;
	{8'd0,8'd252} : s = 429;
	{8'd0,8'd253} : s = 494;
	{8'd0,8'd254} : s = 493;
	{8'd0,8'd255} : s = 510;
	{8'd1,8'd0} : s = 256;
	{8'd1,8'd1} : s = 128;
	{8'd1,8'd2} : s = 384;
	{8'd1,8'd3} : s = 64;
	{8'd1,8'd4} : s = 320;
	{8'd1,8'd5} : s = 288;
	{8'd1,8'd6} : s = 448;
	{8'd1,8'd7} : s = 32;
	{8'd1,8'd8} : s = 272;
	{8'd1,8'd9} : s = 264;
	{8'd1,8'd10} : s = 416;
	{8'd1,8'd11} : s = 260;
	{8'd1,8'd12} : s = 400;
	{8'd1,8'd13} : s = 392;
	{8'd1,8'd14} : s = 480;
	{8'd1,8'd15} : s = 8;
	{8'd1,8'd16} : s = 258;
	{8'd1,8'd17} : s = 257;
	{8'd1,8'd18} : s = 388;
	{8'd1,8'd19} : s = 192;
	{8'd1,8'd20} : s = 386;
	{8'd1,8'd21} : s = 385;
	{8'd1,8'd22} : s = 464;
	{8'd1,8'd23} : s = 160;
	{8'd1,8'd24} : s = 352;
	{8'd1,8'd25} : s = 336;
	{8'd1,8'd26} : s = 456;
	{8'd1,8'd27} : s = 328;
	{8'd1,8'd28} : s = 452;
	{8'd1,8'd29} : s = 450;
	{8'd1,8'd30} : s = 496;
	{8'd1,8'd31} : s = 16;
	{8'd1,8'd32} : s = 144;
	{8'd1,8'd33} : s = 136;
	{8'd1,8'd34} : s = 324;
	{8'd1,8'd35} : s = 132;
	{8'd1,8'd36} : s = 322;
	{8'd1,8'd37} : s = 321;
	{8'd1,8'd38} : s = 449;
	{8'd1,8'd39} : s = 130;
	{8'd1,8'd40} : s = 304;
	{8'd1,8'd41} : s = 296;
	{8'd1,8'd42} : s = 432;
	{8'd1,8'd43} : s = 292;
	{8'd1,8'd44} : s = 424;
	{8'd1,8'd45} : s = 420;
	{8'd1,8'd46} : s = 488;
	{8'd1,8'd47} : s = 129;
	{8'd1,8'd48} : s = 290;
	{8'd1,8'd49} : s = 289;
	{8'd1,8'd50} : s = 418;
	{8'd1,8'd51} : s = 280;
	{8'd1,8'd52} : s = 417;
	{8'd1,8'd53} : s = 408;
	{8'd1,8'd54} : s = 484;
	{8'd1,8'd55} : s = 276;
	{8'd1,8'd56} : s = 404;
	{8'd1,8'd57} : s = 402;
	{8'd1,8'd58} : s = 482;
	{8'd1,8'd59} : s = 401;
	{8'd1,8'd60} : s = 481;
	{8'd1,8'd61} : s = 472;
	{8'd1,8'd62} : s = 504;
	{8'd1,8'd63} : s = 4;
	{8'd1,8'd64} : s = 96;
	{8'd1,8'd65} : s = 80;
	{8'd1,8'd66} : s = 274;
	{8'd1,8'd67} : s = 72;
	{8'd1,8'd68} : s = 273;
	{8'd1,8'd69} : s = 268;
	{8'd1,8'd70} : s = 396;
	{8'd1,8'd71} : s = 68;
	{8'd1,8'd72} : s = 266;
	{8'd1,8'd73} : s = 265;
	{8'd1,8'd74} : s = 394;
	{8'd1,8'd75} : s = 262;
	{8'd1,8'd76} : s = 393;
	{8'd1,8'd77} : s = 390;
	{8'd1,8'd78} : s = 468;
	{8'd1,8'd79} : s = 66;
	{8'd1,8'd80} : s = 261;
	{8'd1,8'd81} : s = 259;
	{8'd1,8'd82} : s = 389;
	{8'd1,8'd83} : s = 224;
	{8'd1,8'd84} : s = 387;
	{8'd1,8'd85} : s = 368;
	{8'd1,8'd86} : s = 466;
	{8'd1,8'd87} : s = 208;
	{8'd1,8'd88} : s = 360;
	{8'd1,8'd89} : s = 356;
	{8'd1,8'd90} : s = 465;
	{8'd1,8'd91} : s = 354;
	{8'd1,8'd92} : s = 460;
	{8'd1,8'd93} : s = 458;
	{8'd1,8'd94} : s = 500;
	{8'd1,8'd95} : s = 65;
	{8'd1,8'd96} : s = 200;
	{8'd1,8'd97} : s = 196;
	{8'd1,8'd98} : s = 353;
	{8'd1,8'd99} : s = 194;
	{8'd1,8'd100} : s = 344;
	{8'd1,8'd101} : s = 340;
	{8'd1,8'd102} : s = 457;
	{8'd1,8'd103} : s = 193;
	{8'd1,8'd104} : s = 338;
	{8'd1,8'd105} : s = 337;
	{8'd1,8'd106} : s = 454;
	{8'd1,8'd107} : s = 332;
	{8'd1,8'd108} : s = 453;
	{8'd1,8'd109} : s = 451;
	{8'd1,8'd110} : s = 498;
	{8'd1,8'd111} : s = 176;
	{8'd1,8'd112} : s = 330;
	{8'd1,8'd113} : s = 329;
	{8'd1,8'd114} : s = 440;
	{8'd1,8'd115} : s = 326;
	{8'd1,8'd116} : s = 436;
	{8'd1,8'd117} : s = 434;
	{8'd1,8'd118} : s = 497;
	{8'd1,8'd119} : s = 325;
	{8'd1,8'd120} : s = 433;
	{8'd1,8'd121} : s = 428;
	{8'd1,8'd122} : s = 492;
	{8'd1,8'd123} : s = 426;
	{8'd1,8'd124} : s = 490;
	{8'd1,8'd125} : s = 489;
	{8'd1,8'd126} : s = 508;
	{8'd1,8'd127} : s = 2;
	{8'd1,8'd128} : s = 48;
	{8'd1,8'd129} : s = 40;
	{8'd1,8'd130} : s = 168;
	{8'd1,8'd131} : s = 36;
	{8'd1,8'd132} : s = 164;
	{8'd1,8'd133} : s = 162;
	{8'd1,8'd134} : s = 323;
	{8'd1,8'd135} : s = 34;
	{8'd1,8'd136} : s = 161;
	{8'd1,8'd137} : s = 152;
	{8'd1,8'd138} : s = 312;
	{8'd1,8'd139} : s = 148;
	{8'd1,8'd140} : s = 308;
	{8'd1,8'd141} : s = 306;
	{8'd1,8'd142} : s = 425;
	{8'd1,8'd143} : s = 33;
	{8'd1,8'd144} : s = 146;
	{8'd1,8'd145} : s = 145;
	{8'd1,8'd146} : s = 305;
	{8'd1,8'd147} : s = 140;
	{8'd1,8'd148} : s = 300;
	{8'd1,8'd149} : s = 298;
	{8'd1,8'd150} : s = 422;
	{8'd1,8'd151} : s = 138;
	{8'd1,8'd152} : s = 297;
	{8'd1,8'd153} : s = 294;
	{8'd1,8'd154} : s = 421;
	{8'd1,8'd155} : s = 293;
	{8'd1,8'd156} : s = 419;
	{8'd1,8'd157} : s = 412;
	{8'd1,8'd158} : s = 486;
	{8'd1,8'd159} : s = 24;
	{8'd1,8'd160} : s = 137;
	{8'd1,8'd161} : s = 134;
	{8'd1,8'd162} : s = 291;
	{8'd1,8'd163} : s = 133;
	{8'd1,8'd164} : s = 284;
	{8'd1,8'd165} : s = 282;
	{8'd1,8'd166} : s = 410;
	{8'd1,8'd167} : s = 131;
	{8'd1,8'd168} : s = 281;
	{8'd1,8'd169} : s = 278;
	{8'd1,8'd170} : s = 409;
	{8'd1,8'd171} : s = 277;
	{8'd1,8'd172} : s = 406;
	{8'd1,8'd173} : s = 405;
	{8'd1,8'd174} : s = 485;
	{8'd1,8'd175} : s = 112;
	{8'd1,8'd176} : s = 275;
	{8'd1,8'd177} : s = 270;
	{8'd1,8'd178} : s = 403;
	{8'd1,8'd179} : s = 269;
	{8'd1,8'd180} : s = 398;
	{8'd1,8'd181} : s = 397;
	{8'd1,8'd182} : s = 483;
	{8'd1,8'd183} : s = 267;
	{8'd1,8'd184} : s = 395;
	{8'd1,8'd185} : s = 391;
	{8'd1,8'd186} : s = 476;
	{8'd1,8'd187} : s = 376;
	{8'd1,8'd188} : s = 474;
	{8'd1,8'd189} : s = 473;
	{8'd1,8'd190} : s = 506;
	{8'd1,8'd191} : s = 20;
	{8'd1,8'd192} : s = 104;
	{8'd1,8'd193} : s = 100;
	{8'd1,8'd194} : s = 263;
	{8'd1,8'd195} : s = 98;
	{8'd1,8'd196} : s = 240;
	{8'd1,8'd197} : s = 232;
	{8'd1,8'd198} : s = 372;
	{8'd1,8'd199} : s = 97;
	{8'd1,8'd200} : s = 228;
	{8'd1,8'd201} : s = 226;
	{8'd1,8'd202} : s = 370;
	{8'd1,8'd203} : s = 225;
	{8'd1,8'd204} : s = 369;
	{8'd1,8'd205} : s = 364;
	{8'd1,8'd206} : s = 470;
	{8'd1,8'd207} : s = 88;
	{8'd1,8'd208} : s = 216;
	{8'd1,8'd209} : s = 212;
	{8'd1,8'd210} : s = 362;
	{8'd1,8'd211} : s = 210;
	{8'd1,8'd212} : s = 361;
	{8'd1,8'd213} : s = 358;
	{8'd1,8'd214} : s = 469;
	{8'd1,8'd215} : s = 209;
	{8'd1,8'd216} : s = 357;
	{8'd1,8'd217} : s = 355;
	{8'd1,8'd218} : s = 467;
	{8'd1,8'd219} : s = 348;
	{8'd1,8'd220} : s = 462;
	{8'd1,8'd221} : s = 461;
	{8'd1,8'd222} : s = 505;
	{8'd1,8'd223} : s = 84;
	{8'd1,8'd224} : s = 204;
	{8'd1,8'd225} : s = 202;
	{8'd1,8'd226} : s = 346;
	{8'd1,8'd227} : s = 201;
	{8'd1,8'd228} : s = 345;
	{8'd1,8'd229} : s = 342;
	{8'd1,8'd230} : s = 459;
	{8'd1,8'd231} : s = 198;
	{8'd1,8'd232} : s = 341;
	{8'd1,8'd233} : s = 339;
	{8'd1,8'd234} : s = 455;
	{8'd1,8'd235} : s = 334;
	{8'd1,8'd236} : s = 444;
	{8'd1,8'd237} : s = 442;
	{8'd1,8'd238} : s = 502;
	{8'd1,8'd239} : s = 197;
	{8'd1,8'd240} : s = 333;
	{8'd1,8'd241} : s = 331;
	{8'd1,8'd242} : s = 441;
	{8'd1,8'd243} : s = 327;
	{8'd1,8'd244} : s = 438;
	{8'd1,8'd245} : s = 437;
	{8'd1,8'd246} : s = 501;
	{8'd1,8'd247} : s = 316;
	{8'd1,8'd248} : s = 435;
	{8'd1,8'd249} : s = 430;
	{8'd1,8'd250} : s = 499;
	{8'd1,8'd251} : s = 429;
	{8'd1,8'd252} : s = 494;
	{8'd1,8'd253} : s = 493;
	{8'd1,8'd254} : s = 510;
	{8'd1,8'd255} : s = 1;
	{8'd2,8'd0} : s = 128;
	{8'd2,8'd1} : s = 384;
	{8'd2,8'd2} : s = 64;
	{8'd2,8'd3} : s = 320;
	{8'd2,8'd4} : s = 288;
	{8'd2,8'd5} : s = 448;
	{8'd2,8'd6} : s = 32;
	{8'd2,8'd7} : s = 272;
	{8'd2,8'd8} : s = 264;
	{8'd2,8'd9} : s = 416;
	{8'd2,8'd10} : s = 260;
	{8'd2,8'd11} : s = 400;
	{8'd2,8'd12} : s = 392;
	{8'd2,8'd13} : s = 480;
	{8'd2,8'd14} : s = 8;
	{8'd2,8'd15} : s = 258;
	{8'd2,8'd16} : s = 257;
	{8'd2,8'd17} : s = 388;
	{8'd2,8'd18} : s = 192;
	{8'd2,8'd19} : s = 386;
	{8'd2,8'd20} : s = 385;
	{8'd2,8'd21} : s = 464;
	{8'd2,8'd22} : s = 160;
	{8'd2,8'd23} : s = 352;
	{8'd2,8'd24} : s = 336;
	{8'd2,8'd25} : s = 456;
	{8'd2,8'd26} : s = 328;
	{8'd2,8'd27} : s = 452;
	{8'd2,8'd28} : s = 450;
	{8'd2,8'd29} : s = 496;
	{8'd2,8'd30} : s = 16;
	{8'd2,8'd31} : s = 144;
	{8'd2,8'd32} : s = 136;
	{8'd2,8'd33} : s = 324;
	{8'd2,8'd34} : s = 132;
	{8'd2,8'd35} : s = 322;
	{8'd2,8'd36} : s = 321;
	{8'd2,8'd37} : s = 449;
	{8'd2,8'd38} : s = 130;
	{8'd2,8'd39} : s = 304;
	{8'd2,8'd40} : s = 296;
	{8'd2,8'd41} : s = 432;
	{8'd2,8'd42} : s = 292;
	{8'd2,8'd43} : s = 424;
	{8'd2,8'd44} : s = 420;
	{8'd2,8'd45} : s = 488;
	{8'd2,8'd46} : s = 129;
	{8'd2,8'd47} : s = 290;
	{8'd2,8'd48} : s = 289;
	{8'd2,8'd49} : s = 418;
	{8'd2,8'd50} : s = 280;
	{8'd2,8'd51} : s = 417;
	{8'd2,8'd52} : s = 408;
	{8'd2,8'd53} : s = 484;
	{8'd2,8'd54} : s = 276;
	{8'd2,8'd55} : s = 404;
	{8'd2,8'd56} : s = 402;
	{8'd2,8'd57} : s = 482;
	{8'd2,8'd58} : s = 401;
	{8'd2,8'd59} : s = 481;
	{8'd2,8'd60} : s = 472;
	{8'd2,8'd61} : s = 504;
	{8'd2,8'd62} : s = 4;
	{8'd2,8'd63} : s = 96;
	{8'd2,8'd64} : s = 80;
	{8'd2,8'd65} : s = 274;
	{8'd2,8'd66} : s = 72;
	{8'd2,8'd67} : s = 273;
	{8'd2,8'd68} : s = 268;
	{8'd2,8'd69} : s = 396;
	{8'd2,8'd70} : s = 68;
	{8'd2,8'd71} : s = 266;
	{8'd2,8'd72} : s = 265;
	{8'd2,8'd73} : s = 394;
	{8'd2,8'd74} : s = 262;
	{8'd2,8'd75} : s = 393;
	{8'd2,8'd76} : s = 390;
	{8'd2,8'd77} : s = 468;
	{8'd2,8'd78} : s = 66;
	{8'd2,8'd79} : s = 261;
	{8'd2,8'd80} : s = 259;
	{8'd2,8'd81} : s = 389;
	{8'd2,8'd82} : s = 224;
	{8'd2,8'd83} : s = 387;
	{8'd2,8'd84} : s = 368;
	{8'd2,8'd85} : s = 466;
	{8'd2,8'd86} : s = 208;
	{8'd2,8'd87} : s = 360;
	{8'd2,8'd88} : s = 356;
	{8'd2,8'd89} : s = 465;
	{8'd2,8'd90} : s = 354;
	{8'd2,8'd91} : s = 460;
	{8'd2,8'd92} : s = 458;
	{8'd2,8'd93} : s = 500;
	{8'd2,8'd94} : s = 65;
	{8'd2,8'd95} : s = 200;
	{8'd2,8'd96} : s = 196;
	{8'd2,8'd97} : s = 353;
	{8'd2,8'd98} : s = 194;
	{8'd2,8'd99} : s = 344;
	{8'd2,8'd100} : s = 340;
	{8'd2,8'd101} : s = 457;
	{8'd2,8'd102} : s = 193;
	{8'd2,8'd103} : s = 338;
	{8'd2,8'd104} : s = 337;
	{8'd2,8'd105} : s = 454;
	{8'd2,8'd106} : s = 332;
	{8'd2,8'd107} : s = 453;
	{8'd2,8'd108} : s = 451;
	{8'd2,8'd109} : s = 498;
	{8'd2,8'd110} : s = 176;
	{8'd2,8'd111} : s = 330;
	{8'd2,8'd112} : s = 329;
	{8'd2,8'd113} : s = 440;
	{8'd2,8'd114} : s = 326;
	{8'd2,8'd115} : s = 436;
	{8'd2,8'd116} : s = 434;
	{8'd2,8'd117} : s = 497;
	{8'd2,8'd118} : s = 325;
	{8'd2,8'd119} : s = 433;
	{8'd2,8'd120} : s = 428;
	{8'd2,8'd121} : s = 492;
	{8'd2,8'd122} : s = 426;
	{8'd2,8'd123} : s = 490;
	{8'd2,8'd124} : s = 489;
	{8'd2,8'd125} : s = 508;
	{8'd2,8'd126} : s = 2;
	{8'd2,8'd127} : s = 48;
	{8'd2,8'd128} : s = 40;
	{8'd2,8'd129} : s = 168;
	{8'd2,8'd130} : s = 36;
	{8'd2,8'd131} : s = 164;
	{8'd2,8'd132} : s = 162;
	{8'd2,8'd133} : s = 323;
	{8'd2,8'd134} : s = 34;
	{8'd2,8'd135} : s = 161;
	{8'd2,8'd136} : s = 152;
	{8'd2,8'd137} : s = 312;
	{8'd2,8'd138} : s = 148;
	{8'd2,8'd139} : s = 308;
	{8'd2,8'd140} : s = 306;
	{8'd2,8'd141} : s = 425;
	{8'd2,8'd142} : s = 33;
	{8'd2,8'd143} : s = 146;
	{8'd2,8'd144} : s = 145;
	{8'd2,8'd145} : s = 305;
	{8'd2,8'd146} : s = 140;
	{8'd2,8'd147} : s = 300;
	{8'd2,8'd148} : s = 298;
	{8'd2,8'd149} : s = 422;
	{8'd2,8'd150} : s = 138;
	{8'd2,8'd151} : s = 297;
	{8'd2,8'd152} : s = 294;
	{8'd2,8'd153} : s = 421;
	{8'd2,8'd154} : s = 293;
	{8'd2,8'd155} : s = 419;
	{8'd2,8'd156} : s = 412;
	{8'd2,8'd157} : s = 486;
	{8'd2,8'd158} : s = 24;
	{8'd2,8'd159} : s = 137;
	{8'd2,8'd160} : s = 134;
	{8'd2,8'd161} : s = 291;
	{8'd2,8'd162} : s = 133;
	{8'd2,8'd163} : s = 284;
	{8'd2,8'd164} : s = 282;
	{8'd2,8'd165} : s = 410;
	{8'd2,8'd166} : s = 131;
	{8'd2,8'd167} : s = 281;
	{8'd2,8'd168} : s = 278;
	{8'd2,8'd169} : s = 409;
	{8'd2,8'd170} : s = 277;
	{8'd2,8'd171} : s = 406;
	{8'd2,8'd172} : s = 405;
	{8'd2,8'd173} : s = 485;
	{8'd2,8'd174} : s = 112;
	{8'd2,8'd175} : s = 275;
	{8'd2,8'd176} : s = 270;
	{8'd2,8'd177} : s = 403;
	{8'd2,8'd178} : s = 269;
	{8'd2,8'd179} : s = 398;
	{8'd2,8'd180} : s = 397;
	{8'd2,8'd181} : s = 483;
	{8'd2,8'd182} : s = 267;
	{8'd2,8'd183} : s = 395;
	{8'd2,8'd184} : s = 391;
	{8'd2,8'd185} : s = 476;
	{8'd2,8'd186} : s = 376;
	{8'd2,8'd187} : s = 474;
	{8'd2,8'd188} : s = 473;
	{8'd2,8'd189} : s = 506;
	{8'd2,8'd190} : s = 20;
	{8'd2,8'd191} : s = 104;
	{8'd2,8'd192} : s = 100;
	{8'd2,8'd193} : s = 263;
	{8'd2,8'd194} : s = 98;
	{8'd2,8'd195} : s = 240;
	{8'd2,8'd196} : s = 232;
	{8'd2,8'd197} : s = 372;
	{8'd2,8'd198} : s = 97;
	{8'd2,8'd199} : s = 228;
	{8'd2,8'd200} : s = 226;
	{8'd2,8'd201} : s = 370;
	{8'd2,8'd202} : s = 225;
	{8'd2,8'd203} : s = 369;
	{8'd2,8'd204} : s = 364;
	{8'd2,8'd205} : s = 470;
	{8'd2,8'd206} : s = 88;
	{8'd2,8'd207} : s = 216;
	{8'd2,8'd208} : s = 212;
	{8'd2,8'd209} : s = 362;
	{8'd2,8'd210} : s = 210;
	{8'd2,8'd211} : s = 361;
	{8'd2,8'd212} : s = 358;
	{8'd2,8'd213} : s = 469;
	{8'd2,8'd214} : s = 209;
	{8'd2,8'd215} : s = 357;
	{8'd2,8'd216} : s = 355;
	{8'd2,8'd217} : s = 467;
	{8'd2,8'd218} : s = 348;
	{8'd2,8'd219} : s = 462;
	{8'd2,8'd220} : s = 461;
	{8'd2,8'd221} : s = 505;
	{8'd2,8'd222} : s = 84;
	{8'd2,8'd223} : s = 204;
	{8'd2,8'd224} : s = 202;
	{8'd2,8'd225} : s = 346;
	{8'd2,8'd226} : s = 201;
	{8'd2,8'd227} : s = 345;
	{8'd2,8'd228} : s = 342;
	{8'd2,8'd229} : s = 459;
	{8'd2,8'd230} : s = 198;
	{8'd2,8'd231} : s = 341;
	{8'd2,8'd232} : s = 339;
	{8'd2,8'd233} : s = 455;
	{8'd2,8'd234} : s = 334;
	{8'd2,8'd235} : s = 444;
	{8'd2,8'd236} : s = 442;
	{8'd2,8'd237} : s = 502;
	{8'd2,8'd238} : s = 197;
	{8'd2,8'd239} : s = 333;
	{8'd2,8'd240} : s = 331;
	{8'd2,8'd241} : s = 441;
	{8'd2,8'd242} : s = 327;
	{8'd2,8'd243} : s = 438;
	{8'd2,8'd244} : s = 437;
	{8'd2,8'd245} : s = 501;
	{8'd2,8'd246} : s = 316;
	{8'd2,8'd247} : s = 435;
	{8'd2,8'd248} : s = 430;
	{8'd2,8'd249} : s = 499;
	{8'd2,8'd250} : s = 429;
	{8'd2,8'd251} : s = 494;
	{8'd2,8'd252} : s = 493;
	{8'd2,8'd253} : s = 510;
	{8'd2,8'd254} : s = 1;
	{8'd2,8'd255} : s = 18;
	{8'd3,8'd0} : s = 384;
	{8'd3,8'd1} : s = 64;
	{8'd3,8'd2} : s = 320;
	{8'd3,8'd3} : s = 288;
	{8'd3,8'd4} : s = 448;
	{8'd3,8'd5} : s = 32;
	{8'd3,8'd6} : s = 272;
	{8'd3,8'd7} : s = 264;
	{8'd3,8'd8} : s = 416;
	{8'd3,8'd9} : s = 260;
	{8'd3,8'd10} : s = 400;
	{8'd3,8'd11} : s = 392;
	{8'd3,8'd12} : s = 480;
	{8'd3,8'd13} : s = 8;
	{8'd3,8'd14} : s = 258;
	{8'd3,8'd15} : s = 257;
	{8'd3,8'd16} : s = 388;
	{8'd3,8'd17} : s = 192;
	{8'd3,8'd18} : s = 386;
	{8'd3,8'd19} : s = 385;
	{8'd3,8'd20} : s = 464;
	{8'd3,8'd21} : s = 160;
	{8'd3,8'd22} : s = 352;
	{8'd3,8'd23} : s = 336;
	{8'd3,8'd24} : s = 456;
	{8'd3,8'd25} : s = 328;
	{8'd3,8'd26} : s = 452;
	{8'd3,8'd27} : s = 450;
	{8'd3,8'd28} : s = 496;
	{8'd3,8'd29} : s = 16;
	{8'd3,8'd30} : s = 144;
	{8'd3,8'd31} : s = 136;
	{8'd3,8'd32} : s = 324;
	{8'd3,8'd33} : s = 132;
	{8'd3,8'd34} : s = 322;
	{8'd3,8'd35} : s = 321;
	{8'd3,8'd36} : s = 449;
	{8'd3,8'd37} : s = 130;
	{8'd3,8'd38} : s = 304;
	{8'd3,8'd39} : s = 296;
	{8'd3,8'd40} : s = 432;
	{8'd3,8'd41} : s = 292;
	{8'd3,8'd42} : s = 424;
	{8'd3,8'd43} : s = 420;
	{8'd3,8'd44} : s = 488;
	{8'd3,8'd45} : s = 129;
	{8'd3,8'd46} : s = 290;
	{8'd3,8'd47} : s = 289;
	{8'd3,8'd48} : s = 418;
	{8'd3,8'd49} : s = 280;
	{8'd3,8'd50} : s = 417;
	{8'd3,8'd51} : s = 408;
	{8'd3,8'd52} : s = 484;
	{8'd3,8'd53} : s = 276;
	{8'd3,8'd54} : s = 404;
	{8'd3,8'd55} : s = 402;
	{8'd3,8'd56} : s = 482;
	{8'd3,8'd57} : s = 401;
	{8'd3,8'd58} : s = 481;
	{8'd3,8'd59} : s = 472;
	{8'd3,8'd60} : s = 504;
	{8'd3,8'd61} : s = 4;
	{8'd3,8'd62} : s = 96;
	{8'd3,8'd63} : s = 80;
	{8'd3,8'd64} : s = 274;
	{8'd3,8'd65} : s = 72;
	{8'd3,8'd66} : s = 273;
	{8'd3,8'd67} : s = 268;
	{8'd3,8'd68} : s = 396;
	{8'd3,8'd69} : s = 68;
	{8'd3,8'd70} : s = 266;
	{8'd3,8'd71} : s = 265;
	{8'd3,8'd72} : s = 394;
	{8'd3,8'd73} : s = 262;
	{8'd3,8'd74} : s = 393;
	{8'd3,8'd75} : s = 390;
	{8'd3,8'd76} : s = 468;
	{8'd3,8'd77} : s = 66;
	{8'd3,8'd78} : s = 261;
	{8'd3,8'd79} : s = 259;
	{8'd3,8'd80} : s = 389;
	{8'd3,8'd81} : s = 224;
	{8'd3,8'd82} : s = 387;
	{8'd3,8'd83} : s = 368;
	{8'd3,8'd84} : s = 466;
	{8'd3,8'd85} : s = 208;
	{8'd3,8'd86} : s = 360;
	{8'd3,8'd87} : s = 356;
	{8'd3,8'd88} : s = 465;
	{8'd3,8'd89} : s = 354;
	{8'd3,8'd90} : s = 460;
	{8'd3,8'd91} : s = 458;
	{8'd3,8'd92} : s = 500;
	{8'd3,8'd93} : s = 65;
	{8'd3,8'd94} : s = 200;
	{8'd3,8'd95} : s = 196;
	{8'd3,8'd96} : s = 353;
	{8'd3,8'd97} : s = 194;
	{8'd3,8'd98} : s = 344;
	{8'd3,8'd99} : s = 340;
	{8'd3,8'd100} : s = 457;
	{8'd3,8'd101} : s = 193;
	{8'd3,8'd102} : s = 338;
	{8'd3,8'd103} : s = 337;
	{8'd3,8'd104} : s = 454;
	{8'd3,8'd105} : s = 332;
	{8'd3,8'd106} : s = 453;
	{8'd3,8'd107} : s = 451;
	{8'd3,8'd108} : s = 498;
	{8'd3,8'd109} : s = 176;
	{8'd3,8'd110} : s = 330;
	{8'd3,8'd111} : s = 329;
	{8'd3,8'd112} : s = 440;
	{8'd3,8'd113} : s = 326;
	{8'd3,8'd114} : s = 436;
	{8'd3,8'd115} : s = 434;
	{8'd3,8'd116} : s = 497;
	{8'd3,8'd117} : s = 325;
	{8'd3,8'd118} : s = 433;
	{8'd3,8'd119} : s = 428;
	{8'd3,8'd120} : s = 492;
	{8'd3,8'd121} : s = 426;
	{8'd3,8'd122} : s = 490;
	{8'd3,8'd123} : s = 489;
	{8'd3,8'd124} : s = 508;
	{8'd3,8'd125} : s = 2;
	{8'd3,8'd126} : s = 48;
	{8'd3,8'd127} : s = 40;
	{8'd3,8'd128} : s = 168;
	{8'd3,8'd129} : s = 36;
	{8'd3,8'd130} : s = 164;
	{8'd3,8'd131} : s = 162;
	{8'd3,8'd132} : s = 323;
	{8'd3,8'd133} : s = 34;
	{8'd3,8'd134} : s = 161;
	{8'd3,8'd135} : s = 152;
	{8'd3,8'd136} : s = 312;
	{8'd3,8'd137} : s = 148;
	{8'd3,8'd138} : s = 308;
	{8'd3,8'd139} : s = 306;
	{8'd3,8'd140} : s = 425;
	{8'd3,8'd141} : s = 33;
	{8'd3,8'd142} : s = 146;
	{8'd3,8'd143} : s = 145;
	{8'd3,8'd144} : s = 305;
	{8'd3,8'd145} : s = 140;
	{8'd3,8'd146} : s = 300;
	{8'd3,8'd147} : s = 298;
	{8'd3,8'd148} : s = 422;
	{8'd3,8'd149} : s = 138;
	{8'd3,8'd150} : s = 297;
	{8'd3,8'd151} : s = 294;
	{8'd3,8'd152} : s = 421;
	{8'd3,8'd153} : s = 293;
	{8'd3,8'd154} : s = 419;
	{8'd3,8'd155} : s = 412;
	{8'd3,8'd156} : s = 486;
	{8'd3,8'd157} : s = 24;
	{8'd3,8'd158} : s = 137;
	{8'd3,8'd159} : s = 134;
	{8'd3,8'd160} : s = 291;
	{8'd3,8'd161} : s = 133;
	{8'd3,8'd162} : s = 284;
	{8'd3,8'd163} : s = 282;
	{8'd3,8'd164} : s = 410;
	{8'd3,8'd165} : s = 131;
	{8'd3,8'd166} : s = 281;
	{8'd3,8'd167} : s = 278;
	{8'd3,8'd168} : s = 409;
	{8'd3,8'd169} : s = 277;
	{8'd3,8'd170} : s = 406;
	{8'd3,8'd171} : s = 405;
	{8'd3,8'd172} : s = 485;
	{8'd3,8'd173} : s = 112;
	{8'd3,8'd174} : s = 275;
	{8'd3,8'd175} : s = 270;
	{8'd3,8'd176} : s = 403;
	{8'd3,8'd177} : s = 269;
	{8'd3,8'd178} : s = 398;
	{8'd3,8'd179} : s = 397;
	{8'd3,8'd180} : s = 483;
	{8'd3,8'd181} : s = 267;
	{8'd3,8'd182} : s = 395;
	{8'd3,8'd183} : s = 391;
	{8'd3,8'd184} : s = 476;
	{8'd3,8'd185} : s = 376;
	{8'd3,8'd186} : s = 474;
	{8'd3,8'd187} : s = 473;
	{8'd3,8'd188} : s = 506;
	{8'd3,8'd189} : s = 20;
	{8'd3,8'd190} : s = 104;
	{8'd3,8'd191} : s = 100;
	{8'd3,8'd192} : s = 263;
	{8'd3,8'd193} : s = 98;
	{8'd3,8'd194} : s = 240;
	{8'd3,8'd195} : s = 232;
	{8'd3,8'd196} : s = 372;
	{8'd3,8'd197} : s = 97;
	{8'd3,8'd198} : s = 228;
	{8'd3,8'd199} : s = 226;
	{8'd3,8'd200} : s = 370;
	{8'd3,8'd201} : s = 225;
	{8'd3,8'd202} : s = 369;
	{8'd3,8'd203} : s = 364;
	{8'd3,8'd204} : s = 470;
	{8'd3,8'd205} : s = 88;
	{8'd3,8'd206} : s = 216;
	{8'd3,8'd207} : s = 212;
	{8'd3,8'd208} : s = 362;
	{8'd3,8'd209} : s = 210;
	{8'd3,8'd210} : s = 361;
	{8'd3,8'd211} : s = 358;
	{8'd3,8'd212} : s = 469;
	{8'd3,8'd213} : s = 209;
	{8'd3,8'd214} : s = 357;
	{8'd3,8'd215} : s = 355;
	{8'd3,8'd216} : s = 467;
	{8'd3,8'd217} : s = 348;
	{8'd3,8'd218} : s = 462;
	{8'd3,8'd219} : s = 461;
	{8'd3,8'd220} : s = 505;
	{8'd3,8'd221} : s = 84;
	{8'd3,8'd222} : s = 204;
	{8'd3,8'd223} : s = 202;
	{8'd3,8'd224} : s = 346;
	{8'd3,8'd225} : s = 201;
	{8'd3,8'd226} : s = 345;
	{8'd3,8'd227} : s = 342;
	{8'd3,8'd228} : s = 459;
	{8'd3,8'd229} : s = 198;
	{8'd3,8'd230} : s = 341;
	{8'd3,8'd231} : s = 339;
	{8'd3,8'd232} : s = 455;
	{8'd3,8'd233} : s = 334;
	{8'd3,8'd234} : s = 444;
	{8'd3,8'd235} : s = 442;
	{8'd3,8'd236} : s = 502;
	{8'd3,8'd237} : s = 197;
	{8'd3,8'd238} : s = 333;
	{8'd3,8'd239} : s = 331;
	{8'd3,8'd240} : s = 441;
	{8'd3,8'd241} : s = 327;
	{8'd3,8'd242} : s = 438;
	{8'd3,8'd243} : s = 437;
	{8'd3,8'd244} : s = 501;
	{8'd3,8'd245} : s = 316;
	{8'd3,8'd246} : s = 435;
	{8'd3,8'd247} : s = 430;
	{8'd3,8'd248} : s = 499;
	{8'd3,8'd249} : s = 429;
	{8'd3,8'd250} : s = 494;
	{8'd3,8'd251} : s = 493;
	{8'd3,8'd252} : s = 510;
	{8'd3,8'd253} : s = 1;
	{8'd3,8'd254} : s = 18;
	{8'd3,8'd255} : s = 17;
	{8'd4,8'd0} : s = 64;
	{8'd4,8'd1} : s = 320;
	{8'd4,8'd2} : s = 288;
	{8'd4,8'd3} : s = 448;
	{8'd4,8'd4} : s = 32;
	{8'd4,8'd5} : s = 272;
	{8'd4,8'd6} : s = 264;
	{8'd4,8'd7} : s = 416;
	{8'd4,8'd8} : s = 260;
	{8'd4,8'd9} : s = 400;
	{8'd4,8'd10} : s = 392;
	{8'd4,8'd11} : s = 480;
	{8'd4,8'd12} : s = 8;
	{8'd4,8'd13} : s = 258;
	{8'd4,8'd14} : s = 257;
	{8'd4,8'd15} : s = 388;
	{8'd4,8'd16} : s = 192;
	{8'd4,8'd17} : s = 386;
	{8'd4,8'd18} : s = 385;
	{8'd4,8'd19} : s = 464;
	{8'd4,8'd20} : s = 160;
	{8'd4,8'd21} : s = 352;
	{8'd4,8'd22} : s = 336;
	{8'd4,8'd23} : s = 456;
	{8'd4,8'd24} : s = 328;
	{8'd4,8'd25} : s = 452;
	{8'd4,8'd26} : s = 450;
	{8'd4,8'd27} : s = 496;
	{8'd4,8'd28} : s = 16;
	{8'd4,8'd29} : s = 144;
	{8'd4,8'd30} : s = 136;
	{8'd4,8'd31} : s = 324;
	{8'd4,8'd32} : s = 132;
	{8'd4,8'd33} : s = 322;
	{8'd4,8'd34} : s = 321;
	{8'd4,8'd35} : s = 449;
	{8'd4,8'd36} : s = 130;
	{8'd4,8'd37} : s = 304;
	{8'd4,8'd38} : s = 296;
	{8'd4,8'd39} : s = 432;
	{8'd4,8'd40} : s = 292;
	{8'd4,8'd41} : s = 424;
	{8'd4,8'd42} : s = 420;
	{8'd4,8'd43} : s = 488;
	{8'd4,8'd44} : s = 129;
	{8'd4,8'd45} : s = 290;
	{8'd4,8'd46} : s = 289;
	{8'd4,8'd47} : s = 418;
	{8'd4,8'd48} : s = 280;
	{8'd4,8'd49} : s = 417;
	{8'd4,8'd50} : s = 408;
	{8'd4,8'd51} : s = 484;
	{8'd4,8'd52} : s = 276;
	{8'd4,8'd53} : s = 404;
	{8'd4,8'd54} : s = 402;
	{8'd4,8'd55} : s = 482;
	{8'd4,8'd56} : s = 401;
	{8'd4,8'd57} : s = 481;
	{8'd4,8'd58} : s = 472;
	{8'd4,8'd59} : s = 504;
	{8'd4,8'd60} : s = 4;
	{8'd4,8'd61} : s = 96;
	{8'd4,8'd62} : s = 80;
	{8'd4,8'd63} : s = 274;
	{8'd4,8'd64} : s = 72;
	{8'd4,8'd65} : s = 273;
	{8'd4,8'd66} : s = 268;
	{8'd4,8'd67} : s = 396;
	{8'd4,8'd68} : s = 68;
	{8'd4,8'd69} : s = 266;
	{8'd4,8'd70} : s = 265;
	{8'd4,8'd71} : s = 394;
	{8'd4,8'd72} : s = 262;
	{8'd4,8'd73} : s = 393;
	{8'd4,8'd74} : s = 390;
	{8'd4,8'd75} : s = 468;
	{8'd4,8'd76} : s = 66;
	{8'd4,8'd77} : s = 261;
	{8'd4,8'd78} : s = 259;
	{8'd4,8'd79} : s = 389;
	{8'd4,8'd80} : s = 224;
	{8'd4,8'd81} : s = 387;
	{8'd4,8'd82} : s = 368;
	{8'd4,8'd83} : s = 466;
	{8'd4,8'd84} : s = 208;
	{8'd4,8'd85} : s = 360;
	{8'd4,8'd86} : s = 356;
	{8'd4,8'd87} : s = 465;
	{8'd4,8'd88} : s = 354;
	{8'd4,8'd89} : s = 460;
	{8'd4,8'd90} : s = 458;
	{8'd4,8'd91} : s = 500;
	{8'd4,8'd92} : s = 65;
	{8'd4,8'd93} : s = 200;
	{8'd4,8'd94} : s = 196;
	{8'd4,8'd95} : s = 353;
	{8'd4,8'd96} : s = 194;
	{8'd4,8'd97} : s = 344;
	{8'd4,8'd98} : s = 340;
	{8'd4,8'd99} : s = 457;
	{8'd4,8'd100} : s = 193;
	{8'd4,8'd101} : s = 338;
	{8'd4,8'd102} : s = 337;
	{8'd4,8'd103} : s = 454;
	{8'd4,8'd104} : s = 332;
	{8'd4,8'd105} : s = 453;
	{8'd4,8'd106} : s = 451;
	{8'd4,8'd107} : s = 498;
	{8'd4,8'd108} : s = 176;
	{8'd4,8'd109} : s = 330;
	{8'd4,8'd110} : s = 329;
	{8'd4,8'd111} : s = 440;
	{8'd4,8'd112} : s = 326;
	{8'd4,8'd113} : s = 436;
	{8'd4,8'd114} : s = 434;
	{8'd4,8'd115} : s = 497;
	{8'd4,8'd116} : s = 325;
	{8'd4,8'd117} : s = 433;
	{8'd4,8'd118} : s = 428;
	{8'd4,8'd119} : s = 492;
	{8'd4,8'd120} : s = 426;
	{8'd4,8'd121} : s = 490;
	{8'd4,8'd122} : s = 489;
	{8'd4,8'd123} : s = 508;
	{8'd4,8'd124} : s = 2;
	{8'd4,8'd125} : s = 48;
	{8'd4,8'd126} : s = 40;
	{8'd4,8'd127} : s = 168;
	{8'd4,8'd128} : s = 36;
	{8'd4,8'd129} : s = 164;
	{8'd4,8'd130} : s = 162;
	{8'd4,8'd131} : s = 323;
	{8'd4,8'd132} : s = 34;
	{8'd4,8'd133} : s = 161;
	{8'd4,8'd134} : s = 152;
	{8'd4,8'd135} : s = 312;
	{8'd4,8'd136} : s = 148;
	{8'd4,8'd137} : s = 308;
	{8'd4,8'd138} : s = 306;
	{8'd4,8'd139} : s = 425;
	{8'd4,8'd140} : s = 33;
	{8'd4,8'd141} : s = 146;
	{8'd4,8'd142} : s = 145;
	{8'd4,8'd143} : s = 305;
	{8'd4,8'd144} : s = 140;
	{8'd4,8'd145} : s = 300;
	{8'd4,8'd146} : s = 298;
	{8'd4,8'd147} : s = 422;
	{8'd4,8'd148} : s = 138;
	{8'd4,8'd149} : s = 297;
	{8'd4,8'd150} : s = 294;
	{8'd4,8'd151} : s = 421;
	{8'd4,8'd152} : s = 293;
	{8'd4,8'd153} : s = 419;
	{8'd4,8'd154} : s = 412;
	{8'd4,8'd155} : s = 486;
	{8'd4,8'd156} : s = 24;
	{8'd4,8'd157} : s = 137;
	{8'd4,8'd158} : s = 134;
	{8'd4,8'd159} : s = 291;
	{8'd4,8'd160} : s = 133;
	{8'd4,8'd161} : s = 284;
	{8'd4,8'd162} : s = 282;
	{8'd4,8'd163} : s = 410;
	{8'd4,8'd164} : s = 131;
	{8'd4,8'd165} : s = 281;
	{8'd4,8'd166} : s = 278;
	{8'd4,8'd167} : s = 409;
	{8'd4,8'd168} : s = 277;
	{8'd4,8'd169} : s = 406;
	{8'd4,8'd170} : s = 405;
	{8'd4,8'd171} : s = 485;
	{8'd4,8'd172} : s = 112;
	{8'd4,8'd173} : s = 275;
	{8'd4,8'd174} : s = 270;
	{8'd4,8'd175} : s = 403;
	{8'd4,8'd176} : s = 269;
	{8'd4,8'd177} : s = 398;
	{8'd4,8'd178} : s = 397;
	{8'd4,8'd179} : s = 483;
	{8'd4,8'd180} : s = 267;
	{8'd4,8'd181} : s = 395;
	{8'd4,8'd182} : s = 391;
	{8'd4,8'd183} : s = 476;
	{8'd4,8'd184} : s = 376;
	{8'd4,8'd185} : s = 474;
	{8'd4,8'd186} : s = 473;
	{8'd4,8'd187} : s = 506;
	{8'd4,8'd188} : s = 20;
	{8'd4,8'd189} : s = 104;
	{8'd4,8'd190} : s = 100;
	{8'd4,8'd191} : s = 263;
	{8'd4,8'd192} : s = 98;
	{8'd4,8'd193} : s = 240;
	{8'd4,8'd194} : s = 232;
	{8'd4,8'd195} : s = 372;
	{8'd4,8'd196} : s = 97;
	{8'd4,8'd197} : s = 228;
	{8'd4,8'd198} : s = 226;
	{8'd4,8'd199} : s = 370;
	{8'd4,8'd200} : s = 225;
	{8'd4,8'd201} : s = 369;
	{8'd4,8'd202} : s = 364;
	{8'd4,8'd203} : s = 470;
	{8'd4,8'd204} : s = 88;
	{8'd4,8'd205} : s = 216;
	{8'd4,8'd206} : s = 212;
	{8'd4,8'd207} : s = 362;
	{8'd4,8'd208} : s = 210;
	{8'd4,8'd209} : s = 361;
	{8'd4,8'd210} : s = 358;
	{8'd4,8'd211} : s = 469;
	{8'd4,8'd212} : s = 209;
	{8'd4,8'd213} : s = 357;
	{8'd4,8'd214} : s = 355;
	{8'd4,8'd215} : s = 467;
	{8'd4,8'd216} : s = 348;
	{8'd4,8'd217} : s = 462;
	{8'd4,8'd218} : s = 461;
	{8'd4,8'd219} : s = 505;
	{8'd4,8'd220} : s = 84;
	{8'd4,8'd221} : s = 204;
	{8'd4,8'd222} : s = 202;
	{8'd4,8'd223} : s = 346;
	{8'd4,8'd224} : s = 201;
	{8'd4,8'd225} : s = 345;
	{8'd4,8'd226} : s = 342;
	{8'd4,8'd227} : s = 459;
	{8'd4,8'd228} : s = 198;
	{8'd4,8'd229} : s = 341;
	{8'd4,8'd230} : s = 339;
	{8'd4,8'd231} : s = 455;
	{8'd4,8'd232} : s = 334;
	{8'd4,8'd233} : s = 444;
	{8'd4,8'd234} : s = 442;
	{8'd4,8'd235} : s = 502;
	{8'd4,8'd236} : s = 197;
	{8'd4,8'd237} : s = 333;
	{8'd4,8'd238} : s = 331;
	{8'd4,8'd239} : s = 441;
	{8'd4,8'd240} : s = 327;
	{8'd4,8'd241} : s = 438;
	{8'd4,8'd242} : s = 437;
	{8'd4,8'd243} : s = 501;
	{8'd4,8'd244} : s = 316;
	{8'd4,8'd245} : s = 435;
	{8'd4,8'd246} : s = 430;
	{8'd4,8'd247} : s = 499;
	{8'd4,8'd248} : s = 429;
	{8'd4,8'd249} : s = 494;
	{8'd4,8'd250} : s = 493;
	{8'd4,8'd251} : s = 510;
	{8'd4,8'd252} : s = 1;
	{8'd4,8'd253} : s = 18;
	{8'd4,8'd254} : s = 17;
	{8'd4,8'd255} : s = 82;
	{8'd5,8'd0} : s = 320;
	{8'd5,8'd1} : s = 288;
	{8'd5,8'd2} : s = 448;
	{8'd5,8'd3} : s = 32;
	{8'd5,8'd4} : s = 272;
	{8'd5,8'd5} : s = 264;
	{8'd5,8'd6} : s = 416;
	{8'd5,8'd7} : s = 260;
	{8'd5,8'd8} : s = 400;
	{8'd5,8'd9} : s = 392;
	{8'd5,8'd10} : s = 480;
	{8'd5,8'd11} : s = 8;
	{8'd5,8'd12} : s = 258;
	{8'd5,8'd13} : s = 257;
	{8'd5,8'd14} : s = 388;
	{8'd5,8'd15} : s = 192;
	{8'd5,8'd16} : s = 386;
	{8'd5,8'd17} : s = 385;
	{8'd5,8'd18} : s = 464;
	{8'd5,8'd19} : s = 160;
	{8'd5,8'd20} : s = 352;
	{8'd5,8'd21} : s = 336;
	{8'd5,8'd22} : s = 456;
	{8'd5,8'd23} : s = 328;
	{8'd5,8'd24} : s = 452;
	{8'd5,8'd25} : s = 450;
	{8'd5,8'd26} : s = 496;
	{8'd5,8'd27} : s = 16;
	{8'd5,8'd28} : s = 144;
	{8'd5,8'd29} : s = 136;
	{8'd5,8'd30} : s = 324;
	{8'd5,8'd31} : s = 132;
	{8'd5,8'd32} : s = 322;
	{8'd5,8'd33} : s = 321;
	{8'd5,8'd34} : s = 449;
	{8'd5,8'd35} : s = 130;
	{8'd5,8'd36} : s = 304;
	{8'd5,8'd37} : s = 296;
	{8'd5,8'd38} : s = 432;
	{8'd5,8'd39} : s = 292;
	{8'd5,8'd40} : s = 424;
	{8'd5,8'd41} : s = 420;
	{8'd5,8'd42} : s = 488;
	{8'd5,8'd43} : s = 129;
	{8'd5,8'd44} : s = 290;
	{8'd5,8'd45} : s = 289;
	{8'd5,8'd46} : s = 418;
	{8'd5,8'd47} : s = 280;
	{8'd5,8'd48} : s = 417;
	{8'd5,8'd49} : s = 408;
	{8'd5,8'd50} : s = 484;
	{8'd5,8'd51} : s = 276;
	{8'd5,8'd52} : s = 404;
	{8'd5,8'd53} : s = 402;
	{8'd5,8'd54} : s = 482;
	{8'd5,8'd55} : s = 401;
	{8'd5,8'd56} : s = 481;
	{8'd5,8'd57} : s = 472;
	{8'd5,8'd58} : s = 504;
	{8'd5,8'd59} : s = 4;
	{8'd5,8'd60} : s = 96;
	{8'd5,8'd61} : s = 80;
	{8'd5,8'd62} : s = 274;
	{8'd5,8'd63} : s = 72;
	{8'd5,8'd64} : s = 273;
	{8'd5,8'd65} : s = 268;
	{8'd5,8'd66} : s = 396;
	{8'd5,8'd67} : s = 68;
	{8'd5,8'd68} : s = 266;
	{8'd5,8'd69} : s = 265;
	{8'd5,8'd70} : s = 394;
	{8'd5,8'd71} : s = 262;
	{8'd5,8'd72} : s = 393;
	{8'd5,8'd73} : s = 390;
	{8'd5,8'd74} : s = 468;
	{8'd5,8'd75} : s = 66;
	{8'd5,8'd76} : s = 261;
	{8'd5,8'd77} : s = 259;
	{8'd5,8'd78} : s = 389;
	{8'd5,8'd79} : s = 224;
	{8'd5,8'd80} : s = 387;
	{8'd5,8'd81} : s = 368;
	{8'd5,8'd82} : s = 466;
	{8'd5,8'd83} : s = 208;
	{8'd5,8'd84} : s = 360;
	{8'd5,8'd85} : s = 356;
	{8'd5,8'd86} : s = 465;
	{8'd5,8'd87} : s = 354;
	{8'd5,8'd88} : s = 460;
	{8'd5,8'd89} : s = 458;
	{8'd5,8'd90} : s = 500;
	{8'd5,8'd91} : s = 65;
	{8'd5,8'd92} : s = 200;
	{8'd5,8'd93} : s = 196;
	{8'd5,8'd94} : s = 353;
	{8'd5,8'd95} : s = 194;
	{8'd5,8'd96} : s = 344;
	{8'd5,8'd97} : s = 340;
	{8'd5,8'd98} : s = 457;
	{8'd5,8'd99} : s = 193;
	{8'd5,8'd100} : s = 338;
	{8'd5,8'd101} : s = 337;
	{8'd5,8'd102} : s = 454;
	{8'd5,8'd103} : s = 332;
	{8'd5,8'd104} : s = 453;
	{8'd5,8'd105} : s = 451;
	{8'd5,8'd106} : s = 498;
	{8'd5,8'd107} : s = 176;
	{8'd5,8'd108} : s = 330;
	{8'd5,8'd109} : s = 329;
	{8'd5,8'd110} : s = 440;
	{8'd5,8'd111} : s = 326;
	{8'd5,8'd112} : s = 436;
	{8'd5,8'd113} : s = 434;
	{8'd5,8'd114} : s = 497;
	{8'd5,8'd115} : s = 325;
	{8'd5,8'd116} : s = 433;
	{8'd5,8'd117} : s = 428;
	{8'd5,8'd118} : s = 492;
	{8'd5,8'd119} : s = 426;
	{8'd5,8'd120} : s = 490;
	{8'd5,8'd121} : s = 489;
	{8'd5,8'd122} : s = 508;
	{8'd5,8'd123} : s = 2;
	{8'd5,8'd124} : s = 48;
	{8'd5,8'd125} : s = 40;
	{8'd5,8'd126} : s = 168;
	{8'd5,8'd127} : s = 36;
	{8'd5,8'd128} : s = 164;
	{8'd5,8'd129} : s = 162;
	{8'd5,8'd130} : s = 323;
	{8'd5,8'd131} : s = 34;
	{8'd5,8'd132} : s = 161;
	{8'd5,8'd133} : s = 152;
	{8'd5,8'd134} : s = 312;
	{8'd5,8'd135} : s = 148;
	{8'd5,8'd136} : s = 308;
	{8'd5,8'd137} : s = 306;
	{8'd5,8'd138} : s = 425;
	{8'd5,8'd139} : s = 33;
	{8'd5,8'd140} : s = 146;
	{8'd5,8'd141} : s = 145;
	{8'd5,8'd142} : s = 305;
	{8'd5,8'd143} : s = 140;
	{8'd5,8'd144} : s = 300;
	{8'd5,8'd145} : s = 298;
	{8'd5,8'd146} : s = 422;
	{8'd5,8'd147} : s = 138;
	{8'd5,8'd148} : s = 297;
	{8'd5,8'd149} : s = 294;
	{8'd5,8'd150} : s = 421;
	{8'd5,8'd151} : s = 293;
	{8'd5,8'd152} : s = 419;
	{8'd5,8'd153} : s = 412;
	{8'd5,8'd154} : s = 486;
	{8'd5,8'd155} : s = 24;
	{8'd5,8'd156} : s = 137;
	{8'd5,8'd157} : s = 134;
	{8'd5,8'd158} : s = 291;
	{8'd5,8'd159} : s = 133;
	{8'd5,8'd160} : s = 284;
	{8'd5,8'd161} : s = 282;
	{8'd5,8'd162} : s = 410;
	{8'd5,8'd163} : s = 131;
	{8'd5,8'd164} : s = 281;
	{8'd5,8'd165} : s = 278;
	{8'd5,8'd166} : s = 409;
	{8'd5,8'd167} : s = 277;
	{8'd5,8'd168} : s = 406;
	{8'd5,8'd169} : s = 405;
	{8'd5,8'd170} : s = 485;
	{8'd5,8'd171} : s = 112;
	{8'd5,8'd172} : s = 275;
	{8'd5,8'd173} : s = 270;
	{8'd5,8'd174} : s = 403;
	{8'd5,8'd175} : s = 269;
	{8'd5,8'd176} : s = 398;
	{8'd5,8'd177} : s = 397;
	{8'd5,8'd178} : s = 483;
	{8'd5,8'd179} : s = 267;
	{8'd5,8'd180} : s = 395;
	{8'd5,8'd181} : s = 391;
	{8'd5,8'd182} : s = 476;
	{8'd5,8'd183} : s = 376;
	{8'd5,8'd184} : s = 474;
	{8'd5,8'd185} : s = 473;
	{8'd5,8'd186} : s = 506;
	{8'd5,8'd187} : s = 20;
	{8'd5,8'd188} : s = 104;
	{8'd5,8'd189} : s = 100;
	{8'd5,8'd190} : s = 263;
	{8'd5,8'd191} : s = 98;
	{8'd5,8'd192} : s = 240;
	{8'd5,8'd193} : s = 232;
	{8'd5,8'd194} : s = 372;
	{8'd5,8'd195} : s = 97;
	{8'd5,8'd196} : s = 228;
	{8'd5,8'd197} : s = 226;
	{8'd5,8'd198} : s = 370;
	{8'd5,8'd199} : s = 225;
	{8'd5,8'd200} : s = 369;
	{8'd5,8'd201} : s = 364;
	{8'd5,8'd202} : s = 470;
	{8'd5,8'd203} : s = 88;
	{8'd5,8'd204} : s = 216;
	{8'd5,8'd205} : s = 212;
	{8'd5,8'd206} : s = 362;
	{8'd5,8'd207} : s = 210;
	{8'd5,8'd208} : s = 361;
	{8'd5,8'd209} : s = 358;
	{8'd5,8'd210} : s = 469;
	{8'd5,8'd211} : s = 209;
	{8'd5,8'd212} : s = 357;
	{8'd5,8'd213} : s = 355;
	{8'd5,8'd214} : s = 467;
	{8'd5,8'd215} : s = 348;
	{8'd5,8'd216} : s = 462;
	{8'd5,8'd217} : s = 461;
	{8'd5,8'd218} : s = 505;
	{8'd5,8'd219} : s = 84;
	{8'd5,8'd220} : s = 204;
	{8'd5,8'd221} : s = 202;
	{8'd5,8'd222} : s = 346;
	{8'd5,8'd223} : s = 201;
	{8'd5,8'd224} : s = 345;
	{8'd5,8'd225} : s = 342;
	{8'd5,8'd226} : s = 459;
	{8'd5,8'd227} : s = 198;
	{8'd5,8'd228} : s = 341;
	{8'd5,8'd229} : s = 339;
	{8'd5,8'd230} : s = 455;
	{8'd5,8'd231} : s = 334;
	{8'd5,8'd232} : s = 444;
	{8'd5,8'd233} : s = 442;
	{8'd5,8'd234} : s = 502;
	{8'd5,8'd235} : s = 197;
	{8'd5,8'd236} : s = 333;
	{8'd5,8'd237} : s = 331;
	{8'd5,8'd238} : s = 441;
	{8'd5,8'd239} : s = 327;
	{8'd5,8'd240} : s = 438;
	{8'd5,8'd241} : s = 437;
	{8'd5,8'd242} : s = 501;
	{8'd5,8'd243} : s = 316;
	{8'd5,8'd244} : s = 435;
	{8'd5,8'd245} : s = 430;
	{8'd5,8'd246} : s = 499;
	{8'd5,8'd247} : s = 429;
	{8'd5,8'd248} : s = 494;
	{8'd5,8'd249} : s = 493;
	{8'd5,8'd250} : s = 510;
	{8'd5,8'd251} : s = 1;
	{8'd5,8'd252} : s = 18;
	{8'd5,8'd253} : s = 17;
	{8'd5,8'd254} : s = 82;
	{8'd5,8'd255} : s = 12;
	{8'd6,8'd0} : s = 288;
	{8'd6,8'd1} : s = 448;
	{8'd6,8'd2} : s = 32;
	{8'd6,8'd3} : s = 272;
	{8'd6,8'd4} : s = 264;
	{8'd6,8'd5} : s = 416;
	{8'd6,8'd6} : s = 260;
	{8'd6,8'd7} : s = 400;
	{8'd6,8'd8} : s = 392;
	{8'd6,8'd9} : s = 480;
	{8'd6,8'd10} : s = 8;
	{8'd6,8'd11} : s = 258;
	{8'd6,8'd12} : s = 257;
	{8'd6,8'd13} : s = 388;
	{8'd6,8'd14} : s = 192;
	{8'd6,8'd15} : s = 386;
	{8'd6,8'd16} : s = 385;
	{8'd6,8'd17} : s = 464;
	{8'd6,8'd18} : s = 160;
	{8'd6,8'd19} : s = 352;
	{8'd6,8'd20} : s = 336;
	{8'd6,8'd21} : s = 456;
	{8'd6,8'd22} : s = 328;
	{8'd6,8'd23} : s = 452;
	{8'd6,8'd24} : s = 450;
	{8'd6,8'd25} : s = 496;
	{8'd6,8'd26} : s = 16;
	{8'd6,8'd27} : s = 144;
	{8'd6,8'd28} : s = 136;
	{8'd6,8'd29} : s = 324;
	{8'd6,8'd30} : s = 132;
	{8'd6,8'd31} : s = 322;
	{8'd6,8'd32} : s = 321;
	{8'd6,8'd33} : s = 449;
	{8'd6,8'd34} : s = 130;
	{8'd6,8'd35} : s = 304;
	{8'd6,8'd36} : s = 296;
	{8'd6,8'd37} : s = 432;
	{8'd6,8'd38} : s = 292;
	{8'd6,8'd39} : s = 424;
	{8'd6,8'd40} : s = 420;
	{8'd6,8'd41} : s = 488;
	{8'd6,8'd42} : s = 129;
	{8'd6,8'd43} : s = 290;
	{8'd6,8'd44} : s = 289;
	{8'd6,8'd45} : s = 418;
	{8'd6,8'd46} : s = 280;
	{8'd6,8'd47} : s = 417;
	{8'd6,8'd48} : s = 408;
	{8'd6,8'd49} : s = 484;
	{8'd6,8'd50} : s = 276;
	{8'd6,8'd51} : s = 404;
	{8'd6,8'd52} : s = 402;
	{8'd6,8'd53} : s = 482;
	{8'd6,8'd54} : s = 401;
	{8'd6,8'd55} : s = 481;
	{8'd6,8'd56} : s = 472;
	{8'd6,8'd57} : s = 504;
	{8'd6,8'd58} : s = 4;
	{8'd6,8'd59} : s = 96;
	{8'd6,8'd60} : s = 80;
	{8'd6,8'd61} : s = 274;
	{8'd6,8'd62} : s = 72;
	{8'd6,8'd63} : s = 273;
	{8'd6,8'd64} : s = 268;
	{8'd6,8'd65} : s = 396;
	{8'd6,8'd66} : s = 68;
	{8'd6,8'd67} : s = 266;
	{8'd6,8'd68} : s = 265;
	{8'd6,8'd69} : s = 394;
	{8'd6,8'd70} : s = 262;
	{8'd6,8'd71} : s = 393;
	{8'd6,8'd72} : s = 390;
	{8'd6,8'd73} : s = 468;
	{8'd6,8'd74} : s = 66;
	{8'd6,8'd75} : s = 261;
	{8'd6,8'd76} : s = 259;
	{8'd6,8'd77} : s = 389;
	{8'd6,8'd78} : s = 224;
	{8'd6,8'd79} : s = 387;
	{8'd6,8'd80} : s = 368;
	{8'd6,8'd81} : s = 466;
	{8'd6,8'd82} : s = 208;
	{8'd6,8'd83} : s = 360;
	{8'd6,8'd84} : s = 356;
	{8'd6,8'd85} : s = 465;
	{8'd6,8'd86} : s = 354;
	{8'd6,8'd87} : s = 460;
	{8'd6,8'd88} : s = 458;
	{8'd6,8'd89} : s = 500;
	{8'd6,8'd90} : s = 65;
	{8'd6,8'd91} : s = 200;
	{8'd6,8'd92} : s = 196;
	{8'd6,8'd93} : s = 353;
	{8'd6,8'd94} : s = 194;
	{8'd6,8'd95} : s = 344;
	{8'd6,8'd96} : s = 340;
	{8'd6,8'd97} : s = 457;
	{8'd6,8'd98} : s = 193;
	{8'd6,8'd99} : s = 338;
	{8'd6,8'd100} : s = 337;
	{8'd6,8'd101} : s = 454;
	{8'd6,8'd102} : s = 332;
	{8'd6,8'd103} : s = 453;
	{8'd6,8'd104} : s = 451;
	{8'd6,8'd105} : s = 498;
	{8'd6,8'd106} : s = 176;
	{8'd6,8'd107} : s = 330;
	{8'd6,8'd108} : s = 329;
	{8'd6,8'd109} : s = 440;
	{8'd6,8'd110} : s = 326;
	{8'd6,8'd111} : s = 436;
	{8'd6,8'd112} : s = 434;
	{8'd6,8'd113} : s = 497;
	{8'd6,8'd114} : s = 325;
	{8'd6,8'd115} : s = 433;
	{8'd6,8'd116} : s = 428;
	{8'd6,8'd117} : s = 492;
	{8'd6,8'd118} : s = 426;
	{8'd6,8'd119} : s = 490;
	{8'd6,8'd120} : s = 489;
	{8'd6,8'd121} : s = 508;
	{8'd6,8'd122} : s = 2;
	{8'd6,8'd123} : s = 48;
	{8'd6,8'd124} : s = 40;
	{8'd6,8'd125} : s = 168;
	{8'd6,8'd126} : s = 36;
	{8'd6,8'd127} : s = 164;
	{8'd6,8'd128} : s = 162;
	{8'd6,8'd129} : s = 323;
	{8'd6,8'd130} : s = 34;
	{8'd6,8'd131} : s = 161;
	{8'd6,8'd132} : s = 152;
	{8'd6,8'd133} : s = 312;
	{8'd6,8'd134} : s = 148;
	{8'd6,8'd135} : s = 308;
	{8'd6,8'd136} : s = 306;
	{8'd6,8'd137} : s = 425;
	{8'd6,8'd138} : s = 33;
	{8'd6,8'd139} : s = 146;
	{8'd6,8'd140} : s = 145;
	{8'd6,8'd141} : s = 305;
	{8'd6,8'd142} : s = 140;
	{8'd6,8'd143} : s = 300;
	{8'd6,8'd144} : s = 298;
	{8'd6,8'd145} : s = 422;
	{8'd6,8'd146} : s = 138;
	{8'd6,8'd147} : s = 297;
	{8'd6,8'd148} : s = 294;
	{8'd6,8'd149} : s = 421;
	{8'd6,8'd150} : s = 293;
	{8'd6,8'd151} : s = 419;
	{8'd6,8'd152} : s = 412;
	{8'd6,8'd153} : s = 486;
	{8'd6,8'd154} : s = 24;
	{8'd6,8'd155} : s = 137;
	{8'd6,8'd156} : s = 134;
	{8'd6,8'd157} : s = 291;
	{8'd6,8'd158} : s = 133;
	{8'd6,8'd159} : s = 284;
	{8'd6,8'd160} : s = 282;
	{8'd6,8'd161} : s = 410;
	{8'd6,8'd162} : s = 131;
	{8'd6,8'd163} : s = 281;
	{8'd6,8'd164} : s = 278;
	{8'd6,8'd165} : s = 409;
	{8'd6,8'd166} : s = 277;
	{8'd6,8'd167} : s = 406;
	{8'd6,8'd168} : s = 405;
	{8'd6,8'd169} : s = 485;
	{8'd6,8'd170} : s = 112;
	{8'd6,8'd171} : s = 275;
	{8'd6,8'd172} : s = 270;
	{8'd6,8'd173} : s = 403;
	{8'd6,8'd174} : s = 269;
	{8'd6,8'd175} : s = 398;
	{8'd6,8'd176} : s = 397;
	{8'd6,8'd177} : s = 483;
	{8'd6,8'd178} : s = 267;
	{8'd6,8'd179} : s = 395;
	{8'd6,8'd180} : s = 391;
	{8'd6,8'd181} : s = 476;
	{8'd6,8'd182} : s = 376;
	{8'd6,8'd183} : s = 474;
	{8'd6,8'd184} : s = 473;
	{8'd6,8'd185} : s = 506;
	{8'd6,8'd186} : s = 20;
	{8'd6,8'd187} : s = 104;
	{8'd6,8'd188} : s = 100;
	{8'd6,8'd189} : s = 263;
	{8'd6,8'd190} : s = 98;
	{8'd6,8'd191} : s = 240;
	{8'd6,8'd192} : s = 232;
	{8'd6,8'd193} : s = 372;
	{8'd6,8'd194} : s = 97;
	{8'd6,8'd195} : s = 228;
	{8'd6,8'd196} : s = 226;
	{8'd6,8'd197} : s = 370;
	{8'd6,8'd198} : s = 225;
	{8'd6,8'd199} : s = 369;
	{8'd6,8'd200} : s = 364;
	{8'd6,8'd201} : s = 470;
	{8'd6,8'd202} : s = 88;
	{8'd6,8'd203} : s = 216;
	{8'd6,8'd204} : s = 212;
	{8'd6,8'd205} : s = 362;
	{8'd6,8'd206} : s = 210;
	{8'd6,8'd207} : s = 361;
	{8'd6,8'd208} : s = 358;
	{8'd6,8'd209} : s = 469;
	{8'd6,8'd210} : s = 209;
	{8'd6,8'd211} : s = 357;
	{8'd6,8'd212} : s = 355;
	{8'd6,8'd213} : s = 467;
	{8'd6,8'd214} : s = 348;
	{8'd6,8'd215} : s = 462;
	{8'd6,8'd216} : s = 461;
	{8'd6,8'd217} : s = 505;
	{8'd6,8'd218} : s = 84;
	{8'd6,8'd219} : s = 204;
	{8'd6,8'd220} : s = 202;
	{8'd6,8'd221} : s = 346;
	{8'd6,8'd222} : s = 201;
	{8'd6,8'd223} : s = 345;
	{8'd6,8'd224} : s = 342;
	{8'd6,8'd225} : s = 459;
	{8'd6,8'd226} : s = 198;
	{8'd6,8'd227} : s = 341;
	{8'd6,8'd228} : s = 339;
	{8'd6,8'd229} : s = 455;
	{8'd6,8'd230} : s = 334;
	{8'd6,8'd231} : s = 444;
	{8'd6,8'd232} : s = 442;
	{8'd6,8'd233} : s = 502;
	{8'd6,8'd234} : s = 197;
	{8'd6,8'd235} : s = 333;
	{8'd6,8'd236} : s = 331;
	{8'd6,8'd237} : s = 441;
	{8'd6,8'd238} : s = 327;
	{8'd6,8'd239} : s = 438;
	{8'd6,8'd240} : s = 437;
	{8'd6,8'd241} : s = 501;
	{8'd6,8'd242} : s = 316;
	{8'd6,8'd243} : s = 435;
	{8'd6,8'd244} : s = 430;
	{8'd6,8'd245} : s = 499;
	{8'd6,8'd246} : s = 429;
	{8'd6,8'd247} : s = 494;
	{8'd6,8'd248} : s = 493;
	{8'd6,8'd249} : s = 510;
	{8'd6,8'd250} : s = 1;
	{8'd6,8'd251} : s = 18;
	{8'd6,8'd252} : s = 17;
	{8'd6,8'd253} : s = 82;
	{8'd6,8'd254} : s = 12;
	{8'd6,8'd255} : s = 81;
	{8'd7,8'd0} : s = 448;
	{8'd7,8'd1} : s = 32;
	{8'd7,8'd2} : s = 272;
	{8'd7,8'd3} : s = 264;
	{8'd7,8'd4} : s = 416;
	{8'd7,8'd5} : s = 260;
	{8'd7,8'd6} : s = 400;
	{8'd7,8'd7} : s = 392;
	{8'd7,8'd8} : s = 480;
	{8'd7,8'd9} : s = 8;
	{8'd7,8'd10} : s = 258;
	{8'd7,8'd11} : s = 257;
	{8'd7,8'd12} : s = 388;
	{8'd7,8'd13} : s = 192;
	{8'd7,8'd14} : s = 386;
	{8'd7,8'd15} : s = 385;
	{8'd7,8'd16} : s = 464;
	{8'd7,8'd17} : s = 160;
	{8'd7,8'd18} : s = 352;
	{8'd7,8'd19} : s = 336;
	{8'd7,8'd20} : s = 456;
	{8'd7,8'd21} : s = 328;
	{8'd7,8'd22} : s = 452;
	{8'd7,8'd23} : s = 450;
	{8'd7,8'd24} : s = 496;
	{8'd7,8'd25} : s = 16;
	{8'd7,8'd26} : s = 144;
	{8'd7,8'd27} : s = 136;
	{8'd7,8'd28} : s = 324;
	{8'd7,8'd29} : s = 132;
	{8'd7,8'd30} : s = 322;
	{8'd7,8'd31} : s = 321;
	{8'd7,8'd32} : s = 449;
	{8'd7,8'd33} : s = 130;
	{8'd7,8'd34} : s = 304;
	{8'd7,8'd35} : s = 296;
	{8'd7,8'd36} : s = 432;
	{8'd7,8'd37} : s = 292;
	{8'd7,8'd38} : s = 424;
	{8'd7,8'd39} : s = 420;
	{8'd7,8'd40} : s = 488;
	{8'd7,8'd41} : s = 129;
	{8'd7,8'd42} : s = 290;
	{8'd7,8'd43} : s = 289;
	{8'd7,8'd44} : s = 418;
	{8'd7,8'd45} : s = 280;
	{8'd7,8'd46} : s = 417;
	{8'd7,8'd47} : s = 408;
	{8'd7,8'd48} : s = 484;
	{8'd7,8'd49} : s = 276;
	{8'd7,8'd50} : s = 404;
	{8'd7,8'd51} : s = 402;
	{8'd7,8'd52} : s = 482;
	{8'd7,8'd53} : s = 401;
	{8'd7,8'd54} : s = 481;
	{8'd7,8'd55} : s = 472;
	{8'd7,8'd56} : s = 504;
	{8'd7,8'd57} : s = 4;
	{8'd7,8'd58} : s = 96;
	{8'd7,8'd59} : s = 80;
	{8'd7,8'd60} : s = 274;
	{8'd7,8'd61} : s = 72;
	{8'd7,8'd62} : s = 273;
	{8'd7,8'd63} : s = 268;
	{8'd7,8'd64} : s = 396;
	{8'd7,8'd65} : s = 68;
	{8'd7,8'd66} : s = 266;
	{8'd7,8'd67} : s = 265;
	{8'd7,8'd68} : s = 394;
	{8'd7,8'd69} : s = 262;
	{8'd7,8'd70} : s = 393;
	{8'd7,8'd71} : s = 390;
	{8'd7,8'd72} : s = 468;
	{8'd7,8'd73} : s = 66;
	{8'd7,8'd74} : s = 261;
	{8'd7,8'd75} : s = 259;
	{8'd7,8'd76} : s = 389;
	{8'd7,8'd77} : s = 224;
	{8'd7,8'd78} : s = 387;
	{8'd7,8'd79} : s = 368;
	{8'd7,8'd80} : s = 466;
	{8'd7,8'd81} : s = 208;
	{8'd7,8'd82} : s = 360;
	{8'd7,8'd83} : s = 356;
	{8'd7,8'd84} : s = 465;
	{8'd7,8'd85} : s = 354;
	{8'd7,8'd86} : s = 460;
	{8'd7,8'd87} : s = 458;
	{8'd7,8'd88} : s = 500;
	{8'd7,8'd89} : s = 65;
	{8'd7,8'd90} : s = 200;
	{8'd7,8'd91} : s = 196;
	{8'd7,8'd92} : s = 353;
	{8'd7,8'd93} : s = 194;
	{8'd7,8'd94} : s = 344;
	{8'd7,8'd95} : s = 340;
	{8'd7,8'd96} : s = 457;
	{8'd7,8'd97} : s = 193;
	{8'd7,8'd98} : s = 338;
	{8'd7,8'd99} : s = 337;
	{8'd7,8'd100} : s = 454;
	{8'd7,8'd101} : s = 332;
	{8'd7,8'd102} : s = 453;
	{8'd7,8'd103} : s = 451;
	{8'd7,8'd104} : s = 498;
	{8'd7,8'd105} : s = 176;
	{8'd7,8'd106} : s = 330;
	{8'd7,8'd107} : s = 329;
	{8'd7,8'd108} : s = 440;
	{8'd7,8'd109} : s = 326;
	{8'd7,8'd110} : s = 436;
	{8'd7,8'd111} : s = 434;
	{8'd7,8'd112} : s = 497;
	{8'd7,8'd113} : s = 325;
	{8'd7,8'd114} : s = 433;
	{8'd7,8'd115} : s = 428;
	{8'd7,8'd116} : s = 492;
	{8'd7,8'd117} : s = 426;
	{8'd7,8'd118} : s = 490;
	{8'd7,8'd119} : s = 489;
	{8'd7,8'd120} : s = 508;
	{8'd7,8'd121} : s = 2;
	{8'd7,8'd122} : s = 48;
	{8'd7,8'd123} : s = 40;
	{8'd7,8'd124} : s = 168;
	{8'd7,8'd125} : s = 36;
	{8'd7,8'd126} : s = 164;
	{8'd7,8'd127} : s = 162;
	{8'd7,8'd128} : s = 323;
	{8'd7,8'd129} : s = 34;
	{8'd7,8'd130} : s = 161;
	{8'd7,8'd131} : s = 152;
	{8'd7,8'd132} : s = 312;
	{8'd7,8'd133} : s = 148;
	{8'd7,8'd134} : s = 308;
	{8'd7,8'd135} : s = 306;
	{8'd7,8'd136} : s = 425;
	{8'd7,8'd137} : s = 33;
	{8'd7,8'd138} : s = 146;
	{8'd7,8'd139} : s = 145;
	{8'd7,8'd140} : s = 305;
	{8'd7,8'd141} : s = 140;
	{8'd7,8'd142} : s = 300;
	{8'd7,8'd143} : s = 298;
	{8'd7,8'd144} : s = 422;
	{8'd7,8'd145} : s = 138;
	{8'd7,8'd146} : s = 297;
	{8'd7,8'd147} : s = 294;
	{8'd7,8'd148} : s = 421;
	{8'd7,8'd149} : s = 293;
	{8'd7,8'd150} : s = 419;
	{8'd7,8'd151} : s = 412;
	{8'd7,8'd152} : s = 486;
	{8'd7,8'd153} : s = 24;
	{8'd7,8'd154} : s = 137;
	{8'd7,8'd155} : s = 134;
	{8'd7,8'd156} : s = 291;
	{8'd7,8'd157} : s = 133;
	{8'd7,8'd158} : s = 284;
	{8'd7,8'd159} : s = 282;
	{8'd7,8'd160} : s = 410;
	{8'd7,8'd161} : s = 131;
	{8'd7,8'd162} : s = 281;
	{8'd7,8'd163} : s = 278;
	{8'd7,8'd164} : s = 409;
	{8'd7,8'd165} : s = 277;
	{8'd7,8'd166} : s = 406;
	{8'd7,8'd167} : s = 405;
	{8'd7,8'd168} : s = 485;
	{8'd7,8'd169} : s = 112;
	{8'd7,8'd170} : s = 275;
	{8'd7,8'd171} : s = 270;
	{8'd7,8'd172} : s = 403;
	{8'd7,8'd173} : s = 269;
	{8'd7,8'd174} : s = 398;
	{8'd7,8'd175} : s = 397;
	{8'd7,8'd176} : s = 483;
	{8'd7,8'd177} : s = 267;
	{8'd7,8'd178} : s = 395;
	{8'd7,8'd179} : s = 391;
	{8'd7,8'd180} : s = 476;
	{8'd7,8'd181} : s = 376;
	{8'd7,8'd182} : s = 474;
	{8'd7,8'd183} : s = 473;
	{8'd7,8'd184} : s = 506;
	{8'd7,8'd185} : s = 20;
	{8'd7,8'd186} : s = 104;
	{8'd7,8'd187} : s = 100;
	{8'd7,8'd188} : s = 263;
	{8'd7,8'd189} : s = 98;
	{8'd7,8'd190} : s = 240;
	{8'd7,8'd191} : s = 232;
	{8'd7,8'd192} : s = 372;
	{8'd7,8'd193} : s = 97;
	{8'd7,8'd194} : s = 228;
	{8'd7,8'd195} : s = 226;
	{8'd7,8'd196} : s = 370;
	{8'd7,8'd197} : s = 225;
	{8'd7,8'd198} : s = 369;
	{8'd7,8'd199} : s = 364;
	{8'd7,8'd200} : s = 470;
	{8'd7,8'd201} : s = 88;
	{8'd7,8'd202} : s = 216;
	{8'd7,8'd203} : s = 212;
	{8'd7,8'd204} : s = 362;
	{8'd7,8'd205} : s = 210;
	{8'd7,8'd206} : s = 361;
	{8'd7,8'd207} : s = 358;
	{8'd7,8'd208} : s = 469;
	{8'd7,8'd209} : s = 209;
	{8'd7,8'd210} : s = 357;
	{8'd7,8'd211} : s = 355;
	{8'd7,8'd212} : s = 467;
	{8'd7,8'd213} : s = 348;
	{8'd7,8'd214} : s = 462;
	{8'd7,8'd215} : s = 461;
	{8'd7,8'd216} : s = 505;
	{8'd7,8'd217} : s = 84;
	{8'd7,8'd218} : s = 204;
	{8'd7,8'd219} : s = 202;
	{8'd7,8'd220} : s = 346;
	{8'd7,8'd221} : s = 201;
	{8'd7,8'd222} : s = 345;
	{8'd7,8'd223} : s = 342;
	{8'd7,8'd224} : s = 459;
	{8'd7,8'd225} : s = 198;
	{8'd7,8'd226} : s = 341;
	{8'd7,8'd227} : s = 339;
	{8'd7,8'd228} : s = 455;
	{8'd7,8'd229} : s = 334;
	{8'd7,8'd230} : s = 444;
	{8'd7,8'd231} : s = 442;
	{8'd7,8'd232} : s = 502;
	{8'd7,8'd233} : s = 197;
	{8'd7,8'd234} : s = 333;
	{8'd7,8'd235} : s = 331;
	{8'd7,8'd236} : s = 441;
	{8'd7,8'd237} : s = 327;
	{8'd7,8'd238} : s = 438;
	{8'd7,8'd239} : s = 437;
	{8'd7,8'd240} : s = 501;
	{8'd7,8'd241} : s = 316;
	{8'd7,8'd242} : s = 435;
	{8'd7,8'd243} : s = 430;
	{8'd7,8'd244} : s = 499;
	{8'd7,8'd245} : s = 429;
	{8'd7,8'd246} : s = 494;
	{8'd7,8'd247} : s = 493;
	{8'd7,8'd248} : s = 510;
	{8'd7,8'd249} : s = 1;
	{8'd7,8'd250} : s = 18;
	{8'd7,8'd251} : s = 17;
	{8'd7,8'd252} : s = 82;
	{8'd7,8'd253} : s = 12;
	{8'd7,8'd254} : s = 81;
	{8'd7,8'd255} : s = 76;
	{8'd8,8'd0} : s = 32;
	{8'd8,8'd1} : s = 272;
	{8'd8,8'd2} : s = 264;
	{8'd8,8'd3} : s = 416;
	{8'd8,8'd4} : s = 260;
	{8'd8,8'd5} : s = 400;
	{8'd8,8'd6} : s = 392;
	{8'd8,8'd7} : s = 480;
	{8'd8,8'd8} : s = 8;
	{8'd8,8'd9} : s = 258;
	{8'd8,8'd10} : s = 257;
	{8'd8,8'd11} : s = 388;
	{8'd8,8'd12} : s = 192;
	{8'd8,8'd13} : s = 386;
	{8'd8,8'd14} : s = 385;
	{8'd8,8'd15} : s = 464;
	{8'd8,8'd16} : s = 160;
	{8'd8,8'd17} : s = 352;
	{8'd8,8'd18} : s = 336;
	{8'd8,8'd19} : s = 456;
	{8'd8,8'd20} : s = 328;
	{8'd8,8'd21} : s = 452;
	{8'd8,8'd22} : s = 450;
	{8'd8,8'd23} : s = 496;
	{8'd8,8'd24} : s = 16;
	{8'd8,8'd25} : s = 144;
	{8'd8,8'd26} : s = 136;
	{8'd8,8'd27} : s = 324;
	{8'd8,8'd28} : s = 132;
	{8'd8,8'd29} : s = 322;
	{8'd8,8'd30} : s = 321;
	{8'd8,8'd31} : s = 449;
	{8'd8,8'd32} : s = 130;
	{8'd8,8'd33} : s = 304;
	{8'd8,8'd34} : s = 296;
	{8'd8,8'd35} : s = 432;
	{8'd8,8'd36} : s = 292;
	{8'd8,8'd37} : s = 424;
	{8'd8,8'd38} : s = 420;
	{8'd8,8'd39} : s = 488;
	{8'd8,8'd40} : s = 129;
	{8'd8,8'd41} : s = 290;
	{8'd8,8'd42} : s = 289;
	{8'd8,8'd43} : s = 418;
	{8'd8,8'd44} : s = 280;
	{8'd8,8'd45} : s = 417;
	{8'd8,8'd46} : s = 408;
	{8'd8,8'd47} : s = 484;
	{8'd8,8'd48} : s = 276;
	{8'd8,8'd49} : s = 404;
	{8'd8,8'd50} : s = 402;
	{8'd8,8'd51} : s = 482;
	{8'd8,8'd52} : s = 401;
	{8'd8,8'd53} : s = 481;
	{8'd8,8'd54} : s = 472;
	{8'd8,8'd55} : s = 504;
	{8'd8,8'd56} : s = 4;
	{8'd8,8'd57} : s = 96;
	{8'd8,8'd58} : s = 80;
	{8'd8,8'd59} : s = 274;
	{8'd8,8'd60} : s = 72;
	{8'd8,8'd61} : s = 273;
	{8'd8,8'd62} : s = 268;
	{8'd8,8'd63} : s = 396;
	{8'd8,8'd64} : s = 68;
	{8'd8,8'd65} : s = 266;
	{8'd8,8'd66} : s = 265;
	{8'd8,8'd67} : s = 394;
	{8'd8,8'd68} : s = 262;
	{8'd8,8'd69} : s = 393;
	{8'd8,8'd70} : s = 390;
	{8'd8,8'd71} : s = 468;
	{8'd8,8'd72} : s = 66;
	{8'd8,8'd73} : s = 261;
	{8'd8,8'd74} : s = 259;
	{8'd8,8'd75} : s = 389;
	{8'd8,8'd76} : s = 224;
	{8'd8,8'd77} : s = 387;
	{8'd8,8'd78} : s = 368;
	{8'd8,8'd79} : s = 466;
	{8'd8,8'd80} : s = 208;
	{8'd8,8'd81} : s = 360;
	{8'd8,8'd82} : s = 356;
	{8'd8,8'd83} : s = 465;
	{8'd8,8'd84} : s = 354;
	{8'd8,8'd85} : s = 460;
	{8'd8,8'd86} : s = 458;
	{8'd8,8'd87} : s = 500;
	{8'd8,8'd88} : s = 65;
	{8'd8,8'd89} : s = 200;
	{8'd8,8'd90} : s = 196;
	{8'd8,8'd91} : s = 353;
	{8'd8,8'd92} : s = 194;
	{8'd8,8'd93} : s = 344;
	{8'd8,8'd94} : s = 340;
	{8'd8,8'd95} : s = 457;
	{8'd8,8'd96} : s = 193;
	{8'd8,8'd97} : s = 338;
	{8'd8,8'd98} : s = 337;
	{8'd8,8'd99} : s = 454;
	{8'd8,8'd100} : s = 332;
	{8'd8,8'd101} : s = 453;
	{8'd8,8'd102} : s = 451;
	{8'd8,8'd103} : s = 498;
	{8'd8,8'd104} : s = 176;
	{8'd8,8'd105} : s = 330;
	{8'd8,8'd106} : s = 329;
	{8'd8,8'd107} : s = 440;
	{8'd8,8'd108} : s = 326;
	{8'd8,8'd109} : s = 436;
	{8'd8,8'd110} : s = 434;
	{8'd8,8'd111} : s = 497;
	{8'd8,8'd112} : s = 325;
	{8'd8,8'd113} : s = 433;
	{8'd8,8'd114} : s = 428;
	{8'd8,8'd115} : s = 492;
	{8'd8,8'd116} : s = 426;
	{8'd8,8'd117} : s = 490;
	{8'd8,8'd118} : s = 489;
	{8'd8,8'd119} : s = 508;
	{8'd8,8'd120} : s = 2;
	{8'd8,8'd121} : s = 48;
	{8'd8,8'd122} : s = 40;
	{8'd8,8'd123} : s = 168;
	{8'd8,8'd124} : s = 36;
	{8'd8,8'd125} : s = 164;
	{8'd8,8'd126} : s = 162;
	{8'd8,8'd127} : s = 323;
	{8'd8,8'd128} : s = 34;
	{8'd8,8'd129} : s = 161;
	{8'd8,8'd130} : s = 152;
	{8'd8,8'd131} : s = 312;
	{8'd8,8'd132} : s = 148;
	{8'd8,8'd133} : s = 308;
	{8'd8,8'd134} : s = 306;
	{8'd8,8'd135} : s = 425;
	{8'd8,8'd136} : s = 33;
	{8'd8,8'd137} : s = 146;
	{8'd8,8'd138} : s = 145;
	{8'd8,8'd139} : s = 305;
	{8'd8,8'd140} : s = 140;
	{8'd8,8'd141} : s = 300;
	{8'd8,8'd142} : s = 298;
	{8'd8,8'd143} : s = 422;
	{8'd8,8'd144} : s = 138;
	{8'd8,8'd145} : s = 297;
	{8'd8,8'd146} : s = 294;
	{8'd8,8'd147} : s = 421;
	{8'd8,8'd148} : s = 293;
	{8'd8,8'd149} : s = 419;
	{8'd8,8'd150} : s = 412;
	{8'd8,8'd151} : s = 486;
	{8'd8,8'd152} : s = 24;
	{8'd8,8'd153} : s = 137;
	{8'd8,8'd154} : s = 134;
	{8'd8,8'd155} : s = 291;
	{8'd8,8'd156} : s = 133;
	{8'd8,8'd157} : s = 284;
	{8'd8,8'd158} : s = 282;
	{8'd8,8'd159} : s = 410;
	{8'd8,8'd160} : s = 131;
	{8'd8,8'd161} : s = 281;
	{8'd8,8'd162} : s = 278;
	{8'd8,8'd163} : s = 409;
	{8'd8,8'd164} : s = 277;
	{8'd8,8'd165} : s = 406;
	{8'd8,8'd166} : s = 405;
	{8'd8,8'd167} : s = 485;
	{8'd8,8'd168} : s = 112;
	{8'd8,8'd169} : s = 275;
	{8'd8,8'd170} : s = 270;
	{8'd8,8'd171} : s = 403;
	{8'd8,8'd172} : s = 269;
	{8'd8,8'd173} : s = 398;
	{8'd8,8'd174} : s = 397;
	{8'd8,8'd175} : s = 483;
	{8'd8,8'd176} : s = 267;
	{8'd8,8'd177} : s = 395;
	{8'd8,8'd178} : s = 391;
	{8'd8,8'd179} : s = 476;
	{8'd8,8'd180} : s = 376;
	{8'd8,8'd181} : s = 474;
	{8'd8,8'd182} : s = 473;
	{8'd8,8'd183} : s = 506;
	{8'd8,8'd184} : s = 20;
	{8'd8,8'd185} : s = 104;
	{8'd8,8'd186} : s = 100;
	{8'd8,8'd187} : s = 263;
	{8'd8,8'd188} : s = 98;
	{8'd8,8'd189} : s = 240;
	{8'd8,8'd190} : s = 232;
	{8'd8,8'd191} : s = 372;
	{8'd8,8'd192} : s = 97;
	{8'd8,8'd193} : s = 228;
	{8'd8,8'd194} : s = 226;
	{8'd8,8'd195} : s = 370;
	{8'd8,8'd196} : s = 225;
	{8'd8,8'd197} : s = 369;
	{8'd8,8'd198} : s = 364;
	{8'd8,8'd199} : s = 470;
	{8'd8,8'd200} : s = 88;
	{8'd8,8'd201} : s = 216;
	{8'd8,8'd202} : s = 212;
	{8'd8,8'd203} : s = 362;
	{8'd8,8'd204} : s = 210;
	{8'd8,8'd205} : s = 361;
	{8'd8,8'd206} : s = 358;
	{8'd8,8'd207} : s = 469;
	{8'd8,8'd208} : s = 209;
	{8'd8,8'd209} : s = 357;
	{8'd8,8'd210} : s = 355;
	{8'd8,8'd211} : s = 467;
	{8'd8,8'd212} : s = 348;
	{8'd8,8'd213} : s = 462;
	{8'd8,8'd214} : s = 461;
	{8'd8,8'd215} : s = 505;
	{8'd8,8'd216} : s = 84;
	{8'd8,8'd217} : s = 204;
	{8'd8,8'd218} : s = 202;
	{8'd8,8'd219} : s = 346;
	{8'd8,8'd220} : s = 201;
	{8'd8,8'd221} : s = 345;
	{8'd8,8'd222} : s = 342;
	{8'd8,8'd223} : s = 459;
	{8'd8,8'd224} : s = 198;
	{8'd8,8'd225} : s = 341;
	{8'd8,8'd226} : s = 339;
	{8'd8,8'd227} : s = 455;
	{8'd8,8'd228} : s = 334;
	{8'd8,8'd229} : s = 444;
	{8'd8,8'd230} : s = 442;
	{8'd8,8'd231} : s = 502;
	{8'd8,8'd232} : s = 197;
	{8'd8,8'd233} : s = 333;
	{8'd8,8'd234} : s = 331;
	{8'd8,8'd235} : s = 441;
	{8'd8,8'd236} : s = 327;
	{8'd8,8'd237} : s = 438;
	{8'd8,8'd238} : s = 437;
	{8'd8,8'd239} : s = 501;
	{8'd8,8'd240} : s = 316;
	{8'd8,8'd241} : s = 435;
	{8'd8,8'd242} : s = 430;
	{8'd8,8'd243} : s = 499;
	{8'd8,8'd244} : s = 429;
	{8'd8,8'd245} : s = 494;
	{8'd8,8'd246} : s = 493;
	{8'd8,8'd247} : s = 510;
	{8'd8,8'd248} : s = 1;
	{8'd8,8'd249} : s = 18;
	{8'd8,8'd250} : s = 17;
	{8'd8,8'd251} : s = 82;
	{8'd8,8'd252} : s = 12;
	{8'd8,8'd253} : s = 81;
	{8'd8,8'd254} : s = 76;
	{8'd8,8'd255} : s = 195;
	{8'd9,8'd0} : s = 272;
	{8'd9,8'd1} : s = 264;
	{8'd9,8'd2} : s = 416;
	{8'd9,8'd3} : s = 260;
	{8'd9,8'd4} : s = 400;
	{8'd9,8'd5} : s = 392;
	{8'd9,8'd6} : s = 480;
	{8'd9,8'd7} : s = 8;
	{8'd9,8'd8} : s = 258;
	{8'd9,8'd9} : s = 257;
	{8'd9,8'd10} : s = 388;
	{8'd9,8'd11} : s = 192;
	{8'd9,8'd12} : s = 386;
	{8'd9,8'd13} : s = 385;
	{8'd9,8'd14} : s = 464;
	{8'd9,8'd15} : s = 160;
	{8'd9,8'd16} : s = 352;
	{8'd9,8'd17} : s = 336;
	{8'd9,8'd18} : s = 456;
	{8'd9,8'd19} : s = 328;
	{8'd9,8'd20} : s = 452;
	{8'd9,8'd21} : s = 450;
	{8'd9,8'd22} : s = 496;
	{8'd9,8'd23} : s = 16;
	{8'd9,8'd24} : s = 144;
	{8'd9,8'd25} : s = 136;
	{8'd9,8'd26} : s = 324;
	{8'd9,8'd27} : s = 132;
	{8'd9,8'd28} : s = 322;
	{8'd9,8'd29} : s = 321;
	{8'd9,8'd30} : s = 449;
	{8'd9,8'd31} : s = 130;
	{8'd9,8'd32} : s = 304;
	{8'd9,8'd33} : s = 296;
	{8'd9,8'd34} : s = 432;
	{8'd9,8'd35} : s = 292;
	{8'd9,8'd36} : s = 424;
	{8'd9,8'd37} : s = 420;
	{8'd9,8'd38} : s = 488;
	{8'd9,8'd39} : s = 129;
	{8'd9,8'd40} : s = 290;
	{8'd9,8'd41} : s = 289;
	{8'd9,8'd42} : s = 418;
	{8'd9,8'd43} : s = 280;
	{8'd9,8'd44} : s = 417;
	{8'd9,8'd45} : s = 408;
	{8'd9,8'd46} : s = 484;
	{8'd9,8'd47} : s = 276;
	{8'd9,8'd48} : s = 404;
	{8'd9,8'd49} : s = 402;
	{8'd9,8'd50} : s = 482;
	{8'd9,8'd51} : s = 401;
	{8'd9,8'd52} : s = 481;
	{8'd9,8'd53} : s = 472;
	{8'd9,8'd54} : s = 504;
	{8'd9,8'd55} : s = 4;
	{8'd9,8'd56} : s = 96;
	{8'd9,8'd57} : s = 80;
	{8'd9,8'd58} : s = 274;
	{8'd9,8'd59} : s = 72;
	{8'd9,8'd60} : s = 273;
	{8'd9,8'd61} : s = 268;
	{8'd9,8'd62} : s = 396;
	{8'd9,8'd63} : s = 68;
	{8'd9,8'd64} : s = 266;
	{8'd9,8'd65} : s = 265;
	{8'd9,8'd66} : s = 394;
	{8'd9,8'd67} : s = 262;
	{8'd9,8'd68} : s = 393;
	{8'd9,8'd69} : s = 390;
	{8'd9,8'd70} : s = 468;
	{8'd9,8'd71} : s = 66;
	{8'd9,8'd72} : s = 261;
	{8'd9,8'd73} : s = 259;
	{8'd9,8'd74} : s = 389;
	{8'd9,8'd75} : s = 224;
	{8'd9,8'd76} : s = 387;
	{8'd9,8'd77} : s = 368;
	{8'd9,8'd78} : s = 466;
	{8'd9,8'd79} : s = 208;
	{8'd9,8'd80} : s = 360;
	{8'd9,8'd81} : s = 356;
	{8'd9,8'd82} : s = 465;
	{8'd9,8'd83} : s = 354;
	{8'd9,8'd84} : s = 460;
	{8'd9,8'd85} : s = 458;
	{8'd9,8'd86} : s = 500;
	{8'd9,8'd87} : s = 65;
	{8'd9,8'd88} : s = 200;
	{8'd9,8'd89} : s = 196;
	{8'd9,8'd90} : s = 353;
	{8'd9,8'd91} : s = 194;
	{8'd9,8'd92} : s = 344;
	{8'd9,8'd93} : s = 340;
	{8'd9,8'd94} : s = 457;
	{8'd9,8'd95} : s = 193;
	{8'd9,8'd96} : s = 338;
	{8'd9,8'd97} : s = 337;
	{8'd9,8'd98} : s = 454;
	{8'd9,8'd99} : s = 332;
	{8'd9,8'd100} : s = 453;
	{8'd9,8'd101} : s = 451;
	{8'd9,8'd102} : s = 498;
	{8'd9,8'd103} : s = 176;
	{8'd9,8'd104} : s = 330;
	{8'd9,8'd105} : s = 329;
	{8'd9,8'd106} : s = 440;
	{8'd9,8'd107} : s = 326;
	{8'd9,8'd108} : s = 436;
	{8'd9,8'd109} : s = 434;
	{8'd9,8'd110} : s = 497;
	{8'd9,8'd111} : s = 325;
	{8'd9,8'd112} : s = 433;
	{8'd9,8'd113} : s = 428;
	{8'd9,8'd114} : s = 492;
	{8'd9,8'd115} : s = 426;
	{8'd9,8'd116} : s = 490;
	{8'd9,8'd117} : s = 489;
	{8'd9,8'd118} : s = 508;
	{8'd9,8'd119} : s = 2;
	{8'd9,8'd120} : s = 48;
	{8'd9,8'd121} : s = 40;
	{8'd9,8'd122} : s = 168;
	{8'd9,8'd123} : s = 36;
	{8'd9,8'd124} : s = 164;
	{8'd9,8'd125} : s = 162;
	{8'd9,8'd126} : s = 323;
	{8'd9,8'd127} : s = 34;
	{8'd9,8'd128} : s = 161;
	{8'd9,8'd129} : s = 152;
	{8'd9,8'd130} : s = 312;
	{8'd9,8'd131} : s = 148;
	{8'd9,8'd132} : s = 308;
	{8'd9,8'd133} : s = 306;
	{8'd9,8'd134} : s = 425;
	{8'd9,8'd135} : s = 33;
	{8'd9,8'd136} : s = 146;
	{8'd9,8'd137} : s = 145;
	{8'd9,8'd138} : s = 305;
	{8'd9,8'd139} : s = 140;
	{8'd9,8'd140} : s = 300;
	{8'd9,8'd141} : s = 298;
	{8'd9,8'd142} : s = 422;
	{8'd9,8'd143} : s = 138;
	{8'd9,8'd144} : s = 297;
	{8'd9,8'd145} : s = 294;
	{8'd9,8'd146} : s = 421;
	{8'd9,8'd147} : s = 293;
	{8'd9,8'd148} : s = 419;
	{8'd9,8'd149} : s = 412;
	{8'd9,8'd150} : s = 486;
	{8'd9,8'd151} : s = 24;
	{8'd9,8'd152} : s = 137;
	{8'd9,8'd153} : s = 134;
	{8'd9,8'd154} : s = 291;
	{8'd9,8'd155} : s = 133;
	{8'd9,8'd156} : s = 284;
	{8'd9,8'd157} : s = 282;
	{8'd9,8'd158} : s = 410;
	{8'd9,8'd159} : s = 131;
	{8'd9,8'd160} : s = 281;
	{8'd9,8'd161} : s = 278;
	{8'd9,8'd162} : s = 409;
	{8'd9,8'd163} : s = 277;
	{8'd9,8'd164} : s = 406;
	{8'd9,8'd165} : s = 405;
	{8'd9,8'd166} : s = 485;
	{8'd9,8'd167} : s = 112;
	{8'd9,8'd168} : s = 275;
	{8'd9,8'd169} : s = 270;
	{8'd9,8'd170} : s = 403;
	{8'd9,8'd171} : s = 269;
	{8'd9,8'd172} : s = 398;
	{8'd9,8'd173} : s = 397;
	{8'd9,8'd174} : s = 483;
	{8'd9,8'd175} : s = 267;
	{8'd9,8'd176} : s = 395;
	{8'd9,8'd177} : s = 391;
	{8'd9,8'd178} : s = 476;
	{8'd9,8'd179} : s = 376;
	{8'd9,8'd180} : s = 474;
	{8'd9,8'd181} : s = 473;
	{8'd9,8'd182} : s = 506;
	{8'd9,8'd183} : s = 20;
	{8'd9,8'd184} : s = 104;
	{8'd9,8'd185} : s = 100;
	{8'd9,8'd186} : s = 263;
	{8'd9,8'd187} : s = 98;
	{8'd9,8'd188} : s = 240;
	{8'd9,8'd189} : s = 232;
	{8'd9,8'd190} : s = 372;
	{8'd9,8'd191} : s = 97;
	{8'd9,8'd192} : s = 228;
	{8'd9,8'd193} : s = 226;
	{8'd9,8'd194} : s = 370;
	{8'd9,8'd195} : s = 225;
	{8'd9,8'd196} : s = 369;
	{8'd9,8'd197} : s = 364;
	{8'd9,8'd198} : s = 470;
	{8'd9,8'd199} : s = 88;
	{8'd9,8'd200} : s = 216;
	{8'd9,8'd201} : s = 212;
	{8'd9,8'd202} : s = 362;
	{8'd9,8'd203} : s = 210;
	{8'd9,8'd204} : s = 361;
	{8'd9,8'd205} : s = 358;
	{8'd9,8'd206} : s = 469;
	{8'd9,8'd207} : s = 209;
	{8'd9,8'd208} : s = 357;
	{8'd9,8'd209} : s = 355;
	{8'd9,8'd210} : s = 467;
	{8'd9,8'd211} : s = 348;
	{8'd9,8'd212} : s = 462;
	{8'd9,8'd213} : s = 461;
	{8'd9,8'd214} : s = 505;
	{8'd9,8'd215} : s = 84;
	{8'd9,8'd216} : s = 204;
	{8'd9,8'd217} : s = 202;
	{8'd9,8'd218} : s = 346;
	{8'd9,8'd219} : s = 201;
	{8'd9,8'd220} : s = 345;
	{8'd9,8'd221} : s = 342;
	{8'd9,8'd222} : s = 459;
	{8'd9,8'd223} : s = 198;
	{8'd9,8'd224} : s = 341;
	{8'd9,8'd225} : s = 339;
	{8'd9,8'd226} : s = 455;
	{8'd9,8'd227} : s = 334;
	{8'd9,8'd228} : s = 444;
	{8'd9,8'd229} : s = 442;
	{8'd9,8'd230} : s = 502;
	{8'd9,8'd231} : s = 197;
	{8'd9,8'd232} : s = 333;
	{8'd9,8'd233} : s = 331;
	{8'd9,8'd234} : s = 441;
	{8'd9,8'd235} : s = 327;
	{8'd9,8'd236} : s = 438;
	{8'd9,8'd237} : s = 437;
	{8'd9,8'd238} : s = 501;
	{8'd9,8'd239} : s = 316;
	{8'd9,8'd240} : s = 435;
	{8'd9,8'd241} : s = 430;
	{8'd9,8'd242} : s = 499;
	{8'd9,8'd243} : s = 429;
	{8'd9,8'd244} : s = 494;
	{8'd9,8'd245} : s = 493;
	{8'd9,8'd246} : s = 510;
	{8'd9,8'd247} : s = 1;
	{8'd9,8'd248} : s = 18;
	{8'd9,8'd249} : s = 17;
	{8'd9,8'd250} : s = 82;
	{8'd9,8'd251} : s = 12;
	{8'd9,8'd252} : s = 81;
	{8'd9,8'd253} : s = 76;
	{8'd9,8'd254} : s = 195;
	{8'd9,8'd255} : s = 10;
	{8'd10,8'd0} : s = 264;
	{8'd10,8'd1} : s = 416;
	{8'd10,8'd2} : s = 260;
	{8'd10,8'd3} : s = 400;
	{8'd10,8'd4} : s = 392;
	{8'd10,8'd5} : s = 480;
	{8'd10,8'd6} : s = 8;
	{8'd10,8'd7} : s = 258;
	{8'd10,8'd8} : s = 257;
	{8'd10,8'd9} : s = 388;
	{8'd10,8'd10} : s = 192;
	{8'd10,8'd11} : s = 386;
	{8'd10,8'd12} : s = 385;
	{8'd10,8'd13} : s = 464;
	{8'd10,8'd14} : s = 160;
	{8'd10,8'd15} : s = 352;
	{8'd10,8'd16} : s = 336;
	{8'd10,8'd17} : s = 456;
	{8'd10,8'd18} : s = 328;
	{8'd10,8'd19} : s = 452;
	{8'd10,8'd20} : s = 450;
	{8'd10,8'd21} : s = 496;
	{8'd10,8'd22} : s = 16;
	{8'd10,8'd23} : s = 144;
	{8'd10,8'd24} : s = 136;
	{8'd10,8'd25} : s = 324;
	{8'd10,8'd26} : s = 132;
	{8'd10,8'd27} : s = 322;
	{8'd10,8'd28} : s = 321;
	{8'd10,8'd29} : s = 449;
	{8'd10,8'd30} : s = 130;
	{8'd10,8'd31} : s = 304;
	{8'd10,8'd32} : s = 296;
	{8'd10,8'd33} : s = 432;
	{8'd10,8'd34} : s = 292;
	{8'd10,8'd35} : s = 424;
	{8'd10,8'd36} : s = 420;
	{8'd10,8'd37} : s = 488;
	{8'd10,8'd38} : s = 129;
	{8'd10,8'd39} : s = 290;
	{8'd10,8'd40} : s = 289;
	{8'd10,8'd41} : s = 418;
	{8'd10,8'd42} : s = 280;
	{8'd10,8'd43} : s = 417;
	{8'd10,8'd44} : s = 408;
	{8'd10,8'd45} : s = 484;
	{8'd10,8'd46} : s = 276;
	{8'd10,8'd47} : s = 404;
	{8'd10,8'd48} : s = 402;
	{8'd10,8'd49} : s = 482;
	{8'd10,8'd50} : s = 401;
	{8'd10,8'd51} : s = 481;
	{8'd10,8'd52} : s = 472;
	{8'd10,8'd53} : s = 504;
	{8'd10,8'd54} : s = 4;
	{8'd10,8'd55} : s = 96;
	{8'd10,8'd56} : s = 80;
	{8'd10,8'd57} : s = 274;
	{8'd10,8'd58} : s = 72;
	{8'd10,8'd59} : s = 273;
	{8'd10,8'd60} : s = 268;
	{8'd10,8'd61} : s = 396;
	{8'd10,8'd62} : s = 68;
	{8'd10,8'd63} : s = 266;
	{8'd10,8'd64} : s = 265;
	{8'd10,8'd65} : s = 394;
	{8'd10,8'd66} : s = 262;
	{8'd10,8'd67} : s = 393;
	{8'd10,8'd68} : s = 390;
	{8'd10,8'd69} : s = 468;
	{8'd10,8'd70} : s = 66;
	{8'd10,8'd71} : s = 261;
	{8'd10,8'd72} : s = 259;
	{8'd10,8'd73} : s = 389;
	{8'd10,8'd74} : s = 224;
	{8'd10,8'd75} : s = 387;
	{8'd10,8'd76} : s = 368;
	{8'd10,8'd77} : s = 466;
	{8'd10,8'd78} : s = 208;
	{8'd10,8'd79} : s = 360;
	{8'd10,8'd80} : s = 356;
	{8'd10,8'd81} : s = 465;
	{8'd10,8'd82} : s = 354;
	{8'd10,8'd83} : s = 460;
	{8'd10,8'd84} : s = 458;
	{8'd10,8'd85} : s = 500;
	{8'd10,8'd86} : s = 65;
	{8'd10,8'd87} : s = 200;
	{8'd10,8'd88} : s = 196;
	{8'd10,8'd89} : s = 353;
	{8'd10,8'd90} : s = 194;
	{8'd10,8'd91} : s = 344;
	{8'd10,8'd92} : s = 340;
	{8'd10,8'd93} : s = 457;
	{8'd10,8'd94} : s = 193;
	{8'd10,8'd95} : s = 338;
	{8'd10,8'd96} : s = 337;
	{8'd10,8'd97} : s = 454;
	{8'd10,8'd98} : s = 332;
	{8'd10,8'd99} : s = 453;
	{8'd10,8'd100} : s = 451;
	{8'd10,8'd101} : s = 498;
	{8'd10,8'd102} : s = 176;
	{8'd10,8'd103} : s = 330;
	{8'd10,8'd104} : s = 329;
	{8'd10,8'd105} : s = 440;
	{8'd10,8'd106} : s = 326;
	{8'd10,8'd107} : s = 436;
	{8'd10,8'd108} : s = 434;
	{8'd10,8'd109} : s = 497;
	{8'd10,8'd110} : s = 325;
	{8'd10,8'd111} : s = 433;
	{8'd10,8'd112} : s = 428;
	{8'd10,8'd113} : s = 492;
	{8'd10,8'd114} : s = 426;
	{8'd10,8'd115} : s = 490;
	{8'd10,8'd116} : s = 489;
	{8'd10,8'd117} : s = 508;
	{8'd10,8'd118} : s = 2;
	{8'd10,8'd119} : s = 48;
	{8'd10,8'd120} : s = 40;
	{8'd10,8'd121} : s = 168;
	{8'd10,8'd122} : s = 36;
	{8'd10,8'd123} : s = 164;
	{8'd10,8'd124} : s = 162;
	{8'd10,8'd125} : s = 323;
	{8'd10,8'd126} : s = 34;
	{8'd10,8'd127} : s = 161;
	{8'd10,8'd128} : s = 152;
	{8'd10,8'd129} : s = 312;
	{8'd10,8'd130} : s = 148;
	{8'd10,8'd131} : s = 308;
	{8'd10,8'd132} : s = 306;
	{8'd10,8'd133} : s = 425;
	{8'd10,8'd134} : s = 33;
	{8'd10,8'd135} : s = 146;
	{8'd10,8'd136} : s = 145;
	{8'd10,8'd137} : s = 305;
	{8'd10,8'd138} : s = 140;
	{8'd10,8'd139} : s = 300;
	{8'd10,8'd140} : s = 298;
	{8'd10,8'd141} : s = 422;
	{8'd10,8'd142} : s = 138;
	{8'd10,8'd143} : s = 297;
	{8'd10,8'd144} : s = 294;
	{8'd10,8'd145} : s = 421;
	{8'd10,8'd146} : s = 293;
	{8'd10,8'd147} : s = 419;
	{8'd10,8'd148} : s = 412;
	{8'd10,8'd149} : s = 486;
	{8'd10,8'd150} : s = 24;
	{8'd10,8'd151} : s = 137;
	{8'd10,8'd152} : s = 134;
	{8'd10,8'd153} : s = 291;
	{8'd10,8'd154} : s = 133;
	{8'd10,8'd155} : s = 284;
	{8'd10,8'd156} : s = 282;
	{8'd10,8'd157} : s = 410;
	{8'd10,8'd158} : s = 131;
	{8'd10,8'd159} : s = 281;
	{8'd10,8'd160} : s = 278;
	{8'd10,8'd161} : s = 409;
	{8'd10,8'd162} : s = 277;
	{8'd10,8'd163} : s = 406;
	{8'd10,8'd164} : s = 405;
	{8'd10,8'd165} : s = 485;
	{8'd10,8'd166} : s = 112;
	{8'd10,8'd167} : s = 275;
	{8'd10,8'd168} : s = 270;
	{8'd10,8'd169} : s = 403;
	{8'd10,8'd170} : s = 269;
	{8'd10,8'd171} : s = 398;
	{8'd10,8'd172} : s = 397;
	{8'd10,8'd173} : s = 483;
	{8'd10,8'd174} : s = 267;
	{8'd10,8'd175} : s = 395;
	{8'd10,8'd176} : s = 391;
	{8'd10,8'd177} : s = 476;
	{8'd10,8'd178} : s = 376;
	{8'd10,8'd179} : s = 474;
	{8'd10,8'd180} : s = 473;
	{8'd10,8'd181} : s = 506;
	{8'd10,8'd182} : s = 20;
	{8'd10,8'd183} : s = 104;
	{8'd10,8'd184} : s = 100;
	{8'd10,8'd185} : s = 263;
	{8'd10,8'd186} : s = 98;
	{8'd10,8'd187} : s = 240;
	{8'd10,8'd188} : s = 232;
	{8'd10,8'd189} : s = 372;
	{8'd10,8'd190} : s = 97;
	{8'd10,8'd191} : s = 228;
	{8'd10,8'd192} : s = 226;
	{8'd10,8'd193} : s = 370;
	{8'd10,8'd194} : s = 225;
	{8'd10,8'd195} : s = 369;
	{8'd10,8'd196} : s = 364;
	{8'd10,8'd197} : s = 470;
	{8'd10,8'd198} : s = 88;
	{8'd10,8'd199} : s = 216;
	{8'd10,8'd200} : s = 212;
	{8'd10,8'd201} : s = 362;
	{8'd10,8'd202} : s = 210;
	{8'd10,8'd203} : s = 361;
	{8'd10,8'd204} : s = 358;
	{8'd10,8'd205} : s = 469;
	{8'd10,8'd206} : s = 209;
	{8'd10,8'd207} : s = 357;
	{8'd10,8'd208} : s = 355;
	{8'd10,8'd209} : s = 467;
	{8'd10,8'd210} : s = 348;
	{8'd10,8'd211} : s = 462;
	{8'd10,8'd212} : s = 461;
	{8'd10,8'd213} : s = 505;
	{8'd10,8'd214} : s = 84;
	{8'd10,8'd215} : s = 204;
	{8'd10,8'd216} : s = 202;
	{8'd10,8'd217} : s = 346;
	{8'd10,8'd218} : s = 201;
	{8'd10,8'd219} : s = 345;
	{8'd10,8'd220} : s = 342;
	{8'd10,8'd221} : s = 459;
	{8'd10,8'd222} : s = 198;
	{8'd10,8'd223} : s = 341;
	{8'd10,8'd224} : s = 339;
	{8'd10,8'd225} : s = 455;
	{8'd10,8'd226} : s = 334;
	{8'd10,8'd227} : s = 444;
	{8'd10,8'd228} : s = 442;
	{8'd10,8'd229} : s = 502;
	{8'd10,8'd230} : s = 197;
	{8'd10,8'd231} : s = 333;
	{8'd10,8'd232} : s = 331;
	{8'd10,8'd233} : s = 441;
	{8'd10,8'd234} : s = 327;
	{8'd10,8'd235} : s = 438;
	{8'd10,8'd236} : s = 437;
	{8'd10,8'd237} : s = 501;
	{8'd10,8'd238} : s = 316;
	{8'd10,8'd239} : s = 435;
	{8'd10,8'd240} : s = 430;
	{8'd10,8'd241} : s = 499;
	{8'd10,8'd242} : s = 429;
	{8'd10,8'd243} : s = 494;
	{8'd10,8'd244} : s = 493;
	{8'd10,8'd245} : s = 510;
	{8'd10,8'd246} : s = 1;
	{8'd10,8'd247} : s = 18;
	{8'd10,8'd248} : s = 17;
	{8'd10,8'd249} : s = 82;
	{8'd10,8'd250} : s = 12;
	{8'd10,8'd251} : s = 81;
	{8'd10,8'd252} : s = 76;
	{8'd10,8'd253} : s = 195;
	{8'd10,8'd254} : s = 10;
	{8'd10,8'd255} : s = 74;
	{8'd11,8'd0} : s = 416;
	{8'd11,8'd1} : s = 260;
	{8'd11,8'd2} : s = 400;
	{8'd11,8'd3} : s = 392;
	{8'd11,8'd4} : s = 480;
	{8'd11,8'd5} : s = 8;
	{8'd11,8'd6} : s = 258;
	{8'd11,8'd7} : s = 257;
	{8'd11,8'd8} : s = 388;
	{8'd11,8'd9} : s = 192;
	{8'd11,8'd10} : s = 386;
	{8'd11,8'd11} : s = 385;
	{8'd11,8'd12} : s = 464;
	{8'd11,8'd13} : s = 160;
	{8'd11,8'd14} : s = 352;
	{8'd11,8'd15} : s = 336;
	{8'd11,8'd16} : s = 456;
	{8'd11,8'd17} : s = 328;
	{8'd11,8'd18} : s = 452;
	{8'd11,8'd19} : s = 450;
	{8'd11,8'd20} : s = 496;
	{8'd11,8'd21} : s = 16;
	{8'd11,8'd22} : s = 144;
	{8'd11,8'd23} : s = 136;
	{8'd11,8'd24} : s = 324;
	{8'd11,8'd25} : s = 132;
	{8'd11,8'd26} : s = 322;
	{8'd11,8'd27} : s = 321;
	{8'd11,8'd28} : s = 449;
	{8'd11,8'd29} : s = 130;
	{8'd11,8'd30} : s = 304;
	{8'd11,8'd31} : s = 296;
	{8'd11,8'd32} : s = 432;
	{8'd11,8'd33} : s = 292;
	{8'd11,8'd34} : s = 424;
	{8'd11,8'd35} : s = 420;
	{8'd11,8'd36} : s = 488;
	{8'd11,8'd37} : s = 129;
	{8'd11,8'd38} : s = 290;
	{8'd11,8'd39} : s = 289;
	{8'd11,8'd40} : s = 418;
	{8'd11,8'd41} : s = 280;
	{8'd11,8'd42} : s = 417;
	{8'd11,8'd43} : s = 408;
	{8'd11,8'd44} : s = 484;
	{8'd11,8'd45} : s = 276;
	{8'd11,8'd46} : s = 404;
	{8'd11,8'd47} : s = 402;
	{8'd11,8'd48} : s = 482;
	{8'd11,8'd49} : s = 401;
	{8'd11,8'd50} : s = 481;
	{8'd11,8'd51} : s = 472;
	{8'd11,8'd52} : s = 504;
	{8'd11,8'd53} : s = 4;
	{8'd11,8'd54} : s = 96;
	{8'd11,8'd55} : s = 80;
	{8'd11,8'd56} : s = 274;
	{8'd11,8'd57} : s = 72;
	{8'd11,8'd58} : s = 273;
	{8'd11,8'd59} : s = 268;
	{8'd11,8'd60} : s = 396;
	{8'd11,8'd61} : s = 68;
	{8'd11,8'd62} : s = 266;
	{8'd11,8'd63} : s = 265;
	{8'd11,8'd64} : s = 394;
	{8'd11,8'd65} : s = 262;
	{8'd11,8'd66} : s = 393;
	{8'd11,8'd67} : s = 390;
	{8'd11,8'd68} : s = 468;
	{8'd11,8'd69} : s = 66;
	{8'd11,8'd70} : s = 261;
	{8'd11,8'd71} : s = 259;
	{8'd11,8'd72} : s = 389;
	{8'd11,8'd73} : s = 224;
	{8'd11,8'd74} : s = 387;
	{8'd11,8'd75} : s = 368;
	{8'd11,8'd76} : s = 466;
	{8'd11,8'd77} : s = 208;
	{8'd11,8'd78} : s = 360;
	{8'd11,8'd79} : s = 356;
	{8'd11,8'd80} : s = 465;
	{8'd11,8'd81} : s = 354;
	{8'd11,8'd82} : s = 460;
	{8'd11,8'd83} : s = 458;
	{8'd11,8'd84} : s = 500;
	{8'd11,8'd85} : s = 65;
	{8'd11,8'd86} : s = 200;
	{8'd11,8'd87} : s = 196;
	{8'd11,8'd88} : s = 353;
	{8'd11,8'd89} : s = 194;
	{8'd11,8'd90} : s = 344;
	{8'd11,8'd91} : s = 340;
	{8'd11,8'd92} : s = 457;
	{8'd11,8'd93} : s = 193;
	{8'd11,8'd94} : s = 338;
	{8'd11,8'd95} : s = 337;
	{8'd11,8'd96} : s = 454;
	{8'd11,8'd97} : s = 332;
	{8'd11,8'd98} : s = 453;
	{8'd11,8'd99} : s = 451;
	{8'd11,8'd100} : s = 498;
	{8'd11,8'd101} : s = 176;
	{8'd11,8'd102} : s = 330;
	{8'd11,8'd103} : s = 329;
	{8'd11,8'd104} : s = 440;
	{8'd11,8'd105} : s = 326;
	{8'd11,8'd106} : s = 436;
	{8'd11,8'd107} : s = 434;
	{8'd11,8'd108} : s = 497;
	{8'd11,8'd109} : s = 325;
	{8'd11,8'd110} : s = 433;
	{8'd11,8'd111} : s = 428;
	{8'd11,8'd112} : s = 492;
	{8'd11,8'd113} : s = 426;
	{8'd11,8'd114} : s = 490;
	{8'd11,8'd115} : s = 489;
	{8'd11,8'd116} : s = 508;
	{8'd11,8'd117} : s = 2;
	{8'd11,8'd118} : s = 48;
	{8'd11,8'd119} : s = 40;
	{8'd11,8'd120} : s = 168;
	{8'd11,8'd121} : s = 36;
	{8'd11,8'd122} : s = 164;
	{8'd11,8'd123} : s = 162;
	{8'd11,8'd124} : s = 323;
	{8'd11,8'd125} : s = 34;
	{8'd11,8'd126} : s = 161;
	{8'd11,8'd127} : s = 152;
	{8'd11,8'd128} : s = 312;
	{8'd11,8'd129} : s = 148;
	{8'd11,8'd130} : s = 308;
	{8'd11,8'd131} : s = 306;
	{8'd11,8'd132} : s = 425;
	{8'd11,8'd133} : s = 33;
	{8'd11,8'd134} : s = 146;
	{8'd11,8'd135} : s = 145;
	{8'd11,8'd136} : s = 305;
	{8'd11,8'd137} : s = 140;
	{8'd11,8'd138} : s = 300;
	{8'd11,8'd139} : s = 298;
	{8'd11,8'd140} : s = 422;
	{8'd11,8'd141} : s = 138;
	{8'd11,8'd142} : s = 297;
	{8'd11,8'd143} : s = 294;
	{8'd11,8'd144} : s = 421;
	{8'd11,8'd145} : s = 293;
	{8'd11,8'd146} : s = 419;
	{8'd11,8'd147} : s = 412;
	{8'd11,8'd148} : s = 486;
	{8'd11,8'd149} : s = 24;
	{8'd11,8'd150} : s = 137;
	{8'd11,8'd151} : s = 134;
	{8'd11,8'd152} : s = 291;
	{8'd11,8'd153} : s = 133;
	{8'd11,8'd154} : s = 284;
	{8'd11,8'd155} : s = 282;
	{8'd11,8'd156} : s = 410;
	{8'd11,8'd157} : s = 131;
	{8'd11,8'd158} : s = 281;
	{8'd11,8'd159} : s = 278;
	{8'd11,8'd160} : s = 409;
	{8'd11,8'd161} : s = 277;
	{8'd11,8'd162} : s = 406;
	{8'd11,8'd163} : s = 405;
	{8'd11,8'd164} : s = 485;
	{8'd11,8'd165} : s = 112;
	{8'd11,8'd166} : s = 275;
	{8'd11,8'd167} : s = 270;
	{8'd11,8'd168} : s = 403;
	{8'd11,8'd169} : s = 269;
	{8'd11,8'd170} : s = 398;
	{8'd11,8'd171} : s = 397;
	{8'd11,8'd172} : s = 483;
	{8'd11,8'd173} : s = 267;
	{8'd11,8'd174} : s = 395;
	{8'd11,8'd175} : s = 391;
	{8'd11,8'd176} : s = 476;
	{8'd11,8'd177} : s = 376;
	{8'd11,8'd178} : s = 474;
	{8'd11,8'd179} : s = 473;
	{8'd11,8'd180} : s = 506;
	{8'd11,8'd181} : s = 20;
	{8'd11,8'd182} : s = 104;
	{8'd11,8'd183} : s = 100;
	{8'd11,8'd184} : s = 263;
	{8'd11,8'd185} : s = 98;
	{8'd11,8'd186} : s = 240;
	{8'd11,8'd187} : s = 232;
	{8'd11,8'd188} : s = 372;
	{8'd11,8'd189} : s = 97;
	{8'd11,8'd190} : s = 228;
	{8'd11,8'd191} : s = 226;
	{8'd11,8'd192} : s = 370;
	{8'd11,8'd193} : s = 225;
	{8'd11,8'd194} : s = 369;
	{8'd11,8'd195} : s = 364;
	{8'd11,8'd196} : s = 470;
	{8'd11,8'd197} : s = 88;
	{8'd11,8'd198} : s = 216;
	{8'd11,8'd199} : s = 212;
	{8'd11,8'd200} : s = 362;
	{8'd11,8'd201} : s = 210;
	{8'd11,8'd202} : s = 361;
	{8'd11,8'd203} : s = 358;
	{8'd11,8'd204} : s = 469;
	{8'd11,8'd205} : s = 209;
	{8'd11,8'd206} : s = 357;
	{8'd11,8'd207} : s = 355;
	{8'd11,8'd208} : s = 467;
	{8'd11,8'd209} : s = 348;
	{8'd11,8'd210} : s = 462;
	{8'd11,8'd211} : s = 461;
	{8'd11,8'd212} : s = 505;
	{8'd11,8'd213} : s = 84;
	{8'd11,8'd214} : s = 204;
	{8'd11,8'd215} : s = 202;
	{8'd11,8'd216} : s = 346;
	{8'd11,8'd217} : s = 201;
	{8'd11,8'd218} : s = 345;
	{8'd11,8'd219} : s = 342;
	{8'd11,8'd220} : s = 459;
	{8'd11,8'd221} : s = 198;
	{8'd11,8'd222} : s = 341;
	{8'd11,8'd223} : s = 339;
	{8'd11,8'd224} : s = 455;
	{8'd11,8'd225} : s = 334;
	{8'd11,8'd226} : s = 444;
	{8'd11,8'd227} : s = 442;
	{8'd11,8'd228} : s = 502;
	{8'd11,8'd229} : s = 197;
	{8'd11,8'd230} : s = 333;
	{8'd11,8'd231} : s = 331;
	{8'd11,8'd232} : s = 441;
	{8'd11,8'd233} : s = 327;
	{8'd11,8'd234} : s = 438;
	{8'd11,8'd235} : s = 437;
	{8'd11,8'd236} : s = 501;
	{8'd11,8'd237} : s = 316;
	{8'd11,8'd238} : s = 435;
	{8'd11,8'd239} : s = 430;
	{8'd11,8'd240} : s = 499;
	{8'd11,8'd241} : s = 429;
	{8'd11,8'd242} : s = 494;
	{8'd11,8'd243} : s = 493;
	{8'd11,8'd244} : s = 510;
	{8'd11,8'd245} : s = 1;
	{8'd11,8'd246} : s = 18;
	{8'd11,8'd247} : s = 17;
	{8'd11,8'd248} : s = 82;
	{8'd11,8'd249} : s = 12;
	{8'd11,8'd250} : s = 81;
	{8'd11,8'd251} : s = 76;
	{8'd11,8'd252} : s = 195;
	{8'd11,8'd253} : s = 10;
	{8'd11,8'd254} : s = 74;
	{8'd11,8'd255} : s = 73;
	{8'd12,8'd0} : s = 260;
	{8'd12,8'd1} : s = 400;
	{8'd12,8'd2} : s = 392;
	{8'd12,8'd3} : s = 480;
	{8'd12,8'd4} : s = 8;
	{8'd12,8'd5} : s = 258;
	{8'd12,8'd6} : s = 257;
	{8'd12,8'd7} : s = 388;
	{8'd12,8'd8} : s = 192;
	{8'd12,8'd9} : s = 386;
	{8'd12,8'd10} : s = 385;
	{8'd12,8'd11} : s = 464;
	{8'd12,8'd12} : s = 160;
	{8'd12,8'd13} : s = 352;
	{8'd12,8'd14} : s = 336;
	{8'd12,8'd15} : s = 456;
	{8'd12,8'd16} : s = 328;
	{8'd12,8'd17} : s = 452;
	{8'd12,8'd18} : s = 450;
	{8'd12,8'd19} : s = 496;
	{8'd12,8'd20} : s = 16;
	{8'd12,8'd21} : s = 144;
	{8'd12,8'd22} : s = 136;
	{8'd12,8'd23} : s = 324;
	{8'd12,8'd24} : s = 132;
	{8'd12,8'd25} : s = 322;
	{8'd12,8'd26} : s = 321;
	{8'd12,8'd27} : s = 449;
	{8'd12,8'd28} : s = 130;
	{8'd12,8'd29} : s = 304;
	{8'd12,8'd30} : s = 296;
	{8'd12,8'd31} : s = 432;
	{8'd12,8'd32} : s = 292;
	{8'd12,8'd33} : s = 424;
	{8'd12,8'd34} : s = 420;
	{8'd12,8'd35} : s = 488;
	{8'd12,8'd36} : s = 129;
	{8'd12,8'd37} : s = 290;
	{8'd12,8'd38} : s = 289;
	{8'd12,8'd39} : s = 418;
	{8'd12,8'd40} : s = 280;
	{8'd12,8'd41} : s = 417;
	{8'd12,8'd42} : s = 408;
	{8'd12,8'd43} : s = 484;
	{8'd12,8'd44} : s = 276;
	{8'd12,8'd45} : s = 404;
	{8'd12,8'd46} : s = 402;
	{8'd12,8'd47} : s = 482;
	{8'd12,8'd48} : s = 401;
	{8'd12,8'd49} : s = 481;
	{8'd12,8'd50} : s = 472;
	{8'd12,8'd51} : s = 504;
	{8'd12,8'd52} : s = 4;
	{8'd12,8'd53} : s = 96;
	{8'd12,8'd54} : s = 80;
	{8'd12,8'd55} : s = 274;
	{8'd12,8'd56} : s = 72;
	{8'd12,8'd57} : s = 273;
	{8'd12,8'd58} : s = 268;
	{8'd12,8'd59} : s = 396;
	{8'd12,8'd60} : s = 68;
	{8'd12,8'd61} : s = 266;
	{8'd12,8'd62} : s = 265;
	{8'd12,8'd63} : s = 394;
	{8'd12,8'd64} : s = 262;
	{8'd12,8'd65} : s = 393;
	{8'd12,8'd66} : s = 390;
	{8'd12,8'd67} : s = 468;
	{8'd12,8'd68} : s = 66;
	{8'd12,8'd69} : s = 261;
	{8'd12,8'd70} : s = 259;
	{8'd12,8'd71} : s = 389;
	{8'd12,8'd72} : s = 224;
	{8'd12,8'd73} : s = 387;
	{8'd12,8'd74} : s = 368;
	{8'd12,8'd75} : s = 466;
	{8'd12,8'd76} : s = 208;
	{8'd12,8'd77} : s = 360;
	{8'd12,8'd78} : s = 356;
	{8'd12,8'd79} : s = 465;
	{8'd12,8'd80} : s = 354;
	{8'd12,8'd81} : s = 460;
	{8'd12,8'd82} : s = 458;
	{8'd12,8'd83} : s = 500;
	{8'd12,8'd84} : s = 65;
	{8'd12,8'd85} : s = 200;
	{8'd12,8'd86} : s = 196;
	{8'd12,8'd87} : s = 353;
	{8'd12,8'd88} : s = 194;
	{8'd12,8'd89} : s = 344;
	{8'd12,8'd90} : s = 340;
	{8'd12,8'd91} : s = 457;
	{8'd12,8'd92} : s = 193;
	{8'd12,8'd93} : s = 338;
	{8'd12,8'd94} : s = 337;
	{8'd12,8'd95} : s = 454;
	{8'd12,8'd96} : s = 332;
	{8'd12,8'd97} : s = 453;
	{8'd12,8'd98} : s = 451;
	{8'd12,8'd99} : s = 498;
	{8'd12,8'd100} : s = 176;
	{8'd12,8'd101} : s = 330;
	{8'd12,8'd102} : s = 329;
	{8'd12,8'd103} : s = 440;
	{8'd12,8'd104} : s = 326;
	{8'd12,8'd105} : s = 436;
	{8'd12,8'd106} : s = 434;
	{8'd12,8'd107} : s = 497;
	{8'd12,8'd108} : s = 325;
	{8'd12,8'd109} : s = 433;
	{8'd12,8'd110} : s = 428;
	{8'd12,8'd111} : s = 492;
	{8'd12,8'd112} : s = 426;
	{8'd12,8'd113} : s = 490;
	{8'd12,8'd114} : s = 489;
	{8'd12,8'd115} : s = 508;
	{8'd12,8'd116} : s = 2;
	{8'd12,8'd117} : s = 48;
	{8'd12,8'd118} : s = 40;
	{8'd12,8'd119} : s = 168;
	{8'd12,8'd120} : s = 36;
	{8'd12,8'd121} : s = 164;
	{8'd12,8'd122} : s = 162;
	{8'd12,8'd123} : s = 323;
	{8'd12,8'd124} : s = 34;
	{8'd12,8'd125} : s = 161;
	{8'd12,8'd126} : s = 152;
	{8'd12,8'd127} : s = 312;
	{8'd12,8'd128} : s = 148;
	{8'd12,8'd129} : s = 308;
	{8'd12,8'd130} : s = 306;
	{8'd12,8'd131} : s = 425;
	{8'd12,8'd132} : s = 33;
	{8'd12,8'd133} : s = 146;
	{8'd12,8'd134} : s = 145;
	{8'd12,8'd135} : s = 305;
	{8'd12,8'd136} : s = 140;
	{8'd12,8'd137} : s = 300;
	{8'd12,8'd138} : s = 298;
	{8'd12,8'd139} : s = 422;
	{8'd12,8'd140} : s = 138;
	{8'd12,8'd141} : s = 297;
	{8'd12,8'd142} : s = 294;
	{8'd12,8'd143} : s = 421;
	{8'd12,8'd144} : s = 293;
	{8'd12,8'd145} : s = 419;
	{8'd12,8'd146} : s = 412;
	{8'd12,8'd147} : s = 486;
	{8'd12,8'd148} : s = 24;
	{8'd12,8'd149} : s = 137;
	{8'd12,8'd150} : s = 134;
	{8'd12,8'd151} : s = 291;
	{8'd12,8'd152} : s = 133;
	{8'd12,8'd153} : s = 284;
	{8'd12,8'd154} : s = 282;
	{8'd12,8'd155} : s = 410;
	{8'd12,8'd156} : s = 131;
	{8'd12,8'd157} : s = 281;
	{8'd12,8'd158} : s = 278;
	{8'd12,8'd159} : s = 409;
	{8'd12,8'd160} : s = 277;
	{8'd12,8'd161} : s = 406;
	{8'd12,8'd162} : s = 405;
	{8'd12,8'd163} : s = 485;
	{8'd12,8'd164} : s = 112;
	{8'd12,8'd165} : s = 275;
	{8'd12,8'd166} : s = 270;
	{8'd12,8'd167} : s = 403;
	{8'd12,8'd168} : s = 269;
	{8'd12,8'd169} : s = 398;
	{8'd12,8'd170} : s = 397;
	{8'd12,8'd171} : s = 483;
	{8'd12,8'd172} : s = 267;
	{8'd12,8'd173} : s = 395;
	{8'd12,8'd174} : s = 391;
	{8'd12,8'd175} : s = 476;
	{8'd12,8'd176} : s = 376;
	{8'd12,8'd177} : s = 474;
	{8'd12,8'd178} : s = 473;
	{8'd12,8'd179} : s = 506;
	{8'd12,8'd180} : s = 20;
	{8'd12,8'd181} : s = 104;
	{8'd12,8'd182} : s = 100;
	{8'd12,8'd183} : s = 263;
	{8'd12,8'd184} : s = 98;
	{8'd12,8'd185} : s = 240;
	{8'd12,8'd186} : s = 232;
	{8'd12,8'd187} : s = 372;
	{8'd12,8'd188} : s = 97;
	{8'd12,8'd189} : s = 228;
	{8'd12,8'd190} : s = 226;
	{8'd12,8'd191} : s = 370;
	{8'd12,8'd192} : s = 225;
	{8'd12,8'd193} : s = 369;
	{8'd12,8'd194} : s = 364;
	{8'd12,8'd195} : s = 470;
	{8'd12,8'd196} : s = 88;
	{8'd12,8'd197} : s = 216;
	{8'd12,8'd198} : s = 212;
	{8'd12,8'd199} : s = 362;
	{8'd12,8'd200} : s = 210;
	{8'd12,8'd201} : s = 361;
	{8'd12,8'd202} : s = 358;
	{8'd12,8'd203} : s = 469;
	{8'd12,8'd204} : s = 209;
	{8'd12,8'd205} : s = 357;
	{8'd12,8'd206} : s = 355;
	{8'd12,8'd207} : s = 467;
	{8'd12,8'd208} : s = 348;
	{8'd12,8'd209} : s = 462;
	{8'd12,8'd210} : s = 461;
	{8'd12,8'd211} : s = 505;
	{8'd12,8'd212} : s = 84;
	{8'd12,8'd213} : s = 204;
	{8'd12,8'd214} : s = 202;
	{8'd12,8'd215} : s = 346;
	{8'd12,8'd216} : s = 201;
	{8'd12,8'd217} : s = 345;
	{8'd12,8'd218} : s = 342;
	{8'd12,8'd219} : s = 459;
	{8'd12,8'd220} : s = 198;
	{8'd12,8'd221} : s = 341;
	{8'd12,8'd222} : s = 339;
	{8'd12,8'd223} : s = 455;
	{8'd12,8'd224} : s = 334;
	{8'd12,8'd225} : s = 444;
	{8'd12,8'd226} : s = 442;
	{8'd12,8'd227} : s = 502;
	{8'd12,8'd228} : s = 197;
	{8'd12,8'd229} : s = 333;
	{8'd12,8'd230} : s = 331;
	{8'd12,8'd231} : s = 441;
	{8'd12,8'd232} : s = 327;
	{8'd12,8'd233} : s = 438;
	{8'd12,8'd234} : s = 437;
	{8'd12,8'd235} : s = 501;
	{8'd12,8'd236} : s = 316;
	{8'd12,8'd237} : s = 435;
	{8'd12,8'd238} : s = 430;
	{8'd12,8'd239} : s = 499;
	{8'd12,8'd240} : s = 429;
	{8'd12,8'd241} : s = 494;
	{8'd12,8'd242} : s = 493;
	{8'd12,8'd243} : s = 510;
	{8'd12,8'd244} : s = 1;
	{8'd12,8'd245} : s = 18;
	{8'd12,8'd246} : s = 17;
	{8'd12,8'd247} : s = 82;
	{8'd12,8'd248} : s = 12;
	{8'd12,8'd249} : s = 81;
	{8'd12,8'd250} : s = 76;
	{8'd12,8'd251} : s = 195;
	{8'd12,8'd252} : s = 10;
	{8'd12,8'd253} : s = 74;
	{8'd12,8'd254} : s = 73;
	{8'd12,8'd255} : s = 184;
	{8'd13,8'd0} : s = 400;
	{8'd13,8'd1} : s = 392;
	{8'd13,8'd2} : s = 480;
	{8'd13,8'd3} : s = 8;
	{8'd13,8'd4} : s = 258;
	{8'd13,8'd5} : s = 257;
	{8'd13,8'd6} : s = 388;
	{8'd13,8'd7} : s = 192;
	{8'd13,8'd8} : s = 386;
	{8'd13,8'd9} : s = 385;
	{8'd13,8'd10} : s = 464;
	{8'd13,8'd11} : s = 160;
	{8'd13,8'd12} : s = 352;
	{8'd13,8'd13} : s = 336;
	{8'd13,8'd14} : s = 456;
	{8'd13,8'd15} : s = 328;
	{8'd13,8'd16} : s = 452;
	{8'd13,8'd17} : s = 450;
	{8'd13,8'd18} : s = 496;
	{8'd13,8'd19} : s = 16;
	{8'd13,8'd20} : s = 144;
	{8'd13,8'd21} : s = 136;
	{8'd13,8'd22} : s = 324;
	{8'd13,8'd23} : s = 132;
	{8'd13,8'd24} : s = 322;
	{8'd13,8'd25} : s = 321;
	{8'd13,8'd26} : s = 449;
	{8'd13,8'd27} : s = 130;
	{8'd13,8'd28} : s = 304;
	{8'd13,8'd29} : s = 296;
	{8'd13,8'd30} : s = 432;
	{8'd13,8'd31} : s = 292;
	{8'd13,8'd32} : s = 424;
	{8'd13,8'd33} : s = 420;
	{8'd13,8'd34} : s = 488;
	{8'd13,8'd35} : s = 129;
	{8'd13,8'd36} : s = 290;
	{8'd13,8'd37} : s = 289;
	{8'd13,8'd38} : s = 418;
	{8'd13,8'd39} : s = 280;
	{8'd13,8'd40} : s = 417;
	{8'd13,8'd41} : s = 408;
	{8'd13,8'd42} : s = 484;
	{8'd13,8'd43} : s = 276;
	{8'd13,8'd44} : s = 404;
	{8'd13,8'd45} : s = 402;
	{8'd13,8'd46} : s = 482;
	{8'd13,8'd47} : s = 401;
	{8'd13,8'd48} : s = 481;
	{8'd13,8'd49} : s = 472;
	{8'd13,8'd50} : s = 504;
	{8'd13,8'd51} : s = 4;
	{8'd13,8'd52} : s = 96;
	{8'd13,8'd53} : s = 80;
	{8'd13,8'd54} : s = 274;
	{8'd13,8'd55} : s = 72;
	{8'd13,8'd56} : s = 273;
	{8'd13,8'd57} : s = 268;
	{8'd13,8'd58} : s = 396;
	{8'd13,8'd59} : s = 68;
	{8'd13,8'd60} : s = 266;
	{8'd13,8'd61} : s = 265;
	{8'd13,8'd62} : s = 394;
	{8'd13,8'd63} : s = 262;
	{8'd13,8'd64} : s = 393;
	{8'd13,8'd65} : s = 390;
	{8'd13,8'd66} : s = 468;
	{8'd13,8'd67} : s = 66;
	{8'd13,8'd68} : s = 261;
	{8'd13,8'd69} : s = 259;
	{8'd13,8'd70} : s = 389;
	{8'd13,8'd71} : s = 224;
	{8'd13,8'd72} : s = 387;
	{8'd13,8'd73} : s = 368;
	{8'd13,8'd74} : s = 466;
	{8'd13,8'd75} : s = 208;
	{8'd13,8'd76} : s = 360;
	{8'd13,8'd77} : s = 356;
	{8'd13,8'd78} : s = 465;
	{8'd13,8'd79} : s = 354;
	{8'd13,8'd80} : s = 460;
	{8'd13,8'd81} : s = 458;
	{8'd13,8'd82} : s = 500;
	{8'd13,8'd83} : s = 65;
	{8'd13,8'd84} : s = 200;
	{8'd13,8'd85} : s = 196;
	{8'd13,8'd86} : s = 353;
	{8'd13,8'd87} : s = 194;
	{8'd13,8'd88} : s = 344;
	{8'd13,8'd89} : s = 340;
	{8'd13,8'd90} : s = 457;
	{8'd13,8'd91} : s = 193;
	{8'd13,8'd92} : s = 338;
	{8'd13,8'd93} : s = 337;
	{8'd13,8'd94} : s = 454;
	{8'd13,8'd95} : s = 332;
	{8'd13,8'd96} : s = 453;
	{8'd13,8'd97} : s = 451;
	{8'd13,8'd98} : s = 498;
	{8'd13,8'd99} : s = 176;
	{8'd13,8'd100} : s = 330;
	{8'd13,8'd101} : s = 329;
	{8'd13,8'd102} : s = 440;
	{8'd13,8'd103} : s = 326;
	{8'd13,8'd104} : s = 436;
	{8'd13,8'd105} : s = 434;
	{8'd13,8'd106} : s = 497;
	{8'd13,8'd107} : s = 325;
	{8'd13,8'd108} : s = 433;
	{8'd13,8'd109} : s = 428;
	{8'd13,8'd110} : s = 492;
	{8'd13,8'd111} : s = 426;
	{8'd13,8'd112} : s = 490;
	{8'd13,8'd113} : s = 489;
	{8'd13,8'd114} : s = 508;
	{8'd13,8'd115} : s = 2;
	{8'd13,8'd116} : s = 48;
	{8'd13,8'd117} : s = 40;
	{8'd13,8'd118} : s = 168;
	{8'd13,8'd119} : s = 36;
	{8'd13,8'd120} : s = 164;
	{8'd13,8'd121} : s = 162;
	{8'd13,8'd122} : s = 323;
	{8'd13,8'd123} : s = 34;
	{8'd13,8'd124} : s = 161;
	{8'd13,8'd125} : s = 152;
	{8'd13,8'd126} : s = 312;
	{8'd13,8'd127} : s = 148;
	{8'd13,8'd128} : s = 308;
	{8'd13,8'd129} : s = 306;
	{8'd13,8'd130} : s = 425;
	{8'd13,8'd131} : s = 33;
	{8'd13,8'd132} : s = 146;
	{8'd13,8'd133} : s = 145;
	{8'd13,8'd134} : s = 305;
	{8'd13,8'd135} : s = 140;
	{8'd13,8'd136} : s = 300;
	{8'd13,8'd137} : s = 298;
	{8'd13,8'd138} : s = 422;
	{8'd13,8'd139} : s = 138;
	{8'd13,8'd140} : s = 297;
	{8'd13,8'd141} : s = 294;
	{8'd13,8'd142} : s = 421;
	{8'd13,8'd143} : s = 293;
	{8'd13,8'd144} : s = 419;
	{8'd13,8'd145} : s = 412;
	{8'd13,8'd146} : s = 486;
	{8'd13,8'd147} : s = 24;
	{8'd13,8'd148} : s = 137;
	{8'd13,8'd149} : s = 134;
	{8'd13,8'd150} : s = 291;
	{8'd13,8'd151} : s = 133;
	{8'd13,8'd152} : s = 284;
	{8'd13,8'd153} : s = 282;
	{8'd13,8'd154} : s = 410;
	{8'd13,8'd155} : s = 131;
	{8'd13,8'd156} : s = 281;
	{8'd13,8'd157} : s = 278;
	{8'd13,8'd158} : s = 409;
	{8'd13,8'd159} : s = 277;
	{8'd13,8'd160} : s = 406;
	{8'd13,8'd161} : s = 405;
	{8'd13,8'd162} : s = 485;
	{8'd13,8'd163} : s = 112;
	{8'd13,8'd164} : s = 275;
	{8'd13,8'd165} : s = 270;
	{8'd13,8'd166} : s = 403;
	{8'd13,8'd167} : s = 269;
	{8'd13,8'd168} : s = 398;
	{8'd13,8'd169} : s = 397;
	{8'd13,8'd170} : s = 483;
	{8'd13,8'd171} : s = 267;
	{8'd13,8'd172} : s = 395;
	{8'd13,8'd173} : s = 391;
	{8'd13,8'd174} : s = 476;
	{8'd13,8'd175} : s = 376;
	{8'd13,8'd176} : s = 474;
	{8'd13,8'd177} : s = 473;
	{8'd13,8'd178} : s = 506;
	{8'd13,8'd179} : s = 20;
	{8'd13,8'd180} : s = 104;
	{8'd13,8'd181} : s = 100;
	{8'd13,8'd182} : s = 263;
	{8'd13,8'd183} : s = 98;
	{8'd13,8'd184} : s = 240;
	{8'd13,8'd185} : s = 232;
	{8'd13,8'd186} : s = 372;
	{8'd13,8'd187} : s = 97;
	{8'd13,8'd188} : s = 228;
	{8'd13,8'd189} : s = 226;
	{8'd13,8'd190} : s = 370;
	{8'd13,8'd191} : s = 225;
	{8'd13,8'd192} : s = 369;
	{8'd13,8'd193} : s = 364;
	{8'd13,8'd194} : s = 470;
	{8'd13,8'd195} : s = 88;
	{8'd13,8'd196} : s = 216;
	{8'd13,8'd197} : s = 212;
	{8'd13,8'd198} : s = 362;
	{8'd13,8'd199} : s = 210;
	{8'd13,8'd200} : s = 361;
	{8'd13,8'd201} : s = 358;
	{8'd13,8'd202} : s = 469;
	{8'd13,8'd203} : s = 209;
	{8'd13,8'd204} : s = 357;
	{8'd13,8'd205} : s = 355;
	{8'd13,8'd206} : s = 467;
	{8'd13,8'd207} : s = 348;
	{8'd13,8'd208} : s = 462;
	{8'd13,8'd209} : s = 461;
	{8'd13,8'd210} : s = 505;
	{8'd13,8'd211} : s = 84;
	{8'd13,8'd212} : s = 204;
	{8'd13,8'd213} : s = 202;
	{8'd13,8'd214} : s = 346;
	{8'd13,8'd215} : s = 201;
	{8'd13,8'd216} : s = 345;
	{8'd13,8'd217} : s = 342;
	{8'd13,8'd218} : s = 459;
	{8'd13,8'd219} : s = 198;
	{8'd13,8'd220} : s = 341;
	{8'd13,8'd221} : s = 339;
	{8'd13,8'd222} : s = 455;
	{8'd13,8'd223} : s = 334;
	{8'd13,8'd224} : s = 444;
	{8'd13,8'd225} : s = 442;
	{8'd13,8'd226} : s = 502;
	{8'd13,8'd227} : s = 197;
	{8'd13,8'd228} : s = 333;
	{8'd13,8'd229} : s = 331;
	{8'd13,8'd230} : s = 441;
	{8'd13,8'd231} : s = 327;
	{8'd13,8'd232} : s = 438;
	{8'd13,8'd233} : s = 437;
	{8'd13,8'd234} : s = 501;
	{8'd13,8'd235} : s = 316;
	{8'd13,8'd236} : s = 435;
	{8'd13,8'd237} : s = 430;
	{8'd13,8'd238} : s = 499;
	{8'd13,8'd239} : s = 429;
	{8'd13,8'd240} : s = 494;
	{8'd13,8'd241} : s = 493;
	{8'd13,8'd242} : s = 510;
	{8'd13,8'd243} : s = 1;
	{8'd13,8'd244} : s = 18;
	{8'd13,8'd245} : s = 17;
	{8'd13,8'd246} : s = 82;
	{8'd13,8'd247} : s = 12;
	{8'd13,8'd248} : s = 81;
	{8'd13,8'd249} : s = 76;
	{8'd13,8'd250} : s = 195;
	{8'd13,8'd251} : s = 10;
	{8'd13,8'd252} : s = 74;
	{8'd13,8'd253} : s = 73;
	{8'd13,8'd254} : s = 184;
	{8'd13,8'd255} : s = 70;
	{8'd14,8'd0} : s = 392;
	{8'd14,8'd1} : s = 480;
	{8'd14,8'd2} : s = 8;
	{8'd14,8'd3} : s = 258;
	{8'd14,8'd4} : s = 257;
	{8'd14,8'd5} : s = 388;
	{8'd14,8'd6} : s = 192;
	{8'd14,8'd7} : s = 386;
	{8'd14,8'd8} : s = 385;
	{8'd14,8'd9} : s = 464;
	{8'd14,8'd10} : s = 160;
	{8'd14,8'd11} : s = 352;
	{8'd14,8'd12} : s = 336;
	{8'd14,8'd13} : s = 456;
	{8'd14,8'd14} : s = 328;
	{8'd14,8'd15} : s = 452;
	{8'd14,8'd16} : s = 450;
	{8'd14,8'd17} : s = 496;
	{8'd14,8'd18} : s = 16;
	{8'd14,8'd19} : s = 144;
	{8'd14,8'd20} : s = 136;
	{8'd14,8'd21} : s = 324;
	{8'd14,8'd22} : s = 132;
	{8'd14,8'd23} : s = 322;
	{8'd14,8'd24} : s = 321;
	{8'd14,8'd25} : s = 449;
	{8'd14,8'd26} : s = 130;
	{8'd14,8'd27} : s = 304;
	{8'd14,8'd28} : s = 296;
	{8'd14,8'd29} : s = 432;
	{8'd14,8'd30} : s = 292;
	{8'd14,8'd31} : s = 424;
	{8'd14,8'd32} : s = 420;
	{8'd14,8'd33} : s = 488;
	{8'd14,8'd34} : s = 129;
	{8'd14,8'd35} : s = 290;
	{8'd14,8'd36} : s = 289;
	{8'd14,8'd37} : s = 418;
	{8'd14,8'd38} : s = 280;
	{8'd14,8'd39} : s = 417;
	{8'd14,8'd40} : s = 408;
	{8'd14,8'd41} : s = 484;
	{8'd14,8'd42} : s = 276;
	{8'd14,8'd43} : s = 404;
	{8'd14,8'd44} : s = 402;
	{8'd14,8'd45} : s = 482;
	{8'd14,8'd46} : s = 401;
	{8'd14,8'd47} : s = 481;
	{8'd14,8'd48} : s = 472;
	{8'd14,8'd49} : s = 504;
	{8'd14,8'd50} : s = 4;
	{8'd14,8'd51} : s = 96;
	{8'd14,8'd52} : s = 80;
	{8'd14,8'd53} : s = 274;
	{8'd14,8'd54} : s = 72;
	{8'd14,8'd55} : s = 273;
	{8'd14,8'd56} : s = 268;
	{8'd14,8'd57} : s = 396;
	{8'd14,8'd58} : s = 68;
	{8'd14,8'd59} : s = 266;
	{8'd14,8'd60} : s = 265;
	{8'd14,8'd61} : s = 394;
	{8'd14,8'd62} : s = 262;
	{8'd14,8'd63} : s = 393;
	{8'd14,8'd64} : s = 390;
	{8'd14,8'd65} : s = 468;
	{8'd14,8'd66} : s = 66;
	{8'd14,8'd67} : s = 261;
	{8'd14,8'd68} : s = 259;
	{8'd14,8'd69} : s = 389;
	{8'd14,8'd70} : s = 224;
	{8'd14,8'd71} : s = 387;
	{8'd14,8'd72} : s = 368;
	{8'd14,8'd73} : s = 466;
	{8'd14,8'd74} : s = 208;
	{8'd14,8'd75} : s = 360;
	{8'd14,8'd76} : s = 356;
	{8'd14,8'd77} : s = 465;
	{8'd14,8'd78} : s = 354;
	{8'd14,8'd79} : s = 460;
	{8'd14,8'd80} : s = 458;
	{8'd14,8'd81} : s = 500;
	{8'd14,8'd82} : s = 65;
	{8'd14,8'd83} : s = 200;
	{8'd14,8'd84} : s = 196;
	{8'd14,8'd85} : s = 353;
	{8'd14,8'd86} : s = 194;
	{8'd14,8'd87} : s = 344;
	{8'd14,8'd88} : s = 340;
	{8'd14,8'd89} : s = 457;
	{8'd14,8'd90} : s = 193;
	{8'd14,8'd91} : s = 338;
	{8'd14,8'd92} : s = 337;
	{8'd14,8'd93} : s = 454;
	{8'd14,8'd94} : s = 332;
	{8'd14,8'd95} : s = 453;
	{8'd14,8'd96} : s = 451;
	{8'd14,8'd97} : s = 498;
	{8'd14,8'd98} : s = 176;
	{8'd14,8'd99} : s = 330;
	{8'd14,8'd100} : s = 329;
	{8'd14,8'd101} : s = 440;
	{8'd14,8'd102} : s = 326;
	{8'd14,8'd103} : s = 436;
	{8'd14,8'd104} : s = 434;
	{8'd14,8'd105} : s = 497;
	{8'd14,8'd106} : s = 325;
	{8'd14,8'd107} : s = 433;
	{8'd14,8'd108} : s = 428;
	{8'd14,8'd109} : s = 492;
	{8'd14,8'd110} : s = 426;
	{8'd14,8'd111} : s = 490;
	{8'd14,8'd112} : s = 489;
	{8'd14,8'd113} : s = 508;
	{8'd14,8'd114} : s = 2;
	{8'd14,8'd115} : s = 48;
	{8'd14,8'd116} : s = 40;
	{8'd14,8'd117} : s = 168;
	{8'd14,8'd118} : s = 36;
	{8'd14,8'd119} : s = 164;
	{8'd14,8'd120} : s = 162;
	{8'd14,8'd121} : s = 323;
	{8'd14,8'd122} : s = 34;
	{8'd14,8'd123} : s = 161;
	{8'd14,8'd124} : s = 152;
	{8'd14,8'd125} : s = 312;
	{8'd14,8'd126} : s = 148;
	{8'd14,8'd127} : s = 308;
	{8'd14,8'd128} : s = 306;
	{8'd14,8'd129} : s = 425;
	{8'd14,8'd130} : s = 33;
	{8'd14,8'd131} : s = 146;
	{8'd14,8'd132} : s = 145;
	{8'd14,8'd133} : s = 305;
	{8'd14,8'd134} : s = 140;
	{8'd14,8'd135} : s = 300;
	{8'd14,8'd136} : s = 298;
	{8'd14,8'd137} : s = 422;
	{8'd14,8'd138} : s = 138;
	{8'd14,8'd139} : s = 297;
	{8'd14,8'd140} : s = 294;
	{8'd14,8'd141} : s = 421;
	{8'd14,8'd142} : s = 293;
	{8'd14,8'd143} : s = 419;
	{8'd14,8'd144} : s = 412;
	{8'd14,8'd145} : s = 486;
	{8'd14,8'd146} : s = 24;
	{8'd14,8'd147} : s = 137;
	{8'd14,8'd148} : s = 134;
	{8'd14,8'd149} : s = 291;
	{8'd14,8'd150} : s = 133;
	{8'd14,8'd151} : s = 284;
	{8'd14,8'd152} : s = 282;
	{8'd14,8'd153} : s = 410;
	{8'd14,8'd154} : s = 131;
	{8'd14,8'd155} : s = 281;
	{8'd14,8'd156} : s = 278;
	{8'd14,8'd157} : s = 409;
	{8'd14,8'd158} : s = 277;
	{8'd14,8'd159} : s = 406;
	{8'd14,8'd160} : s = 405;
	{8'd14,8'd161} : s = 485;
	{8'd14,8'd162} : s = 112;
	{8'd14,8'd163} : s = 275;
	{8'd14,8'd164} : s = 270;
	{8'd14,8'd165} : s = 403;
	{8'd14,8'd166} : s = 269;
	{8'd14,8'd167} : s = 398;
	{8'd14,8'd168} : s = 397;
	{8'd14,8'd169} : s = 483;
	{8'd14,8'd170} : s = 267;
	{8'd14,8'd171} : s = 395;
	{8'd14,8'd172} : s = 391;
	{8'd14,8'd173} : s = 476;
	{8'd14,8'd174} : s = 376;
	{8'd14,8'd175} : s = 474;
	{8'd14,8'd176} : s = 473;
	{8'd14,8'd177} : s = 506;
	{8'd14,8'd178} : s = 20;
	{8'd14,8'd179} : s = 104;
	{8'd14,8'd180} : s = 100;
	{8'd14,8'd181} : s = 263;
	{8'd14,8'd182} : s = 98;
	{8'd14,8'd183} : s = 240;
	{8'd14,8'd184} : s = 232;
	{8'd14,8'd185} : s = 372;
	{8'd14,8'd186} : s = 97;
	{8'd14,8'd187} : s = 228;
	{8'd14,8'd188} : s = 226;
	{8'd14,8'd189} : s = 370;
	{8'd14,8'd190} : s = 225;
	{8'd14,8'd191} : s = 369;
	{8'd14,8'd192} : s = 364;
	{8'd14,8'd193} : s = 470;
	{8'd14,8'd194} : s = 88;
	{8'd14,8'd195} : s = 216;
	{8'd14,8'd196} : s = 212;
	{8'd14,8'd197} : s = 362;
	{8'd14,8'd198} : s = 210;
	{8'd14,8'd199} : s = 361;
	{8'd14,8'd200} : s = 358;
	{8'd14,8'd201} : s = 469;
	{8'd14,8'd202} : s = 209;
	{8'd14,8'd203} : s = 357;
	{8'd14,8'd204} : s = 355;
	{8'd14,8'd205} : s = 467;
	{8'd14,8'd206} : s = 348;
	{8'd14,8'd207} : s = 462;
	{8'd14,8'd208} : s = 461;
	{8'd14,8'd209} : s = 505;
	{8'd14,8'd210} : s = 84;
	{8'd14,8'd211} : s = 204;
	{8'd14,8'd212} : s = 202;
	{8'd14,8'd213} : s = 346;
	{8'd14,8'd214} : s = 201;
	{8'd14,8'd215} : s = 345;
	{8'd14,8'd216} : s = 342;
	{8'd14,8'd217} : s = 459;
	{8'd14,8'd218} : s = 198;
	{8'd14,8'd219} : s = 341;
	{8'd14,8'd220} : s = 339;
	{8'd14,8'd221} : s = 455;
	{8'd14,8'd222} : s = 334;
	{8'd14,8'd223} : s = 444;
	{8'd14,8'd224} : s = 442;
	{8'd14,8'd225} : s = 502;
	{8'd14,8'd226} : s = 197;
	{8'd14,8'd227} : s = 333;
	{8'd14,8'd228} : s = 331;
	{8'd14,8'd229} : s = 441;
	{8'd14,8'd230} : s = 327;
	{8'd14,8'd231} : s = 438;
	{8'd14,8'd232} : s = 437;
	{8'd14,8'd233} : s = 501;
	{8'd14,8'd234} : s = 316;
	{8'd14,8'd235} : s = 435;
	{8'd14,8'd236} : s = 430;
	{8'd14,8'd237} : s = 499;
	{8'd14,8'd238} : s = 429;
	{8'd14,8'd239} : s = 494;
	{8'd14,8'd240} : s = 493;
	{8'd14,8'd241} : s = 510;
	{8'd14,8'd242} : s = 1;
	{8'd14,8'd243} : s = 18;
	{8'd14,8'd244} : s = 17;
	{8'd14,8'd245} : s = 82;
	{8'd14,8'd246} : s = 12;
	{8'd14,8'd247} : s = 81;
	{8'd14,8'd248} : s = 76;
	{8'd14,8'd249} : s = 195;
	{8'd14,8'd250} : s = 10;
	{8'd14,8'd251} : s = 74;
	{8'd14,8'd252} : s = 73;
	{8'd14,8'd253} : s = 184;
	{8'd14,8'd254} : s = 70;
	{8'd14,8'd255} : s = 180;
	{8'd15,8'd0} : s = 480;
	{8'd15,8'd1} : s = 8;
	{8'd15,8'd2} : s = 258;
	{8'd15,8'd3} : s = 257;
	{8'd15,8'd4} : s = 388;
	{8'd15,8'd5} : s = 192;
	{8'd15,8'd6} : s = 386;
	{8'd15,8'd7} : s = 385;
	{8'd15,8'd8} : s = 464;
	{8'd15,8'd9} : s = 160;
	{8'd15,8'd10} : s = 352;
	{8'd15,8'd11} : s = 336;
	{8'd15,8'd12} : s = 456;
	{8'd15,8'd13} : s = 328;
	{8'd15,8'd14} : s = 452;
	{8'd15,8'd15} : s = 450;
	{8'd15,8'd16} : s = 496;
	{8'd15,8'd17} : s = 16;
	{8'd15,8'd18} : s = 144;
	{8'd15,8'd19} : s = 136;
	{8'd15,8'd20} : s = 324;
	{8'd15,8'd21} : s = 132;
	{8'd15,8'd22} : s = 322;
	{8'd15,8'd23} : s = 321;
	{8'd15,8'd24} : s = 449;
	{8'd15,8'd25} : s = 130;
	{8'd15,8'd26} : s = 304;
	{8'd15,8'd27} : s = 296;
	{8'd15,8'd28} : s = 432;
	{8'd15,8'd29} : s = 292;
	{8'd15,8'd30} : s = 424;
	{8'd15,8'd31} : s = 420;
	{8'd15,8'd32} : s = 488;
	{8'd15,8'd33} : s = 129;
	{8'd15,8'd34} : s = 290;
	{8'd15,8'd35} : s = 289;
	{8'd15,8'd36} : s = 418;
	{8'd15,8'd37} : s = 280;
	{8'd15,8'd38} : s = 417;
	{8'd15,8'd39} : s = 408;
	{8'd15,8'd40} : s = 484;
	{8'd15,8'd41} : s = 276;
	{8'd15,8'd42} : s = 404;
	{8'd15,8'd43} : s = 402;
	{8'd15,8'd44} : s = 482;
	{8'd15,8'd45} : s = 401;
	{8'd15,8'd46} : s = 481;
	{8'd15,8'd47} : s = 472;
	{8'd15,8'd48} : s = 504;
	{8'd15,8'd49} : s = 4;
	{8'd15,8'd50} : s = 96;
	{8'd15,8'd51} : s = 80;
	{8'd15,8'd52} : s = 274;
	{8'd15,8'd53} : s = 72;
	{8'd15,8'd54} : s = 273;
	{8'd15,8'd55} : s = 268;
	{8'd15,8'd56} : s = 396;
	{8'd15,8'd57} : s = 68;
	{8'd15,8'd58} : s = 266;
	{8'd15,8'd59} : s = 265;
	{8'd15,8'd60} : s = 394;
	{8'd15,8'd61} : s = 262;
	{8'd15,8'd62} : s = 393;
	{8'd15,8'd63} : s = 390;
	{8'd15,8'd64} : s = 468;
	{8'd15,8'd65} : s = 66;
	{8'd15,8'd66} : s = 261;
	{8'd15,8'd67} : s = 259;
	{8'd15,8'd68} : s = 389;
	{8'd15,8'd69} : s = 224;
	{8'd15,8'd70} : s = 387;
	{8'd15,8'd71} : s = 368;
	{8'd15,8'd72} : s = 466;
	{8'd15,8'd73} : s = 208;
	{8'd15,8'd74} : s = 360;
	{8'd15,8'd75} : s = 356;
	{8'd15,8'd76} : s = 465;
	{8'd15,8'd77} : s = 354;
	{8'd15,8'd78} : s = 460;
	{8'd15,8'd79} : s = 458;
	{8'd15,8'd80} : s = 500;
	{8'd15,8'd81} : s = 65;
	{8'd15,8'd82} : s = 200;
	{8'd15,8'd83} : s = 196;
	{8'd15,8'd84} : s = 353;
	{8'd15,8'd85} : s = 194;
	{8'd15,8'd86} : s = 344;
	{8'd15,8'd87} : s = 340;
	{8'd15,8'd88} : s = 457;
	{8'd15,8'd89} : s = 193;
	{8'd15,8'd90} : s = 338;
	{8'd15,8'd91} : s = 337;
	{8'd15,8'd92} : s = 454;
	{8'd15,8'd93} : s = 332;
	{8'd15,8'd94} : s = 453;
	{8'd15,8'd95} : s = 451;
	{8'd15,8'd96} : s = 498;
	{8'd15,8'd97} : s = 176;
	{8'd15,8'd98} : s = 330;
	{8'd15,8'd99} : s = 329;
	{8'd15,8'd100} : s = 440;
	{8'd15,8'd101} : s = 326;
	{8'd15,8'd102} : s = 436;
	{8'd15,8'd103} : s = 434;
	{8'd15,8'd104} : s = 497;
	{8'd15,8'd105} : s = 325;
	{8'd15,8'd106} : s = 433;
	{8'd15,8'd107} : s = 428;
	{8'd15,8'd108} : s = 492;
	{8'd15,8'd109} : s = 426;
	{8'd15,8'd110} : s = 490;
	{8'd15,8'd111} : s = 489;
	{8'd15,8'd112} : s = 508;
	{8'd15,8'd113} : s = 2;
	{8'd15,8'd114} : s = 48;
	{8'd15,8'd115} : s = 40;
	{8'd15,8'd116} : s = 168;
	{8'd15,8'd117} : s = 36;
	{8'd15,8'd118} : s = 164;
	{8'd15,8'd119} : s = 162;
	{8'd15,8'd120} : s = 323;
	{8'd15,8'd121} : s = 34;
	{8'd15,8'd122} : s = 161;
	{8'd15,8'd123} : s = 152;
	{8'd15,8'd124} : s = 312;
	{8'd15,8'd125} : s = 148;
	{8'd15,8'd126} : s = 308;
	{8'd15,8'd127} : s = 306;
	{8'd15,8'd128} : s = 425;
	{8'd15,8'd129} : s = 33;
	{8'd15,8'd130} : s = 146;
	{8'd15,8'd131} : s = 145;
	{8'd15,8'd132} : s = 305;
	{8'd15,8'd133} : s = 140;
	{8'd15,8'd134} : s = 300;
	{8'd15,8'd135} : s = 298;
	{8'd15,8'd136} : s = 422;
	{8'd15,8'd137} : s = 138;
	{8'd15,8'd138} : s = 297;
	{8'd15,8'd139} : s = 294;
	{8'd15,8'd140} : s = 421;
	{8'd15,8'd141} : s = 293;
	{8'd15,8'd142} : s = 419;
	{8'd15,8'd143} : s = 412;
	{8'd15,8'd144} : s = 486;
	{8'd15,8'd145} : s = 24;
	{8'd15,8'd146} : s = 137;
	{8'd15,8'd147} : s = 134;
	{8'd15,8'd148} : s = 291;
	{8'd15,8'd149} : s = 133;
	{8'd15,8'd150} : s = 284;
	{8'd15,8'd151} : s = 282;
	{8'd15,8'd152} : s = 410;
	{8'd15,8'd153} : s = 131;
	{8'd15,8'd154} : s = 281;
	{8'd15,8'd155} : s = 278;
	{8'd15,8'd156} : s = 409;
	{8'd15,8'd157} : s = 277;
	{8'd15,8'd158} : s = 406;
	{8'd15,8'd159} : s = 405;
	{8'd15,8'd160} : s = 485;
	{8'd15,8'd161} : s = 112;
	{8'd15,8'd162} : s = 275;
	{8'd15,8'd163} : s = 270;
	{8'd15,8'd164} : s = 403;
	{8'd15,8'd165} : s = 269;
	{8'd15,8'd166} : s = 398;
	{8'd15,8'd167} : s = 397;
	{8'd15,8'd168} : s = 483;
	{8'd15,8'd169} : s = 267;
	{8'd15,8'd170} : s = 395;
	{8'd15,8'd171} : s = 391;
	{8'd15,8'd172} : s = 476;
	{8'd15,8'd173} : s = 376;
	{8'd15,8'd174} : s = 474;
	{8'd15,8'd175} : s = 473;
	{8'd15,8'd176} : s = 506;
	{8'd15,8'd177} : s = 20;
	{8'd15,8'd178} : s = 104;
	{8'd15,8'd179} : s = 100;
	{8'd15,8'd180} : s = 263;
	{8'd15,8'd181} : s = 98;
	{8'd15,8'd182} : s = 240;
	{8'd15,8'd183} : s = 232;
	{8'd15,8'd184} : s = 372;
	{8'd15,8'd185} : s = 97;
	{8'd15,8'd186} : s = 228;
	{8'd15,8'd187} : s = 226;
	{8'd15,8'd188} : s = 370;
	{8'd15,8'd189} : s = 225;
	{8'd15,8'd190} : s = 369;
	{8'd15,8'd191} : s = 364;
	{8'd15,8'd192} : s = 470;
	{8'd15,8'd193} : s = 88;
	{8'd15,8'd194} : s = 216;
	{8'd15,8'd195} : s = 212;
	{8'd15,8'd196} : s = 362;
	{8'd15,8'd197} : s = 210;
	{8'd15,8'd198} : s = 361;
	{8'd15,8'd199} : s = 358;
	{8'd15,8'd200} : s = 469;
	{8'd15,8'd201} : s = 209;
	{8'd15,8'd202} : s = 357;
	{8'd15,8'd203} : s = 355;
	{8'd15,8'd204} : s = 467;
	{8'd15,8'd205} : s = 348;
	{8'd15,8'd206} : s = 462;
	{8'd15,8'd207} : s = 461;
	{8'd15,8'd208} : s = 505;
	{8'd15,8'd209} : s = 84;
	{8'd15,8'd210} : s = 204;
	{8'd15,8'd211} : s = 202;
	{8'd15,8'd212} : s = 346;
	{8'd15,8'd213} : s = 201;
	{8'd15,8'd214} : s = 345;
	{8'd15,8'd215} : s = 342;
	{8'd15,8'd216} : s = 459;
	{8'd15,8'd217} : s = 198;
	{8'd15,8'd218} : s = 341;
	{8'd15,8'd219} : s = 339;
	{8'd15,8'd220} : s = 455;
	{8'd15,8'd221} : s = 334;
	{8'd15,8'd222} : s = 444;
	{8'd15,8'd223} : s = 442;
	{8'd15,8'd224} : s = 502;
	{8'd15,8'd225} : s = 197;
	{8'd15,8'd226} : s = 333;
	{8'd15,8'd227} : s = 331;
	{8'd15,8'd228} : s = 441;
	{8'd15,8'd229} : s = 327;
	{8'd15,8'd230} : s = 438;
	{8'd15,8'd231} : s = 437;
	{8'd15,8'd232} : s = 501;
	{8'd15,8'd233} : s = 316;
	{8'd15,8'd234} : s = 435;
	{8'd15,8'd235} : s = 430;
	{8'd15,8'd236} : s = 499;
	{8'd15,8'd237} : s = 429;
	{8'd15,8'd238} : s = 494;
	{8'd15,8'd239} : s = 493;
	{8'd15,8'd240} : s = 510;
	{8'd15,8'd241} : s = 1;
	{8'd15,8'd242} : s = 18;
	{8'd15,8'd243} : s = 17;
	{8'd15,8'd244} : s = 82;
	{8'd15,8'd245} : s = 12;
	{8'd15,8'd246} : s = 81;
	{8'd15,8'd247} : s = 76;
	{8'd15,8'd248} : s = 195;
	{8'd15,8'd249} : s = 10;
	{8'd15,8'd250} : s = 74;
	{8'd15,8'd251} : s = 73;
	{8'd15,8'd252} : s = 184;
	{8'd15,8'd253} : s = 70;
	{8'd15,8'd254} : s = 180;
	{8'd15,8'd255} : s = 178;
	{8'd16,8'd0} : s = 8;
	{8'd16,8'd1} : s = 258;
	{8'd16,8'd2} : s = 257;
	{8'd16,8'd3} : s = 388;
	{8'd16,8'd4} : s = 192;
	{8'd16,8'd5} : s = 386;
	{8'd16,8'd6} : s = 385;
	{8'd16,8'd7} : s = 464;
	{8'd16,8'd8} : s = 160;
	{8'd16,8'd9} : s = 352;
	{8'd16,8'd10} : s = 336;
	{8'd16,8'd11} : s = 456;
	{8'd16,8'd12} : s = 328;
	{8'd16,8'd13} : s = 452;
	{8'd16,8'd14} : s = 450;
	{8'd16,8'd15} : s = 496;
	{8'd16,8'd16} : s = 16;
	{8'd16,8'd17} : s = 144;
	{8'd16,8'd18} : s = 136;
	{8'd16,8'd19} : s = 324;
	{8'd16,8'd20} : s = 132;
	{8'd16,8'd21} : s = 322;
	{8'd16,8'd22} : s = 321;
	{8'd16,8'd23} : s = 449;
	{8'd16,8'd24} : s = 130;
	{8'd16,8'd25} : s = 304;
	{8'd16,8'd26} : s = 296;
	{8'd16,8'd27} : s = 432;
	{8'd16,8'd28} : s = 292;
	{8'd16,8'd29} : s = 424;
	{8'd16,8'd30} : s = 420;
	{8'd16,8'd31} : s = 488;
	{8'd16,8'd32} : s = 129;
	{8'd16,8'd33} : s = 290;
	{8'd16,8'd34} : s = 289;
	{8'd16,8'd35} : s = 418;
	{8'd16,8'd36} : s = 280;
	{8'd16,8'd37} : s = 417;
	{8'd16,8'd38} : s = 408;
	{8'd16,8'd39} : s = 484;
	{8'd16,8'd40} : s = 276;
	{8'd16,8'd41} : s = 404;
	{8'd16,8'd42} : s = 402;
	{8'd16,8'd43} : s = 482;
	{8'd16,8'd44} : s = 401;
	{8'd16,8'd45} : s = 481;
	{8'd16,8'd46} : s = 472;
	{8'd16,8'd47} : s = 504;
	{8'd16,8'd48} : s = 4;
	{8'd16,8'd49} : s = 96;
	{8'd16,8'd50} : s = 80;
	{8'd16,8'd51} : s = 274;
	{8'd16,8'd52} : s = 72;
	{8'd16,8'd53} : s = 273;
	{8'd16,8'd54} : s = 268;
	{8'd16,8'd55} : s = 396;
	{8'd16,8'd56} : s = 68;
	{8'd16,8'd57} : s = 266;
	{8'd16,8'd58} : s = 265;
	{8'd16,8'd59} : s = 394;
	{8'd16,8'd60} : s = 262;
	{8'd16,8'd61} : s = 393;
	{8'd16,8'd62} : s = 390;
	{8'd16,8'd63} : s = 468;
	{8'd16,8'd64} : s = 66;
	{8'd16,8'd65} : s = 261;
	{8'd16,8'd66} : s = 259;
	{8'd16,8'd67} : s = 389;
	{8'd16,8'd68} : s = 224;
	{8'd16,8'd69} : s = 387;
	{8'd16,8'd70} : s = 368;
	{8'd16,8'd71} : s = 466;
	{8'd16,8'd72} : s = 208;
	{8'd16,8'd73} : s = 360;
	{8'd16,8'd74} : s = 356;
	{8'd16,8'd75} : s = 465;
	{8'd16,8'd76} : s = 354;
	{8'd16,8'd77} : s = 460;
	{8'd16,8'd78} : s = 458;
	{8'd16,8'd79} : s = 500;
	{8'd16,8'd80} : s = 65;
	{8'd16,8'd81} : s = 200;
	{8'd16,8'd82} : s = 196;
	{8'd16,8'd83} : s = 353;
	{8'd16,8'd84} : s = 194;
	{8'd16,8'd85} : s = 344;
	{8'd16,8'd86} : s = 340;
	{8'd16,8'd87} : s = 457;
	{8'd16,8'd88} : s = 193;
	{8'd16,8'd89} : s = 338;
	{8'd16,8'd90} : s = 337;
	{8'd16,8'd91} : s = 454;
	{8'd16,8'd92} : s = 332;
	{8'd16,8'd93} : s = 453;
	{8'd16,8'd94} : s = 451;
	{8'd16,8'd95} : s = 498;
	{8'd16,8'd96} : s = 176;
	{8'd16,8'd97} : s = 330;
	{8'd16,8'd98} : s = 329;
	{8'd16,8'd99} : s = 440;
	{8'd16,8'd100} : s = 326;
	{8'd16,8'd101} : s = 436;
	{8'd16,8'd102} : s = 434;
	{8'd16,8'd103} : s = 497;
	{8'd16,8'd104} : s = 325;
	{8'd16,8'd105} : s = 433;
	{8'd16,8'd106} : s = 428;
	{8'd16,8'd107} : s = 492;
	{8'd16,8'd108} : s = 426;
	{8'd16,8'd109} : s = 490;
	{8'd16,8'd110} : s = 489;
	{8'd16,8'd111} : s = 508;
	{8'd16,8'd112} : s = 2;
	{8'd16,8'd113} : s = 48;
	{8'd16,8'd114} : s = 40;
	{8'd16,8'd115} : s = 168;
	{8'd16,8'd116} : s = 36;
	{8'd16,8'd117} : s = 164;
	{8'd16,8'd118} : s = 162;
	{8'd16,8'd119} : s = 323;
	{8'd16,8'd120} : s = 34;
	{8'd16,8'd121} : s = 161;
	{8'd16,8'd122} : s = 152;
	{8'd16,8'd123} : s = 312;
	{8'd16,8'd124} : s = 148;
	{8'd16,8'd125} : s = 308;
	{8'd16,8'd126} : s = 306;
	{8'd16,8'd127} : s = 425;
	{8'd16,8'd128} : s = 33;
	{8'd16,8'd129} : s = 146;
	{8'd16,8'd130} : s = 145;
	{8'd16,8'd131} : s = 305;
	{8'd16,8'd132} : s = 140;
	{8'd16,8'd133} : s = 300;
	{8'd16,8'd134} : s = 298;
	{8'd16,8'd135} : s = 422;
	{8'd16,8'd136} : s = 138;
	{8'd16,8'd137} : s = 297;
	{8'd16,8'd138} : s = 294;
	{8'd16,8'd139} : s = 421;
	{8'd16,8'd140} : s = 293;
	{8'd16,8'd141} : s = 419;
	{8'd16,8'd142} : s = 412;
	{8'd16,8'd143} : s = 486;
	{8'd16,8'd144} : s = 24;
	{8'd16,8'd145} : s = 137;
	{8'd16,8'd146} : s = 134;
	{8'd16,8'd147} : s = 291;
	{8'd16,8'd148} : s = 133;
	{8'd16,8'd149} : s = 284;
	{8'd16,8'd150} : s = 282;
	{8'd16,8'd151} : s = 410;
	{8'd16,8'd152} : s = 131;
	{8'd16,8'd153} : s = 281;
	{8'd16,8'd154} : s = 278;
	{8'd16,8'd155} : s = 409;
	{8'd16,8'd156} : s = 277;
	{8'd16,8'd157} : s = 406;
	{8'd16,8'd158} : s = 405;
	{8'd16,8'd159} : s = 485;
	{8'd16,8'd160} : s = 112;
	{8'd16,8'd161} : s = 275;
	{8'd16,8'd162} : s = 270;
	{8'd16,8'd163} : s = 403;
	{8'd16,8'd164} : s = 269;
	{8'd16,8'd165} : s = 398;
	{8'd16,8'd166} : s = 397;
	{8'd16,8'd167} : s = 483;
	{8'd16,8'd168} : s = 267;
	{8'd16,8'd169} : s = 395;
	{8'd16,8'd170} : s = 391;
	{8'd16,8'd171} : s = 476;
	{8'd16,8'd172} : s = 376;
	{8'd16,8'd173} : s = 474;
	{8'd16,8'd174} : s = 473;
	{8'd16,8'd175} : s = 506;
	{8'd16,8'd176} : s = 20;
	{8'd16,8'd177} : s = 104;
	{8'd16,8'd178} : s = 100;
	{8'd16,8'd179} : s = 263;
	{8'd16,8'd180} : s = 98;
	{8'd16,8'd181} : s = 240;
	{8'd16,8'd182} : s = 232;
	{8'd16,8'd183} : s = 372;
	{8'd16,8'd184} : s = 97;
	{8'd16,8'd185} : s = 228;
	{8'd16,8'd186} : s = 226;
	{8'd16,8'd187} : s = 370;
	{8'd16,8'd188} : s = 225;
	{8'd16,8'd189} : s = 369;
	{8'd16,8'd190} : s = 364;
	{8'd16,8'd191} : s = 470;
	{8'd16,8'd192} : s = 88;
	{8'd16,8'd193} : s = 216;
	{8'd16,8'd194} : s = 212;
	{8'd16,8'd195} : s = 362;
	{8'd16,8'd196} : s = 210;
	{8'd16,8'd197} : s = 361;
	{8'd16,8'd198} : s = 358;
	{8'd16,8'd199} : s = 469;
	{8'd16,8'd200} : s = 209;
	{8'd16,8'd201} : s = 357;
	{8'd16,8'd202} : s = 355;
	{8'd16,8'd203} : s = 467;
	{8'd16,8'd204} : s = 348;
	{8'd16,8'd205} : s = 462;
	{8'd16,8'd206} : s = 461;
	{8'd16,8'd207} : s = 505;
	{8'd16,8'd208} : s = 84;
	{8'd16,8'd209} : s = 204;
	{8'd16,8'd210} : s = 202;
	{8'd16,8'd211} : s = 346;
	{8'd16,8'd212} : s = 201;
	{8'd16,8'd213} : s = 345;
	{8'd16,8'd214} : s = 342;
	{8'd16,8'd215} : s = 459;
	{8'd16,8'd216} : s = 198;
	{8'd16,8'd217} : s = 341;
	{8'd16,8'd218} : s = 339;
	{8'd16,8'd219} : s = 455;
	{8'd16,8'd220} : s = 334;
	{8'd16,8'd221} : s = 444;
	{8'd16,8'd222} : s = 442;
	{8'd16,8'd223} : s = 502;
	{8'd16,8'd224} : s = 197;
	{8'd16,8'd225} : s = 333;
	{8'd16,8'd226} : s = 331;
	{8'd16,8'd227} : s = 441;
	{8'd16,8'd228} : s = 327;
	{8'd16,8'd229} : s = 438;
	{8'd16,8'd230} : s = 437;
	{8'd16,8'd231} : s = 501;
	{8'd16,8'd232} : s = 316;
	{8'd16,8'd233} : s = 435;
	{8'd16,8'd234} : s = 430;
	{8'd16,8'd235} : s = 499;
	{8'd16,8'd236} : s = 429;
	{8'd16,8'd237} : s = 494;
	{8'd16,8'd238} : s = 493;
	{8'd16,8'd239} : s = 510;
	{8'd16,8'd240} : s = 1;
	{8'd16,8'd241} : s = 18;
	{8'd16,8'd242} : s = 17;
	{8'd16,8'd243} : s = 82;
	{8'd16,8'd244} : s = 12;
	{8'd16,8'd245} : s = 81;
	{8'd16,8'd246} : s = 76;
	{8'd16,8'd247} : s = 195;
	{8'd16,8'd248} : s = 10;
	{8'd16,8'd249} : s = 74;
	{8'd16,8'd250} : s = 73;
	{8'd16,8'd251} : s = 184;
	{8'd16,8'd252} : s = 70;
	{8'd16,8'd253} : s = 180;
	{8'd16,8'd254} : s = 178;
	{8'd16,8'd255} : s = 314;
	{8'd17,8'd0} : s = 258;
	{8'd17,8'd1} : s = 257;
	{8'd17,8'd2} : s = 388;
	{8'd17,8'd3} : s = 192;
	{8'd17,8'd4} : s = 386;
	{8'd17,8'd5} : s = 385;
	{8'd17,8'd6} : s = 464;
	{8'd17,8'd7} : s = 160;
	{8'd17,8'd8} : s = 352;
	{8'd17,8'd9} : s = 336;
	{8'd17,8'd10} : s = 456;
	{8'd17,8'd11} : s = 328;
	{8'd17,8'd12} : s = 452;
	{8'd17,8'd13} : s = 450;
	{8'd17,8'd14} : s = 496;
	{8'd17,8'd15} : s = 16;
	{8'd17,8'd16} : s = 144;
	{8'd17,8'd17} : s = 136;
	{8'd17,8'd18} : s = 324;
	{8'd17,8'd19} : s = 132;
	{8'd17,8'd20} : s = 322;
	{8'd17,8'd21} : s = 321;
	{8'd17,8'd22} : s = 449;
	{8'd17,8'd23} : s = 130;
	{8'd17,8'd24} : s = 304;
	{8'd17,8'd25} : s = 296;
	{8'd17,8'd26} : s = 432;
	{8'd17,8'd27} : s = 292;
	{8'd17,8'd28} : s = 424;
	{8'd17,8'd29} : s = 420;
	{8'd17,8'd30} : s = 488;
	{8'd17,8'd31} : s = 129;
	{8'd17,8'd32} : s = 290;
	{8'd17,8'd33} : s = 289;
	{8'd17,8'd34} : s = 418;
	{8'd17,8'd35} : s = 280;
	{8'd17,8'd36} : s = 417;
	{8'd17,8'd37} : s = 408;
	{8'd17,8'd38} : s = 484;
	{8'd17,8'd39} : s = 276;
	{8'd17,8'd40} : s = 404;
	{8'd17,8'd41} : s = 402;
	{8'd17,8'd42} : s = 482;
	{8'd17,8'd43} : s = 401;
	{8'd17,8'd44} : s = 481;
	{8'd17,8'd45} : s = 472;
	{8'd17,8'd46} : s = 504;
	{8'd17,8'd47} : s = 4;
	{8'd17,8'd48} : s = 96;
	{8'd17,8'd49} : s = 80;
	{8'd17,8'd50} : s = 274;
	{8'd17,8'd51} : s = 72;
	{8'd17,8'd52} : s = 273;
	{8'd17,8'd53} : s = 268;
	{8'd17,8'd54} : s = 396;
	{8'd17,8'd55} : s = 68;
	{8'd17,8'd56} : s = 266;
	{8'd17,8'd57} : s = 265;
	{8'd17,8'd58} : s = 394;
	{8'd17,8'd59} : s = 262;
	{8'd17,8'd60} : s = 393;
	{8'd17,8'd61} : s = 390;
	{8'd17,8'd62} : s = 468;
	{8'd17,8'd63} : s = 66;
	{8'd17,8'd64} : s = 261;
	{8'd17,8'd65} : s = 259;
	{8'd17,8'd66} : s = 389;
	{8'd17,8'd67} : s = 224;
	{8'd17,8'd68} : s = 387;
	{8'd17,8'd69} : s = 368;
	{8'd17,8'd70} : s = 466;
	{8'd17,8'd71} : s = 208;
	{8'd17,8'd72} : s = 360;
	{8'd17,8'd73} : s = 356;
	{8'd17,8'd74} : s = 465;
	{8'd17,8'd75} : s = 354;
	{8'd17,8'd76} : s = 460;
	{8'd17,8'd77} : s = 458;
	{8'd17,8'd78} : s = 500;
	{8'd17,8'd79} : s = 65;
	{8'd17,8'd80} : s = 200;
	{8'd17,8'd81} : s = 196;
	{8'd17,8'd82} : s = 353;
	{8'd17,8'd83} : s = 194;
	{8'd17,8'd84} : s = 344;
	{8'd17,8'd85} : s = 340;
	{8'd17,8'd86} : s = 457;
	{8'd17,8'd87} : s = 193;
	{8'd17,8'd88} : s = 338;
	{8'd17,8'd89} : s = 337;
	{8'd17,8'd90} : s = 454;
	{8'd17,8'd91} : s = 332;
	{8'd17,8'd92} : s = 453;
	{8'd17,8'd93} : s = 451;
	{8'd17,8'd94} : s = 498;
	{8'd17,8'd95} : s = 176;
	{8'd17,8'd96} : s = 330;
	{8'd17,8'd97} : s = 329;
	{8'd17,8'd98} : s = 440;
	{8'd17,8'd99} : s = 326;
	{8'd17,8'd100} : s = 436;
	{8'd17,8'd101} : s = 434;
	{8'd17,8'd102} : s = 497;
	{8'd17,8'd103} : s = 325;
	{8'd17,8'd104} : s = 433;
	{8'd17,8'd105} : s = 428;
	{8'd17,8'd106} : s = 492;
	{8'd17,8'd107} : s = 426;
	{8'd17,8'd108} : s = 490;
	{8'd17,8'd109} : s = 489;
	{8'd17,8'd110} : s = 508;
	{8'd17,8'd111} : s = 2;
	{8'd17,8'd112} : s = 48;
	{8'd17,8'd113} : s = 40;
	{8'd17,8'd114} : s = 168;
	{8'd17,8'd115} : s = 36;
	{8'd17,8'd116} : s = 164;
	{8'd17,8'd117} : s = 162;
	{8'd17,8'd118} : s = 323;
	{8'd17,8'd119} : s = 34;
	{8'd17,8'd120} : s = 161;
	{8'd17,8'd121} : s = 152;
	{8'd17,8'd122} : s = 312;
	{8'd17,8'd123} : s = 148;
	{8'd17,8'd124} : s = 308;
	{8'd17,8'd125} : s = 306;
	{8'd17,8'd126} : s = 425;
	{8'd17,8'd127} : s = 33;
	{8'd17,8'd128} : s = 146;
	{8'd17,8'd129} : s = 145;
	{8'd17,8'd130} : s = 305;
	{8'd17,8'd131} : s = 140;
	{8'd17,8'd132} : s = 300;
	{8'd17,8'd133} : s = 298;
	{8'd17,8'd134} : s = 422;
	{8'd17,8'd135} : s = 138;
	{8'd17,8'd136} : s = 297;
	{8'd17,8'd137} : s = 294;
	{8'd17,8'd138} : s = 421;
	{8'd17,8'd139} : s = 293;
	{8'd17,8'd140} : s = 419;
	{8'd17,8'd141} : s = 412;
	{8'd17,8'd142} : s = 486;
	{8'd17,8'd143} : s = 24;
	{8'd17,8'd144} : s = 137;
	{8'd17,8'd145} : s = 134;
	{8'd17,8'd146} : s = 291;
	{8'd17,8'd147} : s = 133;
	{8'd17,8'd148} : s = 284;
	{8'd17,8'd149} : s = 282;
	{8'd17,8'd150} : s = 410;
	{8'd17,8'd151} : s = 131;
	{8'd17,8'd152} : s = 281;
	{8'd17,8'd153} : s = 278;
	{8'd17,8'd154} : s = 409;
	{8'd17,8'd155} : s = 277;
	{8'd17,8'd156} : s = 406;
	{8'd17,8'd157} : s = 405;
	{8'd17,8'd158} : s = 485;
	{8'd17,8'd159} : s = 112;
	{8'd17,8'd160} : s = 275;
	{8'd17,8'd161} : s = 270;
	{8'd17,8'd162} : s = 403;
	{8'd17,8'd163} : s = 269;
	{8'd17,8'd164} : s = 398;
	{8'd17,8'd165} : s = 397;
	{8'd17,8'd166} : s = 483;
	{8'd17,8'd167} : s = 267;
	{8'd17,8'd168} : s = 395;
	{8'd17,8'd169} : s = 391;
	{8'd17,8'd170} : s = 476;
	{8'd17,8'd171} : s = 376;
	{8'd17,8'd172} : s = 474;
	{8'd17,8'd173} : s = 473;
	{8'd17,8'd174} : s = 506;
	{8'd17,8'd175} : s = 20;
	{8'd17,8'd176} : s = 104;
	{8'd17,8'd177} : s = 100;
	{8'd17,8'd178} : s = 263;
	{8'd17,8'd179} : s = 98;
	{8'd17,8'd180} : s = 240;
	{8'd17,8'd181} : s = 232;
	{8'd17,8'd182} : s = 372;
	{8'd17,8'd183} : s = 97;
	{8'd17,8'd184} : s = 228;
	{8'd17,8'd185} : s = 226;
	{8'd17,8'd186} : s = 370;
	{8'd17,8'd187} : s = 225;
	{8'd17,8'd188} : s = 369;
	{8'd17,8'd189} : s = 364;
	{8'd17,8'd190} : s = 470;
	{8'd17,8'd191} : s = 88;
	{8'd17,8'd192} : s = 216;
	{8'd17,8'd193} : s = 212;
	{8'd17,8'd194} : s = 362;
	{8'd17,8'd195} : s = 210;
	{8'd17,8'd196} : s = 361;
	{8'd17,8'd197} : s = 358;
	{8'd17,8'd198} : s = 469;
	{8'd17,8'd199} : s = 209;
	{8'd17,8'd200} : s = 357;
	{8'd17,8'd201} : s = 355;
	{8'd17,8'd202} : s = 467;
	{8'd17,8'd203} : s = 348;
	{8'd17,8'd204} : s = 462;
	{8'd17,8'd205} : s = 461;
	{8'd17,8'd206} : s = 505;
	{8'd17,8'd207} : s = 84;
	{8'd17,8'd208} : s = 204;
	{8'd17,8'd209} : s = 202;
	{8'd17,8'd210} : s = 346;
	{8'd17,8'd211} : s = 201;
	{8'd17,8'd212} : s = 345;
	{8'd17,8'd213} : s = 342;
	{8'd17,8'd214} : s = 459;
	{8'd17,8'd215} : s = 198;
	{8'd17,8'd216} : s = 341;
	{8'd17,8'd217} : s = 339;
	{8'd17,8'd218} : s = 455;
	{8'd17,8'd219} : s = 334;
	{8'd17,8'd220} : s = 444;
	{8'd17,8'd221} : s = 442;
	{8'd17,8'd222} : s = 502;
	{8'd17,8'd223} : s = 197;
	{8'd17,8'd224} : s = 333;
	{8'd17,8'd225} : s = 331;
	{8'd17,8'd226} : s = 441;
	{8'd17,8'd227} : s = 327;
	{8'd17,8'd228} : s = 438;
	{8'd17,8'd229} : s = 437;
	{8'd17,8'd230} : s = 501;
	{8'd17,8'd231} : s = 316;
	{8'd17,8'd232} : s = 435;
	{8'd17,8'd233} : s = 430;
	{8'd17,8'd234} : s = 499;
	{8'd17,8'd235} : s = 429;
	{8'd17,8'd236} : s = 494;
	{8'd17,8'd237} : s = 493;
	{8'd17,8'd238} : s = 510;
	{8'd17,8'd239} : s = 1;
	{8'd17,8'd240} : s = 18;
	{8'd17,8'd241} : s = 17;
	{8'd17,8'd242} : s = 82;
	{8'd17,8'd243} : s = 12;
	{8'd17,8'd244} : s = 81;
	{8'd17,8'd245} : s = 76;
	{8'd17,8'd246} : s = 195;
	{8'd17,8'd247} : s = 10;
	{8'd17,8'd248} : s = 74;
	{8'd17,8'd249} : s = 73;
	{8'd17,8'd250} : s = 184;
	{8'd17,8'd251} : s = 70;
	{8'd17,8'd252} : s = 180;
	{8'd17,8'd253} : s = 178;
	{8'd17,8'd254} : s = 314;
	{8'd17,8'd255} : s = 9;
	{8'd18,8'd0} : s = 257;
	{8'd18,8'd1} : s = 388;
	{8'd18,8'd2} : s = 192;
	{8'd18,8'd3} : s = 386;
	{8'd18,8'd4} : s = 385;
	{8'd18,8'd5} : s = 464;
	{8'd18,8'd6} : s = 160;
	{8'd18,8'd7} : s = 352;
	{8'd18,8'd8} : s = 336;
	{8'd18,8'd9} : s = 456;
	{8'd18,8'd10} : s = 328;
	{8'd18,8'd11} : s = 452;
	{8'd18,8'd12} : s = 450;
	{8'd18,8'd13} : s = 496;
	{8'd18,8'd14} : s = 16;
	{8'd18,8'd15} : s = 144;
	{8'd18,8'd16} : s = 136;
	{8'd18,8'd17} : s = 324;
	{8'd18,8'd18} : s = 132;
	{8'd18,8'd19} : s = 322;
	{8'd18,8'd20} : s = 321;
	{8'd18,8'd21} : s = 449;
	{8'd18,8'd22} : s = 130;
	{8'd18,8'd23} : s = 304;
	{8'd18,8'd24} : s = 296;
	{8'd18,8'd25} : s = 432;
	{8'd18,8'd26} : s = 292;
	{8'd18,8'd27} : s = 424;
	{8'd18,8'd28} : s = 420;
	{8'd18,8'd29} : s = 488;
	{8'd18,8'd30} : s = 129;
	{8'd18,8'd31} : s = 290;
	{8'd18,8'd32} : s = 289;
	{8'd18,8'd33} : s = 418;
	{8'd18,8'd34} : s = 280;
	{8'd18,8'd35} : s = 417;
	{8'd18,8'd36} : s = 408;
	{8'd18,8'd37} : s = 484;
	{8'd18,8'd38} : s = 276;
	{8'd18,8'd39} : s = 404;
	{8'd18,8'd40} : s = 402;
	{8'd18,8'd41} : s = 482;
	{8'd18,8'd42} : s = 401;
	{8'd18,8'd43} : s = 481;
	{8'd18,8'd44} : s = 472;
	{8'd18,8'd45} : s = 504;
	{8'd18,8'd46} : s = 4;
	{8'd18,8'd47} : s = 96;
	{8'd18,8'd48} : s = 80;
	{8'd18,8'd49} : s = 274;
	{8'd18,8'd50} : s = 72;
	{8'd18,8'd51} : s = 273;
	{8'd18,8'd52} : s = 268;
	{8'd18,8'd53} : s = 396;
	{8'd18,8'd54} : s = 68;
	{8'd18,8'd55} : s = 266;
	{8'd18,8'd56} : s = 265;
	{8'd18,8'd57} : s = 394;
	{8'd18,8'd58} : s = 262;
	{8'd18,8'd59} : s = 393;
	{8'd18,8'd60} : s = 390;
	{8'd18,8'd61} : s = 468;
	{8'd18,8'd62} : s = 66;
	{8'd18,8'd63} : s = 261;
	{8'd18,8'd64} : s = 259;
	{8'd18,8'd65} : s = 389;
	{8'd18,8'd66} : s = 224;
	{8'd18,8'd67} : s = 387;
	{8'd18,8'd68} : s = 368;
	{8'd18,8'd69} : s = 466;
	{8'd18,8'd70} : s = 208;
	{8'd18,8'd71} : s = 360;
	{8'd18,8'd72} : s = 356;
	{8'd18,8'd73} : s = 465;
	{8'd18,8'd74} : s = 354;
	{8'd18,8'd75} : s = 460;
	{8'd18,8'd76} : s = 458;
	{8'd18,8'd77} : s = 500;
	{8'd18,8'd78} : s = 65;
	{8'd18,8'd79} : s = 200;
	{8'd18,8'd80} : s = 196;
	{8'd18,8'd81} : s = 353;
	{8'd18,8'd82} : s = 194;
	{8'd18,8'd83} : s = 344;
	{8'd18,8'd84} : s = 340;
	{8'd18,8'd85} : s = 457;
	{8'd18,8'd86} : s = 193;
	{8'd18,8'd87} : s = 338;
	{8'd18,8'd88} : s = 337;
	{8'd18,8'd89} : s = 454;
	{8'd18,8'd90} : s = 332;
	{8'd18,8'd91} : s = 453;
	{8'd18,8'd92} : s = 451;
	{8'd18,8'd93} : s = 498;
	{8'd18,8'd94} : s = 176;
	{8'd18,8'd95} : s = 330;
	{8'd18,8'd96} : s = 329;
	{8'd18,8'd97} : s = 440;
	{8'd18,8'd98} : s = 326;
	{8'd18,8'd99} : s = 436;
	{8'd18,8'd100} : s = 434;
	{8'd18,8'd101} : s = 497;
	{8'd18,8'd102} : s = 325;
	{8'd18,8'd103} : s = 433;
	{8'd18,8'd104} : s = 428;
	{8'd18,8'd105} : s = 492;
	{8'd18,8'd106} : s = 426;
	{8'd18,8'd107} : s = 490;
	{8'd18,8'd108} : s = 489;
	{8'd18,8'd109} : s = 508;
	{8'd18,8'd110} : s = 2;
	{8'd18,8'd111} : s = 48;
	{8'd18,8'd112} : s = 40;
	{8'd18,8'd113} : s = 168;
	{8'd18,8'd114} : s = 36;
	{8'd18,8'd115} : s = 164;
	{8'd18,8'd116} : s = 162;
	{8'd18,8'd117} : s = 323;
	{8'd18,8'd118} : s = 34;
	{8'd18,8'd119} : s = 161;
	{8'd18,8'd120} : s = 152;
	{8'd18,8'd121} : s = 312;
	{8'd18,8'd122} : s = 148;
	{8'd18,8'd123} : s = 308;
	{8'd18,8'd124} : s = 306;
	{8'd18,8'd125} : s = 425;
	{8'd18,8'd126} : s = 33;
	{8'd18,8'd127} : s = 146;
	{8'd18,8'd128} : s = 145;
	{8'd18,8'd129} : s = 305;
	{8'd18,8'd130} : s = 140;
	{8'd18,8'd131} : s = 300;
	{8'd18,8'd132} : s = 298;
	{8'd18,8'd133} : s = 422;
	{8'd18,8'd134} : s = 138;
	{8'd18,8'd135} : s = 297;
	{8'd18,8'd136} : s = 294;
	{8'd18,8'd137} : s = 421;
	{8'd18,8'd138} : s = 293;
	{8'd18,8'd139} : s = 419;
	{8'd18,8'd140} : s = 412;
	{8'd18,8'd141} : s = 486;
	{8'd18,8'd142} : s = 24;
	{8'd18,8'd143} : s = 137;
	{8'd18,8'd144} : s = 134;
	{8'd18,8'd145} : s = 291;
	{8'd18,8'd146} : s = 133;
	{8'd18,8'd147} : s = 284;
	{8'd18,8'd148} : s = 282;
	{8'd18,8'd149} : s = 410;
	{8'd18,8'd150} : s = 131;
	{8'd18,8'd151} : s = 281;
	{8'd18,8'd152} : s = 278;
	{8'd18,8'd153} : s = 409;
	{8'd18,8'd154} : s = 277;
	{8'd18,8'd155} : s = 406;
	{8'd18,8'd156} : s = 405;
	{8'd18,8'd157} : s = 485;
	{8'd18,8'd158} : s = 112;
	{8'd18,8'd159} : s = 275;
	{8'd18,8'd160} : s = 270;
	{8'd18,8'd161} : s = 403;
	{8'd18,8'd162} : s = 269;
	{8'd18,8'd163} : s = 398;
	{8'd18,8'd164} : s = 397;
	{8'd18,8'd165} : s = 483;
	{8'd18,8'd166} : s = 267;
	{8'd18,8'd167} : s = 395;
	{8'd18,8'd168} : s = 391;
	{8'd18,8'd169} : s = 476;
	{8'd18,8'd170} : s = 376;
	{8'd18,8'd171} : s = 474;
	{8'd18,8'd172} : s = 473;
	{8'd18,8'd173} : s = 506;
	{8'd18,8'd174} : s = 20;
	{8'd18,8'd175} : s = 104;
	{8'd18,8'd176} : s = 100;
	{8'd18,8'd177} : s = 263;
	{8'd18,8'd178} : s = 98;
	{8'd18,8'd179} : s = 240;
	{8'd18,8'd180} : s = 232;
	{8'd18,8'd181} : s = 372;
	{8'd18,8'd182} : s = 97;
	{8'd18,8'd183} : s = 228;
	{8'd18,8'd184} : s = 226;
	{8'd18,8'd185} : s = 370;
	{8'd18,8'd186} : s = 225;
	{8'd18,8'd187} : s = 369;
	{8'd18,8'd188} : s = 364;
	{8'd18,8'd189} : s = 470;
	{8'd18,8'd190} : s = 88;
	{8'd18,8'd191} : s = 216;
	{8'd18,8'd192} : s = 212;
	{8'd18,8'd193} : s = 362;
	{8'd18,8'd194} : s = 210;
	{8'd18,8'd195} : s = 361;
	{8'd18,8'd196} : s = 358;
	{8'd18,8'd197} : s = 469;
	{8'd18,8'd198} : s = 209;
	{8'd18,8'd199} : s = 357;
	{8'd18,8'd200} : s = 355;
	{8'd18,8'd201} : s = 467;
	{8'd18,8'd202} : s = 348;
	{8'd18,8'd203} : s = 462;
	{8'd18,8'd204} : s = 461;
	{8'd18,8'd205} : s = 505;
	{8'd18,8'd206} : s = 84;
	{8'd18,8'd207} : s = 204;
	{8'd18,8'd208} : s = 202;
	{8'd18,8'd209} : s = 346;
	{8'd18,8'd210} : s = 201;
	{8'd18,8'd211} : s = 345;
	{8'd18,8'd212} : s = 342;
	{8'd18,8'd213} : s = 459;
	{8'd18,8'd214} : s = 198;
	{8'd18,8'd215} : s = 341;
	{8'd18,8'd216} : s = 339;
	{8'd18,8'd217} : s = 455;
	{8'd18,8'd218} : s = 334;
	{8'd18,8'd219} : s = 444;
	{8'd18,8'd220} : s = 442;
	{8'd18,8'd221} : s = 502;
	{8'd18,8'd222} : s = 197;
	{8'd18,8'd223} : s = 333;
	{8'd18,8'd224} : s = 331;
	{8'd18,8'd225} : s = 441;
	{8'd18,8'd226} : s = 327;
	{8'd18,8'd227} : s = 438;
	{8'd18,8'd228} : s = 437;
	{8'd18,8'd229} : s = 501;
	{8'd18,8'd230} : s = 316;
	{8'd18,8'd231} : s = 435;
	{8'd18,8'd232} : s = 430;
	{8'd18,8'd233} : s = 499;
	{8'd18,8'd234} : s = 429;
	{8'd18,8'd235} : s = 494;
	{8'd18,8'd236} : s = 493;
	{8'd18,8'd237} : s = 510;
	{8'd18,8'd238} : s = 1;
	{8'd18,8'd239} : s = 18;
	{8'd18,8'd240} : s = 17;
	{8'd18,8'd241} : s = 82;
	{8'd18,8'd242} : s = 12;
	{8'd18,8'd243} : s = 81;
	{8'd18,8'd244} : s = 76;
	{8'd18,8'd245} : s = 195;
	{8'd18,8'd246} : s = 10;
	{8'd18,8'd247} : s = 74;
	{8'd18,8'd248} : s = 73;
	{8'd18,8'd249} : s = 184;
	{8'd18,8'd250} : s = 70;
	{8'd18,8'd251} : s = 180;
	{8'd18,8'd252} : s = 178;
	{8'd18,8'd253} : s = 314;
	{8'd18,8'd254} : s = 9;
	{8'd18,8'd255} : s = 69;
	{8'd19,8'd0} : s = 388;
	{8'd19,8'd1} : s = 192;
	{8'd19,8'd2} : s = 386;
	{8'd19,8'd3} : s = 385;
	{8'd19,8'd4} : s = 464;
	{8'd19,8'd5} : s = 160;
	{8'd19,8'd6} : s = 352;
	{8'd19,8'd7} : s = 336;
	{8'd19,8'd8} : s = 456;
	{8'd19,8'd9} : s = 328;
	{8'd19,8'd10} : s = 452;
	{8'd19,8'd11} : s = 450;
	{8'd19,8'd12} : s = 496;
	{8'd19,8'd13} : s = 16;
	{8'd19,8'd14} : s = 144;
	{8'd19,8'd15} : s = 136;
	{8'd19,8'd16} : s = 324;
	{8'd19,8'd17} : s = 132;
	{8'd19,8'd18} : s = 322;
	{8'd19,8'd19} : s = 321;
	{8'd19,8'd20} : s = 449;
	{8'd19,8'd21} : s = 130;
	{8'd19,8'd22} : s = 304;
	{8'd19,8'd23} : s = 296;
	{8'd19,8'd24} : s = 432;
	{8'd19,8'd25} : s = 292;
	{8'd19,8'd26} : s = 424;
	{8'd19,8'd27} : s = 420;
	{8'd19,8'd28} : s = 488;
	{8'd19,8'd29} : s = 129;
	{8'd19,8'd30} : s = 290;
	{8'd19,8'd31} : s = 289;
	{8'd19,8'd32} : s = 418;
	{8'd19,8'd33} : s = 280;
	{8'd19,8'd34} : s = 417;
	{8'd19,8'd35} : s = 408;
	{8'd19,8'd36} : s = 484;
	{8'd19,8'd37} : s = 276;
	{8'd19,8'd38} : s = 404;
	{8'd19,8'd39} : s = 402;
	{8'd19,8'd40} : s = 482;
	{8'd19,8'd41} : s = 401;
	{8'd19,8'd42} : s = 481;
	{8'd19,8'd43} : s = 472;
	{8'd19,8'd44} : s = 504;
	{8'd19,8'd45} : s = 4;
	{8'd19,8'd46} : s = 96;
	{8'd19,8'd47} : s = 80;
	{8'd19,8'd48} : s = 274;
	{8'd19,8'd49} : s = 72;
	{8'd19,8'd50} : s = 273;
	{8'd19,8'd51} : s = 268;
	{8'd19,8'd52} : s = 396;
	{8'd19,8'd53} : s = 68;
	{8'd19,8'd54} : s = 266;
	{8'd19,8'd55} : s = 265;
	{8'd19,8'd56} : s = 394;
	{8'd19,8'd57} : s = 262;
	{8'd19,8'd58} : s = 393;
	{8'd19,8'd59} : s = 390;
	{8'd19,8'd60} : s = 468;
	{8'd19,8'd61} : s = 66;
	{8'd19,8'd62} : s = 261;
	{8'd19,8'd63} : s = 259;
	{8'd19,8'd64} : s = 389;
	{8'd19,8'd65} : s = 224;
	{8'd19,8'd66} : s = 387;
	{8'd19,8'd67} : s = 368;
	{8'd19,8'd68} : s = 466;
	{8'd19,8'd69} : s = 208;
	{8'd19,8'd70} : s = 360;
	{8'd19,8'd71} : s = 356;
	{8'd19,8'd72} : s = 465;
	{8'd19,8'd73} : s = 354;
	{8'd19,8'd74} : s = 460;
	{8'd19,8'd75} : s = 458;
	{8'd19,8'd76} : s = 500;
	{8'd19,8'd77} : s = 65;
	{8'd19,8'd78} : s = 200;
	{8'd19,8'd79} : s = 196;
	{8'd19,8'd80} : s = 353;
	{8'd19,8'd81} : s = 194;
	{8'd19,8'd82} : s = 344;
	{8'd19,8'd83} : s = 340;
	{8'd19,8'd84} : s = 457;
	{8'd19,8'd85} : s = 193;
	{8'd19,8'd86} : s = 338;
	{8'd19,8'd87} : s = 337;
	{8'd19,8'd88} : s = 454;
	{8'd19,8'd89} : s = 332;
	{8'd19,8'd90} : s = 453;
	{8'd19,8'd91} : s = 451;
	{8'd19,8'd92} : s = 498;
	{8'd19,8'd93} : s = 176;
	{8'd19,8'd94} : s = 330;
	{8'd19,8'd95} : s = 329;
	{8'd19,8'd96} : s = 440;
	{8'd19,8'd97} : s = 326;
	{8'd19,8'd98} : s = 436;
	{8'd19,8'd99} : s = 434;
	{8'd19,8'd100} : s = 497;
	{8'd19,8'd101} : s = 325;
	{8'd19,8'd102} : s = 433;
	{8'd19,8'd103} : s = 428;
	{8'd19,8'd104} : s = 492;
	{8'd19,8'd105} : s = 426;
	{8'd19,8'd106} : s = 490;
	{8'd19,8'd107} : s = 489;
	{8'd19,8'd108} : s = 508;
	{8'd19,8'd109} : s = 2;
	{8'd19,8'd110} : s = 48;
	{8'd19,8'd111} : s = 40;
	{8'd19,8'd112} : s = 168;
	{8'd19,8'd113} : s = 36;
	{8'd19,8'd114} : s = 164;
	{8'd19,8'd115} : s = 162;
	{8'd19,8'd116} : s = 323;
	{8'd19,8'd117} : s = 34;
	{8'd19,8'd118} : s = 161;
	{8'd19,8'd119} : s = 152;
	{8'd19,8'd120} : s = 312;
	{8'd19,8'd121} : s = 148;
	{8'd19,8'd122} : s = 308;
	{8'd19,8'd123} : s = 306;
	{8'd19,8'd124} : s = 425;
	{8'd19,8'd125} : s = 33;
	{8'd19,8'd126} : s = 146;
	{8'd19,8'd127} : s = 145;
	{8'd19,8'd128} : s = 305;
	{8'd19,8'd129} : s = 140;
	{8'd19,8'd130} : s = 300;
	{8'd19,8'd131} : s = 298;
	{8'd19,8'd132} : s = 422;
	{8'd19,8'd133} : s = 138;
	{8'd19,8'd134} : s = 297;
	{8'd19,8'd135} : s = 294;
	{8'd19,8'd136} : s = 421;
	{8'd19,8'd137} : s = 293;
	{8'd19,8'd138} : s = 419;
	{8'd19,8'd139} : s = 412;
	{8'd19,8'd140} : s = 486;
	{8'd19,8'd141} : s = 24;
	{8'd19,8'd142} : s = 137;
	{8'd19,8'd143} : s = 134;
	{8'd19,8'd144} : s = 291;
	{8'd19,8'd145} : s = 133;
	{8'd19,8'd146} : s = 284;
	{8'd19,8'd147} : s = 282;
	{8'd19,8'd148} : s = 410;
	{8'd19,8'd149} : s = 131;
	{8'd19,8'd150} : s = 281;
	{8'd19,8'd151} : s = 278;
	{8'd19,8'd152} : s = 409;
	{8'd19,8'd153} : s = 277;
	{8'd19,8'd154} : s = 406;
	{8'd19,8'd155} : s = 405;
	{8'd19,8'd156} : s = 485;
	{8'd19,8'd157} : s = 112;
	{8'd19,8'd158} : s = 275;
	{8'd19,8'd159} : s = 270;
	{8'd19,8'd160} : s = 403;
	{8'd19,8'd161} : s = 269;
	{8'd19,8'd162} : s = 398;
	{8'd19,8'd163} : s = 397;
	{8'd19,8'd164} : s = 483;
	{8'd19,8'd165} : s = 267;
	{8'd19,8'd166} : s = 395;
	{8'd19,8'd167} : s = 391;
	{8'd19,8'd168} : s = 476;
	{8'd19,8'd169} : s = 376;
	{8'd19,8'd170} : s = 474;
	{8'd19,8'd171} : s = 473;
	{8'd19,8'd172} : s = 506;
	{8'd19,8'd173} : s = 20;
	{8'd19,8'd174} : s = 104;
	{8'd19,8'd175} : s = 100;
	{8'd19,8'd176} : s = 263;
	{8'd19,8'd177} : s = 98;
	{8'd19,8'd178} : s = 240;
	{8'd19,8'd179} : s = 232;
	{8'd19,8'd180} : s = 372;
	{8'd19,8'd181} : s = 97;
	{8'd19,8'd182} : s = 228;
	{8'd19,8'd183} : s = 226;
	{8'd19,8'd184} : s = 370;
	{8'd19,8'd185} : s = 225;
	{8'd19,8'd186} : s = 369;
	{8'd19,8'd187} : s = 364;
	{8'd19,8'd188} : s = 470;
	{8'd19,8'd189} : s = 88;
	{8'd19,8'd190} : s = 216;
	{8'd19,8'd191} : s = 212;
	{8'd19,8'd192} : s = 362;
	{8'd19,8'd193} : s = 210;
	{8'd19,8'd194} : s = 361;
	{8'd19,8'd195} : s = 358;
	{8'd19,8'd196} : s = 469;
	{8'd19,8'd197} : s = 209;
	{8'd19,8'd198} : s = 357;
	{8'd19,8'd199} : s = 355;
	{8'd19,8'd200} : s = 467;
	{8'd19,8'd201} : s = 348;
	{8'd19,8'd202} : s = 462;
	{8'd19,8'd203} : s = 461;
	{8'd19,8'd204} : s = 505;
	{8'd19,8'd205} : s = 84;
	{8'd19,8'd206} : s = 204;
	{8'd19,8'd207} : s = 202;
	{8'd19,8'd208} : s = 346;
	{8'd19,8'd209} : s = 201;
	{8'd19,8'd210} : s = 345;
	{8'd19,8'd211} : s = 342;
	{8'd19,8'd212} : s = 459;
	{8'd19,8'd213} : s = 198;
	{8'd19,8'd214} : s = 341;
	{8'd19,8'd215} : s = 339;
	{8'd19,8'd216} : s = 455;
	{8'd19,8'd217} : s = 334;
	{8'd19,8'd218} : s = 444;
	{8'd19,8'd219} : s = 442;
	{8'd19,8'd220} : s = 502;
	{8'd19,8'd221} : s = 197;
	{8'd19,8'd222} : s = 333;
	{8'd19,8'd223} : s = 331;
	{8'd19,8'd224} : s = 441;
	{8'd19,8'd225} : s = 327;
	{8'd19,8'd226} : s = 438;
	{8'd19,8'd227} : s = 437;
	{8'd19,8'd228} : s = 501;
	{8'd19,8'd229} : s = 316;
	{8'd19,8'd230} : s = 435;
	{8'd19,8'd231} : s = 430;
	{8'd19,8'd232} : s = 499;
	{8'd19,8'd233} : s = 429;
	{8'd19,8'd234} : s = 494;
	{8'd19,8'd235} : s = 493;
	{8'd19,8'd236} : s = 510;
	{8'd19,8'd237} : s = 1;
	{8'd19,8'd238} : s = 18;
	{8'd19,8'd239} : s = 17;
	{8'd19,8'd240} : s = 82;
	{8'd19,8'd241} : s = 12;
	{8'd19,8'd242} : s = 81;
	{8'd19,8'd243} : s = 76;
	{8'd19,8'd244} : s = 195;
	{8'd19,8'd245} : s = 10;
	{8'd19,8'd246} : s = 74;
	{8'd19,8'd247} : s = 73;
	{8'd19,8'd248} : s = 184;
	{8'd19,8'd249} : s = 70;
	{8'd19,8'd250} : s = 180;
	{8'd19,8'd251} : s = 178;
	{8'd19,8'd252} : s = 314;
	{8'd19,8'd253} : s = 9;
	{8'd19,8'd254} : s = 69;
	{8'd19,8'd255} : s = 67;
	{8'd20,8'd0} : s = 192;
	{8'd20,8'd1} : s = 386;
	{8'd20,8'd2} : s = 385;
	{8'd20,8'd3} : s = 464;
	{8'd20,8'd4} : s = 160;
	{8'd20,8'd5} : s = 352;
	{8'd20,8'd6} : s = 336;
	{8'd20,8'd7} : s = 456;
	{8'd20,8'd8} : s = 328;
	{8'd20,8'd9} : s = 452;
	{8'd20,8'd10} : s = 450;
	{8'd20,8'd11} : s = 496;
	{8'd20,8'd12} : s = 16;
	{8'd20,8'd13} : s = 144;
	{8'd20,8'd14} : s = 136;
	{8'd20,8'd15} : s = 324;
	{8'd20,8'd16} : s = 132;
	{8'd20,8'd17} : s = 322;
	{8'd20,8'd18} : s = 321;
	{8'd20,8'd19} : s = 449;
	{8'd20,8'd20} : s = 130;
	{8'd20,8'd21} : s = 304;
	{8'd20,8'd22} : s = 296;
	{8'd20,8'd23} : s = 432;
	{8'd20,8'd24} : s = 292;
	{8'd20,8'd25} : s = 424;
	{8'd20,8'd26} : s = 420;
	{8'd20,8'd27} : s = 488;
	{8'd20,8'd28} : s = 129;
	{8'd20,8'd29} : s = 290;
	{8'd20,8'd30} : s = 289;
	{8'd20,8'd31} : s = 418;
	{8'd20,8'd32} : s = 280;
	{8'd20,8'd33} : s = 417;
	{8'd20,8'd34} : s = 408;
	{8'd20,8'd35} : s = 484;
	{8'd20,8'd36} : s = 276;
	{8'd20,8'd37} : s = 404;
	{8'd20,8'd38} : s = 402;
	{8'd20,8'd39} : s = 482;
	{8'd20,8'd40} : s = 401;
	{8'd20,8'd41} : s = 481;
	{8'd20,8'd42} : s = 472;
	{8'd20,8'd43} : s = 504;
	{8'd20,8'd44} : s = 4;
	{8'd20,8'd45} : s = 96;
	{8'd20,8'd46} : s = 80;
	{8'd20,8'd47} : s = 274;
	{8'd20,8'd48} : s = 72;
	{8'd20,8'd49} : s = 273;
	{8'd20,8'd50} : s = 268;
	{8'd20,8'd51} : s = 396;
	{8'd20,8'd52} : s = 68;
	{8'd20,8'd53} : s = 266;
	{8'd20,8'd54} : s = 265;
	{8'd20,8'd55} : s = 394;
	{8'd20,8'd56} : s = 262;
	{8'd20,8'd57} : s = 393;
	{8'd20,8'd58} : s = 390;
	{8'd20,8'd59} : s = 468;
	{8'd20,8'd60} : s = 66;
	{8'd20,8'd61} : s = 261;
	{8'd20,8'd62} : s = 259;
	{8'd20,8'd63} : s = 389;
	{8'd20,8'd64} : s = 224;
	{8'd20,8'd65} : s = 387;
	{8'd20,8'd66} : s = 368;
	{8'd20,8'd67} : s = 466;
	{8'd20,8'd68} : s = 208;
	{8'd20,8'd69} : s = 360;
	{8'd20,8'd70} : s = 356;
	{8'd20,8'd71} : s = 465;
	{8'd20,8'd72} : s = 354;
	{8'd20,8'd73} : s = 460;
	{8'd20,8'd74} : s = 458;
	{8'd20,8'd75} : s = 500;
	{8'd20,8'd76} : s = 65;
	{8'd20,8'd77} : s = 200;
	{8'd20,8'd78} : s = 196;
	{8'd20,8'd79} : s = 353;
	{8'd20,8'd80} : s = 194;
	{8'd20,8'd81} : s = 344;
	{8'd20,8'd82} : s = 340;
	{8'd20,8'd83} : s = 457;
	{8'd20,8'd84} : s = 193;
	{8'd20,8'd85} : s = 338;
	{8'd20,8'd86} : s = 337;
	{8'd20,8'd87} : s = 454;
	{8'd20,8'd88} : s = 332;
	{8'd20,8'd89} : s = 453;
	{8'd20,8'd90} : s = 451;
	{8'd20,8'd91} : s = 498;
	{8'd20,8'd92} : s = 176;
	{8'd20,8'd93} : s = 330;
	{8'd20,8'd94} : s = 329;
	{8'd20,8'd95} : s = 440;
	{8'd20,8'd96} : s = 326;
	{8'd20,8'd97} : s = 436;
	{8'd20,8'd98} : s = 434;
	{8'd20,8'd99} : s = 497;
	{8'd20,8'd100} : s = 325;
	{8'd20,8'd101} : s = 433;
	{8'd20,8'd102} : s = 428;
	{8'd20,8'd103} : s = 492;
	{8'd20,8'd104} : s = 426;
	{8'd20,8'd105} : s = 490;
	{8'd20,8'd106} : s = 489;
	{8'd20,8'd107} : s = 508;
	{8'd20,8'd108} : s = 2;
	{8'd20,8'd109} : s = 48;
	{8'd20,8'd110} : s = 40;
	{8'd20,8'd111} : s = 168;
	{8'd20,8'd112} : s = 36;
	{8'd20,8'd113} : s = 164;
	{8'd20,8'd114} : s = 162;
	{8'd20,8'd115} : s = 323;
	{8'd20,8'd116} : s = 34;
	{8'd20,8'd117} : s = 161;
	{8'd20,8'd118} : s = 152;
	{8'd20,8'd119} : s = 312;
	{8'd20,8'd120} : s = 148;
	{8'd20,8'd121} : s = 308;
	{8'd20,8'd122} : s = 306;
	{8'd20,8'd123} : s = 425;
	{8'd20,8'd124} : s = 33;
	{8'd20,8'd125} : s = 146;
	{8'd20,8'd126} : s = 145;
	{8'd20,8'd127} : s = 305;
	{8'd20,8'd128} : s = 140;
	{8'd20,8'd129} : s = 300;
	{8'd20,8'd130} : s = 298;
	{8'd20,8'd131} : s = 422;
	{8'd20,8'd132} : s = 138;
	{8'd20,8'd133} : s = 297;
	{8'd20,8'd134} : s = 294;
	{8'd20,8'd135} : s = 421;
	{8'd20,8'd136} : s = 293;
	{8'd20,8'd137} : s = 419;
	{8'd20,8'd138} : s = 412;
	{8'd20,8'd139} : s = 486;
	{8'd20,8'd140} : s = 24;
	{8'd20,8'd141} : s = 137;
	{8'd20,8'd142} : s = 134;
	{8'd20,8'd143} : s = 291;
	{8'd20,8'd144} : s = 133;
	{8'd20,8'd145} : s = 284;
	{8'd20,8'd146} : s = 282;
	{8'd20,8'd147} : s = 410;
	{8'd20,8'd148} : s = 131;
	{8'd20,8'd149} : s = 281;
	{8'd20,8'd150} : s = 278;
	{8'd20,8'd151} : s = 409;
	{8'd20,8'd152} : s = 277;
	{8'd20,8'd153} : s = 406;
	{8'd20,8'd154} : s = 405;
	{8'd20,8'd155} : s = 485;
	{8'd20,8'd156} : s = 112;
	{8'd20,8'd157} : s = 275;
	{8'd20,8'd158} : s = 270;
	{8'd20,8'd159} : s = 403;
	{8'd20,8'd160} : s = 269;
	{8'd20,8'd161} : s = 398;
	{8'd20,8'd162} : s = 397;
	{8'd20,8'd163} : s = 483;
	{8'd20,8'd164} : s = 267;
	{8'd20,8'd165} : s = 395;
	{8'd20,8'd166} : s = 391;
	{8'd20,8'd167} : s = 476;
	{8'd20,8'd168} : s = 376;
	{8'd20,8'd169} : s = 474;
	{8'd20,8'd170} : s = 473;
	{8'd20,8'd171} : s = 506;
	{8'd20,8'd172} : s = 20;
	{8'd20,8'd173} : s = 104;
	{8'd20,8'd174} : s = 100;
	{8'd20,8'd175} : s = 263;
	{8'd20,8'd176} : s = 98;
	{8'd20,8'd177} : s = 240;
	{8'd20,8'd178} : s = 232;
	{8'd20,8'd179} : s = 372;
	{8'd20,8'd180} : s = 97;
	{8'd20,8'd181} : s = 228;
	{8'd20,8'd182} : s = 226;
	{8'd20,8'd183} : s = 370;
	{8'd20,8'd184} : s = 225;
	{8'd20,8'd185} : s = 369;
	{8'd20,8'd186} : s = 364;
	{8'd20,8'd187} : s = 470;
	{8'd20,8'd188} : s = 88;
	{8'd20,8'd189} : s = 216;
	{8'd20,8'd190} : s = 212;
	{8'd20,8'd191} : s = 362;
	{8'd20,8'd192} : s = 210;
	{8'd20,8'd193} : s = 361;
	{8'd20,8'd194} : s = 358;
	{8'd20,8'd195} : s = 469;
	{8'd20,8'd196} : s = 209;
	{8'd20,8'd197} : s = 357;
	{8'd20,8'd198} : s = 355;
	{8'd20,8'd199} : s = 467;
	{8'd20,8'd200} : s = 348;
	{8'd20,8'd201} : s = 462;
	{8'd20,8'd202} : s = 461;
	{8'd20,8'd203} : s = 505;
	{8'd20,8'd204} : s = 84;
	{8'd20,8'd205} : s = 204;
	{8'd20,8'd206} : s = 202;
	{8'd20,8'd207} : s = 346;
	{8'd20,8'd208} : s = 201;
	{8'd20,8'd209} : s = 345;
	{8'd20,8'd210} : s = 342;
	{8'd20,8'd211} : s = 459;
	{8'd20,8'd212} : s = 198;
	{8'd20,8'd213} : s = 341;
	{8'd20,8'd214} : s = 339;
	{8'd20,8'd215} : s = 455;
	{8'd20,8'd216} : s = 334;
	{8'd20,8'd217} : s = 444;
	{8'd20,8'd218} : s = 442;
	{8'd20,8'd219} : s = 502;
	{8'd20,8'd220} : s = 197;
	{8'd20,8'd221} : s = 333;
	{8'd20,8'd222} : s = 331;
	{8'd20,8'd223} : s = 441;
	{8'd20,8'd224} : s = 327;
	{8'd20,8'd225} : s = 438;
	{8'd20,8'd226} : s = 437;
	{8'd20,8'd227} : s = 501;
	{8'd20,8'd228} : s = 316;
	{8'd20,8'd229} : s = 435;
	{8'd20,8'd230} : s = 430;
	{8'd20,8'd231} : s = 499;
	{8'd20,8'd232} : s = 429;
	{8'd20,8'd233} : s = 494;
	{8'd20,8'd234} : s = 493;
	{8'd20,8'd235} : s = 510;
	{8'd20,8'd236} : s = 1;
	{8'd20,8'd237} : s = 18;
	{8'd20,8'd238} : s = 17;
	{8'd20,8'd239} : s = 82;
	{8'd20,8'd240} : s = 12;
	{8'd20,8'd241} : s = 81;
	{8'd20,8'd242} : s = 76;
	{8'd20,8'd243} : s = 195;
	{8'd20,8'd244} : s = 10;
	{8'd20,8'd245} : s = 74;
	{8'd20,8'd246} : s = 73;
	{8'd20,8'd247} : s = 184;
	{8'd20,8'd248} : s = 70;
	{8'd20,8'd249} : s = 180;
	{8'd20,8'd250} : s = 178;
	{8'd20,8'd251} : s = 314;
	{8'd20,8'd252} : s = 9;
	{8'd20,8'd253} : s = 69;
	{8'd20,8'd254} : s = 67;
	{8'd20,8'd255} : s = 177;
	{8'd21,8'd0} : s = 386;
	{8'd21,8'd1} : s = 385;
	{8'd21,8'd2} : s = 464;
	{8'd21,8'd3} : s = 160;
	{8'd21,8'd4} : s = 352;
	{8'd21,8'd5} : s = 336;
	{8'd21,8'd6} : s = 456;
	{8'd21,8'd7} : s = 328;
	{8'd21,8'd8} : s = 452;
	{8'd21,8'd9} : s = 450;
	{8'd21,8'd10} : s = 496;
	{8'd21,8'd11} : s = 16;
	{8'd21,8'd12} : s = 144;
	{8'd21,8'd13} : s = 136;
	{8'd21,8'd14} : s = 324;
	{8'd21,8'd15} : s = 132;
	{8'd21,8'd16} : s = 322;
	{8'd21,8'd17} : s = 321;
	{8'd21,8'd18} : s = 449;
	{8'd21,8'd19} : s = 130;
	{8'd21,8'd20} : s = 304;
	{8'd21,8'd21} : s = 296;
	{8'd21,8'd22} : s = 432;
	{8'd21,8'd23} : s = 292;
	{8'd21,8'd24} : s = 424;
	{8'd21,8'd25} : s = 420;
	{8'd21,8'd26} : s = 488;
	{8'd21,8'd27} : s = 129;
	{8'd21,8'd28} : s = 290;
	{8'd21,8'd29} : s = 289;
	{8'd21,8'd30} : s = 418;
	{8'd21,8'd31} : s = 280;
	{8'd21,8'd32} : s = 417;
	{8'd21,8'd33} : s = 408;
	{8'd21,8'd34} : s = 484;
	{8'd21,8'd35} : s = 276;
	{8'd21,8'd36} : s = 404;
	{8'd21,8'd37} : s = 402;
	{8'd21,8'd38} : s = 482;
	{8'd21,8'd39} : s = 401;
	{8'd21,8'd40} : s = 481;
	{8'd21,8'd41} : s = 472;
	{8'd21,8'd42} : s = 504;
	{8'd21,8'd43} : s = 4;
	{8'd21,8'd44} : s = 96;
	{8'd21,8'd45} : s = 80;
	{8'd21,8'd46} : s = 274;
	{8'd21,8'd47} : s = 72;
	{8'd21,8'd48} : s = 273;
	{8'd21,8'd49} : s = 268;
	{8'd21,8'd50} : s = 396;
	{8'd21,8'd51} : s = 68;
	{8'd21,8'd52} : s = 266;
	{8'd21,8'd53} : s = 265;
	{8'd21,8'd54} : s = 394;
	{8'd21,8'd55} : s = 262;
	{8'd21,8'd56} : s = 393;
	{8'd21,8'd57} : s = 390;
	{8'd21,8'd58} : s = 468;
	{8'd21,8'd59} : s = 66;
	{8'd21,8'd60} : s = 261;
	{8'd21,8'd61} : s = 259;
	{8'd21,8'd62} : s = 389;
	{8'd21,8'd63} : s = 224;
	{8'd21,8'd64} : s = 387;
	{8'd21,8'd65} : s = 368;
	{8'd21,8'd66} : s = 466;
	{8'd21,8'd67} : s = 208;
	{8'd21,8'd68} : s = 360;
	{8'd21,8'd69} : s = 356;
	{8'd21,8'd70} : s = 465;
	{8'd21,8'd71} : s = 354;
	{8'd21,8'd72} : s = 460;
	{8'd21,8'd73} : s = 458;
	{8'd21,8'd74} : s = 500;
	{8'd21,8'd75} : s = 65;
	{8'd21,8'd76} : s = 200;
	{8'd21,8'd77} : s = 196;
	{8'd21,8'd78} : s = 353;
	{8'd21,8'd79} : s = 194;
	{8'd21,8'd80} : s = 344;
	{8'd21,8'd81} : s = 340;
	{8'd21,8'd82} : s = 457;
	{8'd21,8'd83} : s = 193;
	{8'd21,8'd84} : s = 338;
	{8'd21,8'd85} : s = 337;
	{8'd21,8'd86} : s = 454;
	{8'd21,8'd87} : s = 332;
	{8'd21,8'd88} : s = 453;
	{8'd21,8'd89} : s = 451;
	{8'd21,8'd90} : s = 498;
	{8'd21,8'd91} : s = 176;
	{8'd21,8'd92} : s = 330;
	{8'd21,8'd93} : s = 329;
	{8'd21,8'd94} : s = 440;
	{8'd21,8'd95} : s = 326;
	{8'd21,8'd96} : s = 436;
	{8'd21,8'd97} : s = 434;
	{8'd21,8'd98} : s = 497;
	{8'd21,8'd99} : s = 325;
	{8'd21,8'd100} : s = 433;
	{8'd21,8'd101} : s = 428;
	{8'd21,8'd102} : s = 492;
	{8'd21,8'd103} : s = 426;
	{8'd21,8'd104} : s = 490;
	{8'd21,8'd105} : s = 489;
	{8'd21,8'd106} : s = 508;
	{8'd21,8'd107} : s = 2;
	{8'd21,8'd108} : s = 48;
	{8'd21,8'd109} : s = 40;
	{8'd21,8'd110} : s = 168;
	{8'd21,8'd111} : s = 36;
	{8'd21,8'd112} : s = 164;
	{8'd21,8'd113} : s = 162;
	{8'd21,8'd114} : s = 323;
	{8'd21,8'd115} : s = 34;
	{8'd21,8'd116} : s = 161;
	{8'd21,8'd117} : s = 152;
	{8'd21,8'd118} : s = 312;
	{8'd21,8'd119} : s = 148;
	{8'd21,8'd120} : s = 308;
	{8'd21,8'd121} : s = 306;
	{8'd21,8'd122} : s = 425;
	{8'd21,8'd123} : s = 33;
	{8'd21,8'd124} : s = 146;
	{8'd21,8'd125} : s = 145;
	{8'd21,8'd126} : s = 305;
	{8'd21,8'd127} : s = 140;
	{8'd21,8'd128} : s = 300;
	{8'd21,8'd129} : s = 298;
	{8'd21,8'd130} : s = 422;
	{8'd21,8'd131} : s = 138;
	{8'd21,8'd132} : s = 297;
	{8'd21,8'd133} : s = 294;
	{8'd21,8'd134} : s = 421;
	{8'd21,8'd135} : s = 293;
	{8'd21,8'd136} : s = 419;
	{8'd21,8'd137} : s = 412;
	{8'd21,8'd138} : s = 486;
	{8'd21,8'd139} : s = 24;
	{8'd21,8'd140} : s = 137;
	{8'd21,8'd141} : s = 134;
	{8'd21,8'd142} : s = 291;
	{8'd21,8'd143} : s = 133;
	{8'd21,8'd144} : s = 284;
	{8'd21,8'd145} : s = 282;
	{8'd21,8'd146} : s = 410;
	{8'd21,8'd147} : s = 131;
	{8'd21,8'd148} : s = 281;
	{8'd21,8'd149} : s = 278;
	{8'd21,8'd150} : s = 409;
	{8'd21,8'd151} : s = 277;
	{8'd21,8'd152} : s = 406;
	{8'd21,8'd153} : s = 405;
	{8'd21,8'd154} : s = 485;
	{8'd21,8'd155} : s = 112;
	{8'd21,8'd156} : s = 275;
	{8'd21,8'd157} : s = 270;
	{8'd21,8'd158} : s = 403;
	{8'd21,8'd159} : s = 269;
	{8'd21,8'd160} : s = 398;
	{8'd21,8'd161} : s = 397;
	{8'd21,8'd162} : s = 483;
	{8'd21,8'd163} : s = 267;
	{8'd21,8'd164} : s = 395;
	{8'd21,8'd165} : s = 391;
	{8'd21,8'd166} : s = 476;
	{8'd21,8'd167} : s = 376;
	{8'd21,8'd168} : s = 474;
	{8'd21,8'd169} : s = 473;
	{8'd21,8'd170} : s = 506;
	{8'd21,8'd171} : s = 20;
	{8'd21,8'd172} : s = 104;
	{8'd21,8'd173} : s = 100;
	{8'd21,8'd174} : s = 263;
	{8'd21,8'd175} : s = 98;
	{8'd21,8'd176} : s = 240;
	{8'd21,8'd177} : s = 232;
	{8'd21,8'd178} : s = 372;
	{8'd21,8'd179} : s = 97;
	{8'd21,8'd180} : s = 228;
	{8'd21,8'd181} : s = 226;
	{8'd21,8'd182} : s = 370;
	{8'd21,8'd183} : s = 225;
	{8'd21,8'd184} : s = 369;
	{8'd21,8'd185} : s = 364;
	{8'd21,8'd186} : s = 470;
	{8'd21,8'd187} : s = 88;
	{8'd21,8'd188} : s = 216;
	{8'd21,8'd189} : s = 212;
	{8'd21,8'd190} : s = 362;
	{8'd21,8'd191} : s = 210;
	{8'd21,8'd192} : s = 361;
	{8'd21,8'd193} : s = 358;
	{8'd21,8'd194} : s = 469;
	{8'd21,8'd195} : s = 209;
	{8'd21,8'd196} : s = 357;
	{8'd21,8'd197} : s = 355;
	{8'd21,8'd198} : s = 467;
	{8'd21,8'd199} : s = 348;
	{8'd21,8'd200} : s = 462;
	{8'd21,8'd201} : s = 461;
	{8'd21,8'd202} : s = 505;
	{8'd21,8'd203} : s = 84;
	{8'd21,8'd204} : s = 204;
	{8'd21,8'd205} : s = 202;
	{8'd21,8'd206} : s = 346;
	{8'd21,8'd207} : s = 201;
	{8'd21,8'd208} : s = 345;
	{8'd21,8'd209} : s = 342;
	{8'd21,8'd210} : s = 459;
	{8'd21,8'd211} : s = 198;
	{8'd21,8'd212} : s = 341;
	{8'd21,8'd213} : s = 339;
	{8'd21,8'd214} : s = 455;
	{8'd21,8'd215} : s = 334;
	{8'd21,8'd216} : s = 444;
	{8'd21,8'd217} : s = 442;
	{8'd21,8'd218} : s = 502;
	{8'd21,8'd219} : s = 197;
	{8'd21,8'd220} : s = 333;
	{8'd21,8'd221} : s = 331;
	{8'd21,8'd222} : s = 441;
	{8'd21,8'd223} : s = 327;
	{8'd21,8'd224} : s = 438;
	{8'd21,8'd225} : s = 437;
	{8'd21,8'd226} : s = 501;
	{8'd21,8'd227} : s = 316;
	{8'd21,8'd228} : s = 435;
	{8'd21,8'd229} : s = 430;
	{8'd21,8'd230} : s = 499;
	{8'd21,8'd231} : s = 429;
	{8'd21,8'd232} : s = 494;
	{8'd21,8'd233} : s = 493;
	{8'd21,8'd234} : s = 510;
	{8'd21,8'd235} : s = 1;
	{8'd21,8'd236} : s = 18;
	{8'd21,8'd237} : s = 17;
	{8'd21,8'd238} : s = 82;
	{8'd21,8'd239} : s = 12;
	{8'd21,8'd240} : s = 81;
	{8'd21,8'd241} : s = 76;
	{8'd21,8'd242} : s = 195;
	{8'd21,8'd243} : s = 10;
	{8'd21,8'd244} : s = 74;
	{8'd21,8'd245} : s = 73;
	{8'd21,8'd246} : s = 184;
	{8'd21,8'd247} : s = 70;
	{8'd21,8'd248} : s = 180;
	{8'd21,8'd249} : s = 178;
	{8'd21,8'd250} : s = 314;
	{8'd21,8'd251} : s = 9;
	{8'd21,8'd252} : s = 69;
	{8'd21,8'd253} : s = 67;
	{8'd21,8'd254} : s = 177;
	{8'd21,8'd255} : s = 56;
	{8'd22,8'd0} : s = 385;
	{8'd22,8'd1} : s = 464;
	{8'd22,8'd2} : s = 160;
	{8'd22,8'd3} : s = 352;
	{8'd22,8'd4} : s = 336;
	{8'd22,8'd5} : s = 456;
	{8'd22,8'd6} : s = 328;
	{8'd22,8'd7} : s = 452;
	{8'd22,8'd8} : s = 450;
	{8'd22,8'd9} : s = 496;
	{8'd22,8'd10} : s = 16;
	{8'd22,8'd11} : s = 144;
	{8'd22,8'd12} : s = 136;
	{8'd22,8'd13} : s = 324;
	{8'd22,8'd14} : s = 132;
	{8'd22,8'd15} : s = 322;
	{8'd22,8'd16} : s = 321;
	{8'd22,8'd17} : s = 449;
	{8'd22,8'd18} : s = 130;
	{8'd22,8'd19} : s = 304;
	{8'd22,8'd20} : s = 296;
	{8'd22,8'd21} : s = 432;
	{8'd22,8'd22} : s = 292;
	{8'd22,8'd23} : s = 424;
	{8'd22,8'd24} : s = 420;
	{8'd22,8'd25} : s = 488;
	{8'd22,8'd26} : s = 129;
	{8'd22,8'd27} : s = 290;
	{8'd22,8'd28} : s = 289;
	{8'd22,8'd29} : s = 418;
	{8'd22,8'd30} : s = 280;
	{8'd22,8'd31} : s = 417;
	{8'd22,8'd32} : s = 408;
	{8'd22,8'd33} : s = 484;
	{8'd22,8'd34} : s = 276;
	{8'd22,8'd35} : s = 404;
	{8'd22,8'd36} : s = 402;
	{8'd22,8'd37} : s = 482;
	{8'd22,8'd38} : s = 401;
	{8'd22,8'd39} : s = 481;
	{8'd22,8'd40} : s = 472;
	{8'd22,8'd41} : s = 504;
	{8'd22,8'd42} : s = 4;
	{8'd22,8'd43} : s = 96;
	{8'd22,8'd44} : s = 80;
	{8'd22,8'd45} : s = 274;
	{8'd22,8'd46} : s = 72;
	{8'd22,8'd47} : s = 273;
	{8'd22,8'd48} : s = 268;
	{8'd22,8'd49} : s = 396;
	{8'd22,8'd50} : s = 68;
	{8'd22,8'd51} : s = 266;
	{8'd22,8'd52} : s = 265;
	{8'd22,8'd53} : s = 394;
	{8'd22,8'd54} : s = 262;
	{8'd22,8'd55} : s = 393;
	{8'd22,8'd56} : s = 390;
	{8'd22,8'd57} : s = 468;
	{8'd22,8'd58} : s = 66;
	{8'd22,8'd59} : s = 261;
	{8'd22,8'd60} : s = 259;
	{8'd22,8'd61} : s = 389;
	{8'd22,8'd62} : s = 224;
	{8'd22,8'd63} : s = 387;
	{8'd22,8'd64} : s = 368;
	{8'd22,8'd65} : s = 466;
	{8'd22,8'd66} : s = 208;
	{8'd22,8'd67} : s = 360;
	{8'd22,8'd68} : s = 356;
	{8'd22,8'd69} : s = 465;
	{8'd22,8'd70} : s = 354;
	{8'd22,8'd71} : s = 460;
	{8'd22,8'd72} : s = 458;
	{8'd22,8'd73} : s = 500;
	{8'd22,8'd74} : s = 65;
	{8'd22,8'd75} : s = 200;
	{8'd22,8'd76} : s = 196;
	{8'd22,8'd77} : s = 353;
	{8'd22,8'd78} : s = 194;
	{8'd22,8'd79} : s = 344;
	{8'd22,8'd80} : s = 340;
	{8'd22,8'd81} : s = 457;
	{8'd22,8'd82} : s = 193;
	{8'd22,8'd83} : s = 338;
	{8'd22,8'd84} : s = 337;
	{8'd22,8'd85} : s = 454;
	{8'd22,8'd86} : s = 332;
	{8'd22,8'd87} : s = 453;
	{8'd22,8'd88} : s = 451;
	{8'd22,8'd89} : s = 498;
	{8'd22,8'd90} : s = 176;
	{8'd22,8'd91} : s = 330;
	{8'd22,8'd92} : s = 329;
	{8'd22,8'd93} : s = 440;
	{8'd22,8'd94} : s = 326;
	{8'd22,8'd95} : s = 436;
	{8'd22,8'd96} : s = 434;
	{8'd22,8'd97} : s = 497;
	{8'd22,8'd98} : s = 325;
	{8'd22,8'd99} : s = 433;
	{8'd22,8'd100} : s = 428;
	{8'd22,8'd101} : s = 492;
	{8'd22,8'd102} : s = 426;
	{8'd22,8'd103} : s = 490;
	{8'd22,8'd104} : s = 489;
	{8'd22,8'd105} : s = 508;
	{8'd22,8'd106} : s = 2;
	{8'd22,8'd107} : s = 48;
	{8'd22,8'd108} : s = 40;
	{8'd22,8'd109} : s = 168;
	{8'd22,8'd110} : s = 36;
	{8'd22,8'd111} : s = 164;
	{8'd22,8'd112} : s = 162;
	{8'd22,8'd113} : s = 323;
	{8'd22,8'd114} : s = 34;
	{8'd22,8'd115} : s = 161;
	{8'd22,8'd116} : s = 152;
	{8'd22,8'd117} : s = 312;
	{8'd22,8'd118} : s = 148;
	{8'd22,8'd119} : s = 308;
	{8'd22,8'd120} : s = 306;
	{8'd22,8'd121} : s = 425;
	{8'd22,8'd122} : s = 33;
	{8'd22,8'd123} : s = 146;
	{8'd22,8'd124} : s = 145;
	{8'd22,8'd125} : s = 305;
	{8'd22,8'd126} : s = 140;
	{8'd22,8'd127} : s = 300;
	{8'd22,8'd128} : s = 298;
	{8'd22,8'd129} : s = 422;
	{8'd22,8'd130} : s = 138;
	{8'd22,8'd131} : s = 297;
	{8'd22,8'd132} : s = 294;
	{8'd22,8'd133} : s = 421;
	{8'd22,8'd134} : s = 293;
	{8'd22,8'd135} : s = 419;
	{8'd22,8'd136} : s = 412;
	{8'd22,8'd137} : s = 486;
	{8'd22,8'd138} : s = 24;
	{8'd22,8'd139} : s = 137;
	{8'd22,8'd140} : s = 134;
	{8'd22,8'd141} : s = 291;
	{8'd22,8'd142} : s = 133;
	{8'd22,8'd143} : s = 284;
	{8'd22,8'd144} : s = 282;
	{8'd22,8'd145} : s = 410;
	{8'd22,8'd146} : s = 131;
	{8'd22,8'd147} : s = 281;
	{8'd22,8'd148} : s = 278;
	{8'd22,8'd149} : s = 409;
	{8'd22,8'd150} : s = 277;
	{8'd22,8'd151} : s = 406;
	{8'd22,8'd152} : s = 405;
	{8'd22,8'd153} : s = 485;
	{8'd22,8'd154} : s = 112;
	{8'd22,8'd155} : s = 275;
	{8'd22,8'd156} : s = 270;
	{8'd22,8'd157} : s = 403;
	{8'd22,8'd158} : s = 269;
	{8'd22,8'd159} : s = 398;
	{8'd22,8'd160} : s = 397;
	{8'd22,8'd161} : s = 483;
	{8'd22,8'd162} : s = 267;
	{8'd22,8'd163} : s = 395;
	{8'd22,8'd164} : s = 391;
	{8'd22,8'd165} : s = 476;
	{8'd22,8'd166} : s = 376;
	{8'd22,8'd167} : s = 474;
	{8'd22,8'd168} : s = 473;
	{8'd22,8'd169} : s = 506;
	{8'd22,8'd170} : s = 20;
	{8'd22,8'd171} : s = 104;
	{8'd22,8'd172} : s = 100;
	{8'd22,8'd173} : s = 263;
	{8'd22,8'd174} : s = 98;
	{8'd22,8'd175} : s = 240;
	{8'd22,8'd176} : s = 232;
	{8'd22,8'd177} : s = 372;
	{8'd22,8'd178} : s = 97;
	{8'd22,8'd179} : s = 228;
	{8'd22,8'd180} : s = 226;
	{8'd22,8'd181} : s = 370;
	{8'd22,8'd182} : s = 225;
	{8'd22,8'd183} : s = 369;
	{8'd22,8'd184} : s = 364;
	{8'd22,8'd185} : s = 470;
	{8'd22,8'd186} : s = 88;
	{8'd22,8'd187} : s = 216;
	{8'd22,8'd188} : s = 212;
	{8'd22,8'd189} : s = 362;
	{8'd22,8'd190} : s = 210;
	{8'd22,8'd191} : s = 361;
	{8'd22,8'd192} : s = 358;
	{8'd22,8'd193} : s = 469;
	{8'd22,8'd194} : s = 209;
	{8'd22,8'd195} : s = 357;
	{8'd22,8'd196} : s = 355;
	{8'd22,8'd197} : s = 467;
	{8'd22,8'd198} : s = 348;
	{8'd22,8'd199} : s = 462;
	{8'd22,8'd200} : s = 461;
	{8'd22,8'd201} : s = 505;
	{8'd22,8'd202} : s = 84;
	{8'd22,8'd203} : s = 204;
	{8'd22,8'd204} : s = 202;
	{8'd22,8'd205} : s = 346;
	{8'd22,8'd206} : s = 201;
	{8'd22,8'd207} : s = 345;
	{8'd22,8'd208} : s = 342;
	{8'd22,8'd209} : s = 459;
	{8'd22,8'd210} : s = 198;
	{8'd22,8'd211} : s = 341;
	{8'd22,8'd212} : s = 339;
	{8'd22,8'd213} : s = 455;
	{8'd22,8'd214} : s = 334;
	{8'd22,8'd215} : s = 444;
	{8'd22,8'd216} : s = 442;
	{8'd22,8'd217} : s = 502;
	{8'd22,8'd218} : s = 197;
	{8'd22,8'd219} : s = 333;
	{8'd22,8'd220} : s = 331;
	{8'd22,8'd221} : s = 441;
	{8'd22,8'd222} : s = 327;
	{8'd22,8'd223} : s = 438;
	{8'd22,8'd224} : s = 437;
	{8'd22,8'd225} : s = 501;
	{8'd22,8'd226} : s = 316;
	{8'd22,8'd227} : s = 435;
	{8'd22,8'd228} : s = 430;
	{8'd22,8'd229} : s = 499;
	{8'd22,8'd230} : s = 429;
	{8'd22,8'd231} : s = 494;
	{8'd22,8'd232} : s = 493;
	{8'd22,8'd233} : s = 510;
	{8'd22,8'd234} : s = 1;
	{8'd22,8'd235} : s = 18;
	{8'd22,8'd236} : s = 17;
	{8'd22,8'd237} : s = 82;
	{8'd22,8'd238} : s = 12;
	{8'd22,8'd239} : s = 81;
	{8'd22,8'd240} : s = 76;
	{8'd22,8'd241} : s = 195;
	{8'd22,8'd242} : s = 10;
	{8'd22,8'd243} : s = 74;
	{8'd22,8'd244} : s = 73;
	{8'd22,8'd245} : s = 184;
	{8'd22,8'd246} : s = 70;
	{8'd22,8'd247} : s = 180;
	{8'd22,8'd248} : s = 178;
	{8'd22,8'd249} : s = 314;
	{8'd22,8'd250} : s = 9;
	{8'd22,8'd251} : s = 69;
	{8'd22,8'd252} : s = 67;
	{8'd22,8'd253} : s = 177;
	{8'd22,8'd254} : s = 56;
	{8'd22,8'd255} : s = 172;
	{8'd23,8'd0} : s = 464;
	{8'd23,8'd1} : s = 160;
	{8'd23,8'd2} : s = 352;
	{8'd23,8'd3} : s = 336;
	{8'd23,8'd4} : s = 456;
	{8'd23,8'd5} : s = 328;
	{8'd23,8'd6} : s = 452;
	{8'd23,8'd7} : s = 450;
	{8'd23,8'd8} : s = 496;
	{8'd23,8'd9} : s = 16;
	{8'd23,8'd10} : s = 144;
	{8'd23,8'd11} : s = 136;
	{8'd23,8'd12} : s = 324;
	{8'd23,8'd13} : s = 132;
	{8'd23,8'd14} : s = 322;
	{8'd23,8'd15} : s = 321;
	{8'd23,8'd16} : s = 449;
	{8'd23,8'd17} : s = 130;
	{8'd23,8'd18} : s = 304;
	{8'd23,8'd19} : s = 296;
	{8'd23,8'd20} : s = 432;
	{8'd23,8'd21} : s = 292;
	{8'd23,8'd22} : s = 424;
	{8'd23,8'd23} : s = 420;
	{8'd23,8'd24} : s = 488;
	{8'd23,8'd25} : s = 129;
	{8'd23,8'd26} : s = 290;
	{8'd23,8'd27} : s = 289;
	{8'd23,8'd28} : s = 418;
	{8'd23,8'd29} : s = 280;
	{8'd23,8'd30} : s = 417;
	{8'd23,8'd31} : s = 408;
	{8'd23,8'd32} : s = 484;
	{8'd23,8'd33} : s = 276;
	{8'd23,8'd34} : s = 404;
	{8'd23,8'd35} : s = 402;
	{8'd23,8'd36} : s = 482;
	{8'd23,8'd37} : s = 401;
	{8'd23,8'd38} : s = 481;
	{8'd23,8'd39} : s = 472;
	{8'd23,8'd40} : s = 504;
	{8'd23,8'd41} : s = 4;
	{8'd23,8'd42} : s = 96;
	{8'd23,8'd43} : s = 80;
	{8'd23,8'd44} : s = 274;
	{8'd23,8'd45} : s = 72;
	{8'd23,8'd46} : s = 273;
	{8'd23,8'd47} : s = 268;
	{8'd23,8'd48} : s = 396;
	{8'd23,8'd49} : s = 68;
	{8'd23,8'd50} : s = 266;
	{8'd23,8'd51} : s = 265;
	{8'd23,8'd52} : s = 394;
	{8'd23,8'd53} : s = 262;
	{8'd23,8'd54} : s = 393;
	{8'd23,8'd55} : s = 390;
	{8'd23,8'd56} : s = 468;
	{8'd23,8'd57} : s = 66;
	{8'd23,8'd58} : s = 261;
	{8'd23,8'd59} : s = 259;
	{8'd23,8'd60} : s = 389;
	{8'd23,8'd61} : s = 224;
	{8'd23,8'd62} : s = 387;
	{8'd23,8'd63} : s = 368;
	{8'd23,8'd64} : s = 466;
	{8'd23,8'd65} : s = 208;
	{8'd23,8'd66} : s = 360;
	{8'd23,8'd67} : s = 356;
	{8'd23,8'd68} : s = 465;
	{8'd23,8'd69} : s = 354;
	{8'd23,8'd70} : s = 460;
	{8'd23,8'd71} : s = 458;
	{8'd23,8'd72} : s = 500;
	{8'd23,8'd73} : s = 65;
	{8'd23,8'd74} : s = 200;
	{8'd23,8'd75} : s = 196;
	{8'd23,8'd76} : s = 353;
	{8'd23,8'd77} : s = 194;
	{8'd23,8'd78} : s = 344;
	{8'd23,8'd79} : s = 340;
	{8'd23,8'd80} : s = 457;
	{8'd23,8'd81} : s = 193;
	{8'd23,8'd82} : s = 338;
	{8'd23,8'd83} : s = 337;
	{8'd23,8'd84} : s = 454;
	{8'd23,8'd85} : s = 332;
	{8'd23,8'd86} : s = 453;
	{8'd23,8'd87} : s = 451;
	{8'd23,8'd88} : s = 498;
	{8'd23,8'd89} : s = 176;
	{8'd23,8'd90} : s = 330;
	{8'd23,8'd91} : s = 329;
	{8'd23,8'd92} : s = 440;
	{8'd23,8'd93} : s = 326;
	{8'd23,8'd94} : s = 436;
	{8'd23,8'd95} : s = 434;
	{8'd23,8'd96} : s = 497;
	{8'd23,8'd97} : s = 325;
	{8'd23,8'd98} : s = 433;
	{8'd23,8'd99} : s = 428;
	{8'd23,8'd100} : s = 492;
	{8'd23,8'd101} : s = 426;
	{8'd23,8'd102} : s = 490;
	{8'd23,8'd103} : s = 489;
	{8'd23,8'd104} : s = 508;
	{8'd23,8'd105} : s = 2;
	{8'd23,8'd106} : s = 48;
	{8'd23,8'd107} : s = 40;
	{8'd23,8'd108} : s = 168;
	{8'd23,8'd109} : s = 36;
	{8'd23,8'd110} : s = 164;
	{8'd23,8'd111} : s = 162;
	{8'd23,8'd112} : s = 323;
	{8'd23,8'd113} : s = 34;
	{8'd23,8'd114} : s = 161;
	{8'd23,8'd115} : s = 152;
	{8'd23,8'd116} : s = 312;
	{8'd23,8'd117} : s = 148;
	{8'd23,8'd118} : s = 308;
	{8'd23,8'd119} : s = 306;
	{8'd23,8'd120} : s = 425;
	{8'd23,8'd121} : s = 33;
	{8'd23,8'd122} : s = 146;
	{8'd23,8'd123} : s = 145;
	{8'd23,8'd124} : s = 305;
	{8'd23,8'd125} : s = 140;
	{8'd23,8'd126} : s = 300;
	{8'd23,8'd127} : s = 298;
	{8'd23,8'd128} : s = 422;
	{8'd23,8'd129} : s = 138;
	{8'd23,8'd130} : s = 297;
	{8'd23,8'd131} : s = 294;
	{8'd23,8'd132} : s = 421;
	{8'd23,8'd133} : s = 293;
	{8'd23,8'd134} : s = 419;
	{8'd23,8'd135} : s = 412;
	{8'd23,8'd136} : s = 486;
	{8'd23,8'd137} : s = 24;
	{8'd23,8'd138} : s = 137;
	{8'd23,8'd139} : s = 134;
	{8'd23,8'd140} : s = 291;
	{8'd23,8'd141} : s = 133;
	{8'd23,8'd142} : s = 284;
	{8'd23,8'd143} : s = 282;
	{8'd23,8'd144} : s = 410;
	{8'd23,8'd145} : s = 131;
	{8'd23,8'd146} : s = 281;
	{8'd23,8'd147} : s = 278;
	{8'd23,8'd148} : s = 409;
	{8'd23,8'd149} : s = 277;
	{8'd23,8'd150} : s = 406;
	{8'd23,8'd151} : s = 405;
	{8'd23,8'd152} : s = 485;
	{8'd23,8'd153} : s = 112;
	{8'd23,8'd154} : s = 275;
	{8'd23,8'd155} : s = 270;
	{8'd23,8'd156} : s = 403;
	{8'd23,8'd157} : s = 269;
	{8'd23,8'd158} : s = 398;
	{8'd23,8'd159} : s = 397;
	{8'd23,8'd160} : s = 483;
	{8'd23,8'd161} : s = 267;
	{8'd23,8'd162} : s = 395;
	{8'd23,8'd163} : s = 391;
	{8'd23,8'd164} : s = 476;
	{8'd23,8'd165} : s = 376;
	{8'd23,8'd166} : s = 474;
	{8'd23,8'd167} : s = 473;
	{8'd23,8'd168} : s = 506;
	{8'd23,8'd169} : s = 20;
	{8'd23,8'd170} : s = 104;
	{8'd23,8'd171} : s = 100;
	{8'd23,8'd172} : s = 263;
	{8'd23,8'd173} : s = 98;
	{8'd23,8'd174} : s = 240;
	{8'd23,8'd175} : s = 232;
	{8'd23,8'd176} : s = 372;
	{8'd23,8'd177} : s = 97;
	{8'd23,8'd178} : s = 228;
	{8'd23,8'd179} : s = 226;
	{8'd23,8'd180} : s = 370;
	{8'd23,8'd181} : s = 225;
	{8'd23,8'd182} : s = 369;
	{8'd23,8'd183} : s = 364;
	{8'd23,8'd184} : s = 470;
	{8'd23,8'd185} : s = 88;
	{8'd23,8'd186} : s = 216;
	{8'd23,8'd187} : s = 212;
	{8'd23,8'd188} : s = 362;
	{8'd23,8'd189} : s = 210;
	{8'd23,8'd190} : s = 361;
	{8'd23,8'd191} : s = 358;
	{8'd23,8'd192} : s = 469;
	{8'd23,8'd193} : s = 209;
	{8'd23,8'd194} : s = 357;
	{8'd23,8'd195} : s = 355;
	{8'd23,8'd196} : s = 467;
	{8'd23,8'd197} : s = 348;
	{8'd23,8'd198} : s = 462;
	{8'd23,8'd199} : s = 461;
	{8'd23,8'd200} : s = 505;
	{8'd23,8'd201} : s = 84;
	{8'd23,8'd202} : s = 204;
	{8'd23,8'd203} : s = 202;
	{8'd23,8'd204} : s = 346;
	{8'd23,8'd205} : s = 201;
	{8'd23,8'd206} : s = 345;
	{8'd23,8'd207} : s = 342;
	{8'd23,8'd208} : s = 459;
	{8'd23,8'd209} : s = 198;
	{8'd23,8'd210} : s = 341;
	{8'd23,8'd211} : s = 339;
	{8'd23,8'd212} : s = 455;
	{8'd23,8'd213} : s = 334;
	{8'd23,8'd214} : s = 444;
	{8'd23,8'd215} : s = 442;
	{8'd23,8'd216} : s = 502;
	{8'd23,8'd217} : s = 197;
	{8'd23,8'd218} : s = 333;
	{8'd23,8'd219} : s = 331;
	{8'd23,8'd220} : s = 441;
	{8'd23,8'd221} : s = 327;
	{8'd23,8'd222} : s = 438;
	{8'd23,8'd223} : s = 437;
	{8'd23,8'd224} : s = 501;
	{8'd23,8'd225} : s = 316;
	{8'd23,8'd226} : s = 435;
	{8'd23,8'd227} : s = 430;
	{8'd23,8'd228} : s = 499;
	{8'd23,8'd229} : s = 429;
	{8'd23,8'd230} : s = 494;
	{8'd23,8'd231} : s = 493;
	{8'd23,8'd232} : s = 510;
	{8'd23,8'd233} : s = 1;
	{8'd23,8'd234} : s = 18;
	{8'd23,8'd235} : s = 17;
	{8'd23,8'd236} : s = 82;
	{8'd23,8'd237} : s = 12;
	{8'd23,8'd238} : s = 81;
	{8'd23,8'd239} : s = 76;
	{8'd23,8'd240} : s = 195;
	{8'd23,8'd241} : s = 10;
	{8'd23,8'd242} : s = 74;
	{8'd23,8'd243} : s = 73;
	{8'd23,8'd244} : s = 184;
	{8'd23,8'd245} : s = 70;
	{8'd23,8'd246} : s = 180;
	{8'd23,8'd247} : s = 178;
	{8'd23,8'd248} : s = 314;
	{8'd23,8'd249} : s = 9;
	{8'd23,8'd250} : s = 69;
	{8'd23,8'd251} : s = 67;
	{8'd23,8'd252} : s = 177;
	{8'd23,8'd253} : s = 56;
	{8'd23,8'd254} : s = 172;
	{8'd23,8'd255} : s = 170;
	{8'd24,8'd0} : s = 160;
	{8'd24,8'd1} : s = 352;
	{8'd24,8'd2} : s = 336;
	{8'd24,8'd3} : s = 456;
	{8'd24,8'd4} : s = 328;
	{8'd24,8'd5} : s = 452;
	{8'd24,8'd6} : s = 450;
	{8'd24,8'd7} : s = 496;
	{8'd24,8'd8} : s = 16;
	{8'd24,8'd9} : s = 144;
	{8'd24,8'd10} : s = 136;
	{8'd24,8'd11} : s = 324;
	{8'd24,8'd12} : s = 132;
	{8'd24,8'd13} : s = 322;
	{8'd24,8'd14} : s = 321;
	{8'd24,8'd15} : s = 449;
	{8'd24,8'd16} : s = 130;
	{8'd24,8'd17} : s = 304;
	{8'd24,8'd18} : s = 296;
	{8'd24,8'd19} : s = 432;
	{8'd24,8'd20} : s = 292;
	{8'd24,8'd21} : s = 424;
	{8'd24,8'd22} : s = 420;
	{8'd24,8'd23} : s = 488;
	{8'd24,8'd24} : s = 129;
	{8'd24,8'd25} : s = 290;
	{8'd24,8'd26} : s = 289;
	{8'd24,8'd27} : s = 418;
	{8'd24,8'd28} : s = 280;
	{8'd24,8'd29} : s = 417;
	{8'd24,8'd30} : s = 408;
	{8'd24,8'd31} : s = 484;
	{8'd24,8'd32} : s = 276;
	{8'd24,8'd33} : s = 404;
	{8'd24,8'd34} : s = 402;
	{8'd24,8'd35} : s = 482;
	{8'd24,8'd36} : s = 401;
	{8'd24,8'd37} : s = 481;
	{8'd24,8'd38} : s = 472;
	{8'd24,8'd39} : s = 504;
	{8'd24,8'd40} : s = 4;
	{8'd24,8'd41} : s = 96;
	{8'd24,8'd42} : s = 80;
	{8'd24,8'd43} : s = 274;
	{8'd24,8'd44} : s = 72;
	{8'd24,8'd45} : s = 273;
	{8'd24,8'd46} : s = 268;
	{8'd24,8'd47} : s = 396;
	{8'd24,8'd48} : s = 68;
	{8'd24,8'd49} : s = 266;
	{8'd24,8'd50} : s = 265;
	{8'd24,8'd51} : s = 394;
	{8'd24,8'd52} : s = 262;
	{8'd24,8'd53} : s = 393;
	{8'd24,8'd54} : s = 390;
	{8'd24,8'd55} : s = 468;
	{8'd24,8'd56} : s = 66;
	{8'd24,8'd57} : s = 261;
	{8'd24,8'd58} : s = 259;
	{8'd24,8'd59} : s = 389;
	{8'd24,8'd60} : s = 224;
	{8'd24,8'd61} : s = 387;
	{8'd24,8'd62} : s = 368;
	{8'd24,8'd63} : s = 466;
	{8'd24,8'd64} : s = 208;
	{8'd24,8'd65} : s = 360;
	{8'd24,8'd66} : s = 356;
	{8'd24,8'd67} : s = 465;
	{8'd24,8'd68} : s = 354;
	{8'd24,8'd69} : s = 460;
	{8'd24,8'd70} : s = 458;
	{8'd24,8'd71} : s = 500;
	{8'd24,8'd72} : s = 65;
	{8'd24,8'd73} : s = 200;
	{8'd24,8'd74} : s = 196;
	{8'd24,8'd75} : s = 353;
	{8'd24,8'd76} : s = 194;
	{8'd24,8'd77} : s = 344;
	{8'd24,8'd78} : s = 340;
	{8'd24,8'd79} : s = 457;
	{8'd24,8'd80} : s = 193;
	{8'd24,8'd81} : s = 338;
	{8'd24,8'd82} : s = 337;
	{8'd24,8'd83} : s = 454;
	{8'd24,8'd84} : s = 332;
	{8'd24,8'd85} : s = 453;
	{8'd24,8'd86} : s = 451;
	{8'd24,8'd87} : s = 498;
	{8'd24,8'd88} : s = 176;
	{8'd24,8'd89} : s = 330;
	{8'd24,8'd90} : s = 329;
	{8'd24,8'd91} : s = 440;
	{8'd24,8'd92} : s = 326;
	{8'd24,8'd93} : s = 436;
	{8'd24,8'd94} : s = 434;
	{8'd24,8'd95} : s = 497;
	{8'd24,8'd96} : s = 325;
	{8'd24,8'd97} : s = 433;
	{8'd24,8'd98} : s = 428;
	{8'd24,8'd99} : s = 492;
	{8'd24,8'd100} : s = 426;
	{8'd24,8'd101} : s = 490;
	{8'd24,8'd102} : s = 489;
	{8'd24,8'd103} : s = 508;
	{8'd24,8'd104} : s = 2;
	{8'd24,8'd105} : s = 48;
	{8'd24,8'd106} : s = 40;
	{8'd24,8'd107} : s = 168;
	{8'd24,8'd108} : s = 36;
	{8'd24,8'd109} : s = 164;
	{8'd24,8'd110} : s = 162;
	{8'd24,8'd111} : s = 323;
	{8'd24,8'd112} : s = 34;
	{8'd24,8'd113} : s = 161;
	{8'd24,8'd114} : s = 152;
	{8'd24,8'd115} : s = 312;
	{8'd24,8'd116} : s = 148;
	{8'd24,8'd117} : s = 308;
	{8'd24,8'd118} : s = 306;
	{8'd24,8'd119} : s = 425;
	{8'd24,8'd120} : s = 33;
	{8'd24,8'd121} : s = 146;
	{8'd24,8'd122} : s = 145;
	{8'd24,8'd123} : s = 305;
	{8'd24,8'd124} : s = 140;
	{8'd24,8'd125} : s = 300;
	{8'd24,8'd126} : s = 298;
	{8'd24,8'd127} : s = 422;
	{8'd24,8'd128} : s = 138;
	{8'd24,8'd129} : s = 297;
	{8'd24,8'd130} : s = 294;
	{8'd24,8'd131} : s = 421;
	{8'd24,8'd132} : s = 293;
	{8'd24,8'd133} : s = 419;
	{8'd24,8'd134} : s = 412;
	{8'd24,8'd135} : s = 486;
	{8'd24,8'd136} : s = 24;
	{8'd24,8'd137} : s = 137;
	{8'd24,8'd138} : s = 134;
	{8'd24,8'd139} : s = 291;
	{8'd24,8'd140} : s = 133;
	{8'd24,8'd141} : s = 284;
	{8'd24,8'd142} : s = 282;
	{8'd24,8'd143} : s = 410;
	{8'd24,8'd144} : s = 131;
	{8'd24,8'd145} : s = 281;
	{8'd24,8'd146} : s = 278;
	{8'd24,8'd147} : s = 409;
	{8'd24,8'd148} : s = 277;
	{8'd24,8'd149} : s = 406;
	{8'd24,8'd150} : s = 405;
	{8'd24,8'd151} : s = 485;
	{8'd24,8'd152} : s = 112;
	{8'd24,8'd153} : s = 275;
	{8'd24,8'd154} : s = 270;
	{8'd24,8'd155} : s = 403;
	{8'd24,8'd156} : s = 269;
	{8'd24,8'd157} : s = 398;
	{8'd24,8'd158} : s = 397;
	{8'd24,8'd159} : s = 483;
	{8'd24,8'd160} : s = 267;
	{8'd24,8'd161} : s = 395;
	{8'd24,8'd162} : s = 391;
	{8'd24,8'd163} : s = 476;
	{8'd24,8'd164} : s = 376;
	{8'd24,8'd165} : s = 474;
	{8'd24,8'd166} : s = 473;
	{8'd24,8'd167} : s = 506;
	{8'd24,8'd168} : s = 20;
	{8'd24,8'd169} : s = 104;
	{8'd24,8'd170} : s = 100;
	{8'd24,8'd171} : s = 263;
	{8'd24,8'd172} : s = 98;
	{8'd24,8'd173} : s = 240;
	{8'd24,8'd174} : s = 232;
	{8'd24,8'd175} : s = 372;
	{8'd24,8'd176} : s = 97;
	{8'd24,8'd177} : s = 228;
	{8'd24,8'd178} : s = 226;
	{8'd24,8'd179} : s = 370;
	{8'd24,8'd180} : s = 225;
	{8'd24,8'd181} : s = 369;
	{8'd24,8'd182} : s = 364;
	{8'd24,8'd183} : s = 470;
	{8'd24,8'd184} : s = 88;
	{8'd24,8'd185} : s = 216;
	{8'd24,8'd186} : s = 212;
	{8'd24,8'd187} : s = 362;
	{8'd24,8'd188} : s = 210;
	{8'd24,8'd189} : s = 361;
	{8'd24,8'd190} : s = 358;
	{8'd24,8'd191} : s = 469;
	{8'd24,8'd192} : s = 209;
	{8'd24,8'd193} : s = 357;
	{8'd24,8'd194} : s = 355;
	{8'd24,8'd195} : s = 467;
	{8'd24,8'd196} : s = 348;
	{8'd24,8'd197} : s = 462;
	{8'd24,8'd198} : s = 461;
	{8'd24,8'd199} : s = 505;
	{8'd24,8'd200} : s = 84;
	{8'd24,8'd201} : s = 204;
	{8'd24,8'd202} : s = 202;
	{8'd24,8'd203} : s = 346;
	{8'd24,8'd204} : s = 201;
	{8'd24,8'd205} : s = 345;
	{8'd24,8'd206} : s = 342;
	{8'd24,8'd207} : s = 459;
	{8'd24,8'd208} : s = 198;
	{8'd24,8'd209} : s = 341;
	{8'd24,8'd210} : s = 339;
	{8'd24,8'd211} : s = 455;
	{8'd24,8'd212} : s = 334;
	{8'd24,8'd213} : s = 444;
	{8'd24,8'd214} : s = 442;
	{8'd24,8'd215} : s = 502;
	{8'd24,8'd216} : s = 197;
	{8'd24,8'd217} : s = 333;
	{8'd24,8'd218} : s = 331;
	{8'd24,8'd219} : s = 441;
	{8'd24,8'd220} : s = 327;
	{8'd24,8'd221} : s = 438;
	{8'd24,8'd222} : s = 437;
	{8'd24,8'd223} : s = 501;
	{8'd24,8'd224} : s = 316;
	{8'd24,8'd225} : s = 435;
	{8'd24,8'd226} : s = 430;
	{8'd24,8'd227} : s = 499;
	{8'd24,8'd228} : s = 429;
	{8'd24,8'd229} : s = 494;
	{8'd24,8'd230} : s = 493;
	{8'd24,8'd231} : s = 510;
	{8'd24,8'd232} : s = 1;
	{8'd24,8'd233} : s = 18;
	{8'd24,8'd234} : s = 17;
	{8'd24,8'd235} : s = 82;
	{8'd24,8'd236} : s = 12;
	{8'd24,8'd237} : s = 81;
	{8'd24,8'd238} : s = 76;
	{8'd24,8'd239} : s = 195;
	{8'd24,8'd240} : s = 10;
	{8'd24,8'd241} : s = 74;
	{8'd24,8'd242} : s = 73;
	{8'd24,8'd243} : s = 184;
	{8'd24,8'd244} : s = 70;
	{8'd24,8'd245} : s = 180;
	{8'd24,8'd246} : s = 178;
	{8'd24,8'd247} : s = 314;
	{8'd24,8'd248} : s = 9;
	{8'd24,8'd249} : s = 69;
	{8'd24,8'd250} : s = 67;
	{8'd24,8'd251} : s = 177;
	{8'd24,8'd252} : s = 56;
	{8'd24,8'd253} : s = 172;
	{8'd24,8'd254} : s = 170;
	{8'd24,8'd255} : s = 313;
	{8'd25,8'd0} : s = 352;
	{8'd25,8'd1} : s = 336;
	{8'd25,8'd2} : s = 456;
	{8'd25,8'd3} : s = 328;
	{8'd25,8'd4} : s = 452;
	{8'd25,8'd5} : s = 450;
	{8'd25,8'd6} : s = 496;
	{8'd25,8'd7} : s = 16;
	{8'd25,8'd8} : s = 144;
	{8'd25,8'd9} : s = 136;
	{8'd25,8'd10} : s = 324;
	{8'd25,8'd11} : s = 132;
	{8'd25,8'd12} : s = 322;
	{8'd25,8'd13} : s = 321;
	{8'd25,8'd14} : s = 449;
	{8'd25,8'd15} : s = 130;
	{8'd25,8'd16} : s = 304;
	{8'd25,8'd17} : s = 296;
	{8'd25,8'd18} : s = 432;
	{8'd25,8'd19} : s = 292;
	{8'd25,8'd20} : s = 424;
	{8'd25,8'd21} : s = 420;
	{8'd25,8'd22} : s = 488;
	{8'd25,8'd23} : s = 129;
	{8'd25,8'd24} : s = 290;
	{8'd25,8'd25} : s = 289;
	{8'd25,8'd26} : s = 418;
	{8'd25,8'd27} : s = 280;
	{8'd25,8'd28} : s = 417;
	{8'd25,8'd29} : s = 408;
	{8'd25,8'd30} : s = 484;
	{8'd25,8'd31} : s = 276;
	{8'd25,8'd32} : s = 404;
	{8'd25,8'd33} : s = 402;
	{8'd25,8'd34} : s = 482;
	{8'd25,8'd35} : s = 401;
	{8'd25,8'd36} : s = 481;
	{8'd25,8'd37} : s = 472;
	{8'd25,8'd38} : s = 504;
	{8'd25,8'd39} : s = 4;
	{8'd25,8'd40} : s = 96;
	{8'd25,8'd41} : s = 80;
	{8'd25,8'd42} : s = 274;
	{8'd25,8'd43} : s = 72;
	{8'd25,8'd44} : s = 273;
	{8'd25,8'd45} : s = 268;
	{8'd25,8'd46} : s = 396;
	{8'd25,8'd47} : s = 68;
	{8'd25,8'd48} : s = 266;
	{8'd25,8'd49} : s = 265;
	{8'd25,8'd50} : s = 394;
	{8'd25,8'd51} : s = 262;
	{8'd25,8'd52} : s = 393;
	{8'd25,8'd53} : s = 390;
	{8'd25,8'd54} : s = 468;
	{8'd25,8'd55} : s = 66;
	{8'd25,8'd56} : s = 261;
	{8'd25,8'd57} : s = 259;
	{8'd25,8'd58} : s = 389;
	{8'd25,8'd59} : s = 224;
	{8'd25,8'd60} : s = 387;
	{8'd25,8'd61} : s = 368;
	{8'd25,8'd62} : s = 466;
	{8'd25,8'd63} : s = 208;
	{8'd25,8'd64} : s = 360;
	{8'd25,8'd65} : s = 356;
	{8'd25,8'd66} : s = 465;
	{8'd25,8'd67} : s = 354;
	{8'd25,8'd68} : s = 460;
	{8'd25,8'd69} : s = 458;
	{8'd25,8'd70} : s = 500;
	{8'd25,8'd71} : s = 65;
	{8'd25,8'd72} : s = 200;
	{8'd25,8'd73} : s = 196;
	{8'd25,8'd74} : s = 353;
	{8'd25,8'd75} : s = 194;
	{8'd25,8'd76} : s = 344;
	{8'd25,8'd77} : s = 340;
	{8'd25,8'd78} : s = 457;
	{8'd25,8'd79} : s = 193;
	{8'd25,8'd80} : s = 338;
	{8'd25,8'd81} : s = 337;
	{8'd25,8'd82} : s = 454;
	{8'd25,8'd83} : s = 332;
	{8'd25,8'd84} : s = 453;
	{8'd25,8'd85} : s = 451;
	{8'd25,8'd86} : s = 498;
	{8'd25,8'd87} : s = 176;
	{8'd25,8'd88} : s = 330;
	{8'd25,8'd89} : s = 329;
	{8'd25,8'd90} : s = 440;
	{8'd25,8'd91} : s = 326;
	{8'd25,8'd92} : s = 436;
	{8'd25,8'd93} : s = 434;
	{8'd25,8'd94} : s = 497;
	{8'd25,8'd95} : s = 325;
	{8'd25,8'd96} : s = 433;
	{8'd25,8'd97} : s = 428;
	{8'd25,8'd98} : s = 492;
	{8'd25,8'd99} : s = 426;
	{8'd25,8'd100} : s = 490;
	{8'd25,8'd101} : s = 489;
	{8'd25,8'd102} : s = 508;
	{8'd25,8'd103} : s = 2;
	{8'd25,8'd104} : s = 48;
	{8'd25,8'd105} : s = 40;
	{8'd25,8'd106} : s = 168;
	{8'd25,8'd107} : s = 36;
	{8'd25,8'd108} : s = 164;
	{8'd25,8'd109} : s = 162;
	{8'd25,8'd110} : s = 323;
	{8'd25,8'd111} : s = 34;
	{8'd25,8'd112} : s = 161;
	{8'd25,8'd113} : s = 152;
	{8'd25,8'd114} : s = 312;
	{8'd25,8'd115} : s = 148;
	{8'd25,8'd116} : s = 308;
	{8'd25,8'd117} : s = 306;
	{8'd25,8'd118} : s = 425;
	{8'd25,8'd119} : s = 33;
	{8'd25,8'd120} : s = 146;
	{8'd25,8'd121} : s = 145;
	{8'd25,8'd122} : s = 305;
	{8'd25,8'd123} : s = 140;
	{8'd25,8'd124} : s = 300;
	{8'd25,8'd125} : s = 298;
	{8'd25,8'd126} : s = 422;
	{8'd25,8'd127} : s = 138;
	{8'd25,8'd128} : s = 297;
	{8'd25,8'd129} : s = 294;
	{8'd25,8'd130} : s = 421;
	{8'd25,8'd131} : s = 293;
	{8'd25,8'd132} : s = 419;
	{8'd25,8'd133} : s = 412;
	{8'd25,8'd134} : s = 486;
	{8'd25,8'd135} : s = 24;
	{8'd25,8'd136} : s = 137;
	{8'd25,8'd137} : s = 134;
	{8'd25,8'd138} : s = 291;
	{8'd25,8'd139} : s = 133;
	{8'd25,8'd140} : s = 284;
	{8'd25,8'd141} : s = 282;
	{8'd25,8'd142} : s = 410;
	{8'd25,8'd143} : s = 131;
	{8'd25,8'd144} : s = 281;
	{8'd25,8'd145} : s = 278;
	{8'd25,8'd146} : s = 409;
	{8'd25,8'd147} : s = 277;
	{8'd25,8'd148} : s = 406;
	{8'd25,8'd149} : s = 405;
	{8'd25,8'd150} : s = 485;
	{8'd25,8'd151} : s = 112;
	{8'd25,8'd152} : s = 275;
	{8'd25,8'd153} : s = 270;
	{8'd25,8'd154} : s = 403;
	{8'd25,8'd155} : s = 269;
	{8'd25,8'd156} : s = 398;
	{8'd25,8'd157} : s = 397;
	{8'd25,8'd158} : s = 483;
	{8'd25,8'd159} : s = 267;
	{8'd25,8'd160} : s = 395;
	{8'd25,8'd161} : s = 391;
	{8'd25,8'd162} : s = 476;
	{8'd25,8'd163} : s = 376;
	{8'd25,8'd164} : s = 474;
	{8'd25,8'd165} : s = 473;
	{8'd25,8'd166} : s = 506;
	{8'd25,8'd167} : s = 20;
	{8'd25,8'd168} : s = 104;
	{8'd25,8'd169} : s = 100;
	{8'd25,8'd170} : s = 263;
	{8'd25,8'd171} : s = 98;
	{8'd25,8'd172} : s = 240;
	{8'd25,8'd173} : s = 232;
	{8'd25,8'd174} : s = 372;
	{8'd25,8'd175} : s = 97;
	{8'd25,8'd176} : s = 228;
	{8'd25,8'd177} : s = 226;
	{8'd25,8'd178} : s = 370;
	{8'd25,8'd179} : s = 225;
	{8'd25,8'd180} : s = 369;
	{8'd25,8'd181} : s = 364;
	{8'd25,8'd182} : s = 470;
	{8'd25,8'd183} : s = 88;
	{8'd25,8'd184} : s = 216;
	{8'd25,8'd185} : s = 212;
	{8'd25,8'd186} : s = 362;
	{8'd25,8'd187} : s = 210;
	{8'd25,8'd188} : s = 361;
	{8'd25,8'd189} : s = 358;
	{8'd25,8'd190} : s = 469;
	{8'd25,8'd191} : s = 209;
	{8'd25,8'd192} : s = 357;
	{8'd25,8'd193} : s = 355;
	{8'd25,8'd194} : s = 467;
	{8'd25,8'd195} : s = 348;
	{8'd25,8'd196} : s = 462;
	{8'd25,8'd197} : s = 461;
	{8'd25,8'd198} : s = 505;
	{8'd25,8'd199} : s = 84;
	{8'd25,8'd200} : s = 204;
	{8'd25,8'd201} : s = 202;
	{8'd25,8'd202} : s = 346;
	{8'd25,8'd203} : s = 201;
	{8'd25,8'd204} : s = 345;
	{8'd25,8'd205} : s = 342;
	{8'd25,8'd206} : s = 459;
	{8'd25,8'd207} : s = 198;
	{8'd25,8'd208} : s = 341;
	{8'd25,8'd209} : s = 339;
	{8'd25,8'd210} : s = 455;
	{8'd25,8'd211} : s = 334;
	{8'd25,8'd212} : s = 444;
	{8'd25,8'd213} : s = 442;
	{8'd25,8'd214} : s = 502;
	{8'd25,8'd215} : s = 197;
	{8'd25,8'd216} : s = 333;
	{8'd25,8'd217} : s = 331;
	{8'd25,8'd218} : s = 441;
	{8'd25,8'd219} : s = 327;
	{8'd25,8'd220} : s = 438;
	{8'd25,8'd221} : s = 437;
	{8'd25,8'd222} : s = 501;
	{8'd25,8'd223} : s = 316;
	{8'd25,8'd224} : s = 435;
	{8'd25,8'd225} : s = 430;
	{8'd25,8'd226} : s = 499;
	{8'd25,8'd227} : s = 429;
	{8'd25,8'd228} : s = 494;
	{8'd25,8'd229} : s = 493;
	{8'd25,8'd230} : s = 510;
	{8'd25,8'd231} : s = 1;
	{8'd25,8'd232} : s = 18;
	{8'd25,8'd233} : s = 17;
	{8'd25,8'd234} : s = 82;
	{8'd25,8'd235} : s = 12;
	{8'd25,8'd236} : s = 81;
	{8'd25,8'd237} : s = 76;
	{8'd25,8'd238} : s = 195;
	{8'd25,8'd239} : s = 10;
	{8'd25,8'd240} : s = 74;
	{8'd25,8'd241} : s = 73;
	{8'd25,8'd242} : s = 184;
	{8'd25,8'd243} : s = 70;
	{8'd25,8'd244} : s = 180;
	{8'd25,8'd245} : s = 178;
	{8'd25,8'd246} : s = 314;
	{8'd25,8'd247} : s = 9;
	{8'd25,8'd248} : s = 69;
	{8'd25,8'd249} : s = 67;
	{8'd25,8'd250} : s = 177;
	{8'd25,8'd251} : s = 56;
	{8'd25,8'd252} : s = 172;
	{8'd25,8'd253} : s = 170;
	{8'd25,8'd254} : s = 313;
	{8'd25,8'd255} : s = 52;
	{8'd26,8'd0} : s = 336;
	{8'd26,8'd1} : s = 456;
	{8'd26,8'd2} : s = 328;
	{8'd26,8'd3} : s = 452;
	{8'd26,8'd4} : s = 450;
	{8'd26,8'd5} : s = 496;
	{8'd26,8'd6} : s = 16;
	{8'd26,8'd7} : s = 144;
	{8'd26,8'd8} : s = 136;
	{8'd26,8'd9} : s = 324;
	{8'd26,8'd10} : s = 132;
	{8'd26,8'd11} : s = 322;
	{8'd26,8'd12} : s = 321;
	{8'd26,8'd13} : s = 449;
	{8'd26,8'd14} : s = 130;
	{8'd26,8'd15} : s = 304;
	{8'd26,8'd16} : s = 296;
	{8'd26,8'd17} : s = 432;
	{8'd26,8'd18} : s = 292;
	{8'd26,8'd19} : s = 424;
	{8'd26,8'd20} : s = 420;
	{8'd26,8'd21} : s = 488;
	{8'd26,8'd22} : s = 129;
	{8'd26,8'd23} : s = 290;
	{8'd26,8'd24} : s = 289;
	{8'd26,8'd25} : s = 418;
	{8'd26,8'd26} : s = 280;
	{8'd26,8'd27} : s = 417;
	{8'd26,8'd28} : s = 408;
	{8'd26,8'd29} : s = 484;
	{8'd26,8'd30} : s = 276;
	{8'd26,8'd31} : s = 404;
	{8'd26,8'd32} : s = 402;
	{8'd26,8'd33} : s = 482;
	{8'd26,8'd34} : s = 401;
	{8'd26,8'd35} : s = 481;
	{8'd26,8'd36} : s = 472;
	{8'd26,8'd37} : s = 504;
	{8'd26,8'd38} : s = 4;
	{8'd26,8'd39} : s = 96;
	{8'd26,8'd40} : s = 80;
	{8'd26,8'd41} : s = 274;
	{8'd26,8'd42} : s = 72;
	{8'd26,8'd43} : s = 273;
	{8'd26,8'd44} : s = 268;
	{8'd26,8'd45} : s = 396;
	{8'd26,8'd46} : s = 68;
	{8'd26,8'd47} : s = 266;
	{8'd26,8'd48} : s = 265;
	{8'd26,8'd49} : s = 394;
	{8'd26,8'd50} : s = 262;
	{8'd26,8'd51} : s = 393;
	{8'd26,8'd52} : s = 390;
	{8'd26,8'd53} : s = 468;
	{8'd26,8'd54} : s = 66;
	{8'd26,8'd55} : s = 261;
	{8'd26,8'd56} : s = 259;
	{8'd26,8'd57} : s = 389;
	{8'd26,8'd58} : s = 224;
	{8'd26,8'd59} : s = 387;
	{8'd26,8'd60} : s = 368;
	{8'd26,8'd61} : s = 466;
	{8'd26,8'd62} : s = 208;
	{8'd26,8'd63} : s = 360;
	{8'd26,8'd64} : s = 356;
	{8'd26,8'd65} : s = 465;
	{8'd26,8'd66} : s = 354;
	{8'd26,8'd67} : s = 460;
	{8'd26,8'd68} : s = 458;
	{8'd26,8'd69} : s = 500;
	{8'd26,8'd70} : s = 65;
	{8'd26,8'd71} : s = 200;
	{8'd26,8'd72} : s = 196;
	{8'd26,8'd73} : s = 353;
	{8'd26,8'd74} : s = 194;
	{8'd26,8'd75} : s = 344;
	{8'd26,8'd76} : s = 340;
	{8'd26,8'd77} : s = 457;
	{8'd26,8'd78} : s = 193;
	{8'd26,8'd79} : s = 338;
	{8'd26,8'd80} : s = 337;
	{8'd26,8'd81} : s = 454;
	{8'd26,8'd82} : s = 332;
	{8'd26,8'd83} : s = 453;
	{8'd26,8'd84} : s = 451;
	{8'd26,8'd85} : s = 498;
	{8'd26,8'd86} : s = 176;
	{8'd26,8'd87} : s = 330;
	{8'd26,8'd88} : s = 329;
	{8'd26,8'd89} : s = 440;
	{8'd26,8'd90} : s = 326;
	{8'd26,8'd91} : s = 436;
	{8'd26,8'd92} : s = 434;
	{8'd26,8'd93} : s = 497;
	{8'd26,8'd94} : s = 325;
	{8'd26,8'd95} : s = 433;
	{8'd26,8'd96} : s = 428;
	{8'd26,8'd97} : s = 492;
	{8'd26,8'd98} : s = 426;
	{8'd26,8'd99} : s = 490;
	{8'd26,8'd100} : s = 489;
	{8'd26,8'd101} : s = 508;
	{8'd26,8'd102} : s = 2;
	{8'd26,8'd103} : s = 48;
	{8'd26,8'd104} : s = 40;
	{8'd26,8'd105} : s = 168;
	{8'd26,8'd106} : s = 36;
	{8'd26,8'd107} : s = 164;
	{8'd26,8'd108} : s = 162;
	{8'd26,8'd109} : s = 323;
	{8'd26,8'd110} : s = 34;
	{8'd26,8'd111} : s = 161;
	{8'd26,8'd112} : s = 152;
	{8'd26,8'd113} : s = 312;
	{8'd26,8'd114} : s = 148;
	{8'd26,8'd115} : s = 308;
	{8'd26,8'd116} : s = 306;
	{8'd26,8'd117} : s = 425;
	{8'd26,8'd118} : s = 33;
	{8'd26,8'd119} : s = 146;
	{8'd26,8'd120} : s = 145;
	{8'd26,8'd121} : s = 305;
	{8'd26,8'd122} : s = 140;
	{8'd26,8'd123} : s = 300;
	{8'd26,8'd124} : s = 298;
	{8'd26,8'd125} : s = 422;
	{8'd26,8'd126} : s = 138;
	{8'd26,8'd127} : s = 297;
	{8'd26,8'd128} : s = 294;
	{8'd26,8'd129} : s = 421;
	{8'd26,8'd130} : s = 293;
	{8'd26,8'd131} : s = 419;
	{8'd26,8'd132} : s = 412;
	{8'd26,8'd133} : s = 486;
	{8'd26,8'd134} : s = 24;
	{8'd26,8'd135} : s = 137;
	{8'd26,8'd136} : s = 134;
	{8'd26,8'd137} : s = 291;
	{8'd26,8'd138} : s = 133;
	{8'd26,8'd139} : s = 284;
	{8'd26,8'd140} : s = 282;
	{8'd26,8'd141} : s = 410;
	{8'd26,8'd142} : s = 131;
	{8'd26,8'd143} : s = 281;
	{8'd26,8'd144} : s = 278;
	{8'd26,8'd145} : s = 409;
	{8'd26,8'd146} : s = 277;
	{8'd26,8'd147} : s = 406;
	{8'd26,8'd148} : s = 405;
	{8'd26,8'd149} : s = 485;
	{8'd26,8'd150} : s = 112;
	{8'd26,8'd151} : s = 275;
	{8'd26,8'd152} : s = 270;
	{8'd26,8'd153} : s = 403;
	{8'd26,8'd154} : s = 269;
	{8'd26,8'd155} : s = 398;
	{8'd26,8'd156} : s = 397;
	{8'd26,8'd157} : s = 483;
	{8'd26,8'd158} : s = 267;
	{8'd26,8'd159} : s = 395;
	{8'd26,8'd160} : s = 391;
	{8'd26,8'd161} : s = 476;
	{8'd26,8'd162} : s = 376;
	{8'd26,8'd163} : s = 474;
	{8'd26,8'd164} : s = 473;
	{8'd26,8'd165} : s = 506;
	{8'd26,8'd166} : s = 20;
	{8'd26,8'd167} : s = 104;
	{8'd26,8'd168} : s = 100;
	{8'd26,8'd169} : s = 263;
	{8'd26,8'd170} : s = 98;
	{8'd26,8'd171} : s = 240;
	{8'd26,8'd172} : s = 232;
	{8'd26,8'd173} : s = 372;
	{8'd26,8'd174} : s = 97;
	{8'd26,8'd175} : s = 228;
	{8'd26,8'd176} : s = 226;
	{8'd26,8'd177} : s = 370;
	{8'd26,8'd178} : s = 225;
	{8'd26,8'd179} : s = 369;
	{8'd26,8'd180} : s = 364;
	{8'd26,8'd181} : s = 470;
	{8'd26,8'd182} : s = 88;
	{8'd26,8'd183} : s = 216;
	{8'd26,8'd184} : s = 212;
	{8'd26,8'd185} : s = 362;
	{8'd26,8'd186} : s = 210;
	{8'd26,8'd187} : s = 361;
	{8'd26,8'd188} : s = 358;
	{8'd26,8'd189} : s = 469;
	{8'd26,8'd190} : s = 209;
	{8'd26,8'd191} : s = 357;
	{8'd26,8'd192} : s = 355;
	{8'd26,8'd193} : s = 467;
	{8'd26,8'd194} : s = 348;
	{8'd26,8'd195} : s = 462;
	{8'd26,8'd196} : s = 461;
	{8'd26,8'd197} : s = 505;
	{8'd26,8'd198} : s = 84;
	{8'd26,8'd199} : s = 204;
	{8'd26,8'd200} : s = 202;
	{8'd26,8'd201} : s = 346;
	{8'd26,8'd202} : s = 201;
	{8'd26,8'd203} : s = 345;
	{8'd26,8'd204} : s = 342;
	{8'd26,8'd205} : s = 459;
	{8'd26,8'd206} : s = 198;
	{8'd26,8'd207} : s = 341;
	{8'd26,8'd208} : s = 339;
	{8'd26,8'd209} : s = 455;
	{8'd26,8'd210} : s = 334;
	{8'd26,8'd211} : s = 444;
	{8'd26,8'd212} : s = 442;
	{8'd26,8'd213} : s = 502;
	{8'd26,8'd214} : s = 197;
	{8'd26,8'd215} : s = 333;
	{8'd26,8'd216} : s = 331;
	{8'd26,8'd217} : s = 441;
	{8'd26,8'd218} : s = 327;
	{8'd26,8'd219} : s = 438;
	{8'd26,8'd220} : s = 437;
	{8'd26,8'd221} : s = 501;
	{8'd26,8'd222} : s = 316;
	{8'd26,8'd223} : s = 435;
	{8'd26,8'd224} : s = 430;
	{8'd26,8'd225} : s = 499;
	{8'd26,8'd226} : s = 429;
	{8'd26,8'd227} : s = 494;
	{8'd26,8'd228} : s = 493;
	{8'd26,8'd229} : s = 510;
	{8'd26,8'd230} : s = 1;
	{8'd26,8'd231} : s = 18;
	{8'd26,8'd232} : s = 17;
	{8'd26,8'd233} : s = 82;
	{8'd26,8'd234} : s = 12;
	{8'd26,8'd235} : s = 81;
	{8'd26,8'd236} : s = 76;
	{8'd26,8'd237} : s = 195;
	{8'd26,8'd238} : s = 10;
	{8'd26,8'd239} : s = 74;
	{8'd26,8'd240} : s = 73;
	{8'd26,8'd241} : s = 184;
	{8'd26,8'd242} : s = 70;
	{8'd26,8'd243} : s = 180;
	{8'd26,8'd244} : s = 178;
	{8'd26,8'd245} : s = 314;
	{8'd26,8'd246} : s = 9;
	{8'd26,8'd247} : s = 69;
	{8'd26,8'd248} : s = 67;
	{8'd26,8'd249} : s = 177;
	{8'd26,8'd250} : s = 56;
	{8'd26,8'd251} : s = 172;
	{8'd26,8'd252} : s = 170;
	{8'd26,8'd253} : s = 313;
	{8'd26,8'd254} : s = 52;
	{8'd26,8'd255} : s = 169;
	{8'd27,8'd0} : s = 456;
	{8'd27,8'd1} : s = 328;
	{8'd27,8'd2} : s = 452;
	{8'd27,8'd3} : s = 450;
	{8'd27,8'd4} : s = 496;
	{8'd27,8'd5} : s = 16;
	{8'd27,8'd6} : s = 144;
	{8'd27,8'd7} : s = 136;
	{8'd27,8'd8} : s = 324;
	{8'd27,8'd9} : s = 132;
	{8'd27,8'd10} : s = 322;
	{8'd27,8'd11} : s = 321;
	{8'd27,8'd12} : s = 449;
	{8'd27,8'd13} : s = 130;
	{8'd27,8'd14} : s = 304;
	{8'd27,8'd15} : s = 296;
	{8'd27,8'd16} : s = 432;
	{8'd27,8'd17} : s = 292;
	{8'd27,8'd18} : s = 424;
	{8'd27,8'd19} : s = 420;
	{8'd27,8'd20} : s = 488;
	{8'd27,8'd21} : s = 129;
	{8'd27,8'd22} : s = 290;
	{8'd27,8'd23} : s = 289;
	{8'd27,8'd24} : s = 418;
	{8'd27,8'd25} : s = 280;
	{8'd27,8'd26} : s = 417;
	{8'd27,8'd27} : s = 408;
	{8'd27,8'd28} : s = 484;
	{8'd27,8'd29} : s = 276;
	{8'd27,8'd30} : s = 404;
	{8'd27,8'd31} : s = 402;
	{8'd27,8'd32} : s = 482;
	{8'd27,8'd33} : s = 401;
	{8'd27,8'd34} : s = 481;
	{8'd27,8'd35} : s = 472;
	{8'd27,8'd36} : s = 504;
	{8'd27,8'd37} : s = 4;
	{8'd27,8'd38} : s = 96;
	{8'd27,8'd39} : s = 80;
	{8'd27,8'd40} : s = 274;
	{8'd27,8'd41} : s = 72;
	{8'd27,8'd42} : s = 273;
	{8'd27,8'd43} : s = 268;
	{8'd27,8'd44} : s = 396;
	{8'd27,8'd45} : s = 68;
	{8'd27,8'd46} : s = 266;
	{8'd27,8'd47} : s = 265;
	{8'd27,8'd48} : s = 394;
	{8'd27,8'd49} : s = 262;
	{8'd27,8'd50} : s = 393;
	{8'd27,8'd51} : s = 390;
	{8'd27,8'd52} : s = 468;
	{8'd27,8'd53} : s = 66;
	{8'd27,8'd54} : s = 261;
	{8'd27,8'd55} : s = 259;
	{8'd27,8'd56} : s = 389;
	{8'd27,8'd57} : s = 224;
	{8'd27,8'd58} : s = 387;
	{8'd27,8'd59} : s = 368;
	{8'd27,8'd60} : s = 466;
	{8'd27,8'd61} : s = 208;
	{8'd27,8'd62} : s = 360;
	{8'd27,8'd63} : s = 356;
	{8'd27,8'd64} : s = 465;
	{8'd27,8'd65} : s = 354;
	{8'd27,8'd66} : s = 460;
	{8'd27,8'd67} : s = 458;
	{8'd27,8'd68} : s = 500;
	{8'd27,8'd69} : s = 65;
	{8'd27,8'd70} : s = 200;
	{8'd27,8'd71} : s = 196;
	{8'd27,8'd72} : s = 353;
	{8'd27,8'd73} : s = 194;
	{8'd27,8'd74} : s = 344;
	{8'd27,8'd75} : s = 340;
	{8'd27,8'd76} : s = 457;
	{8'd27,8'd77} : s = 193;
	{8'd27,8'd78} : s = 338;
	{8'd27,8'd79} : s = 337;
	{8'd27,8'd80} : s = 454;
	{8'd27,8'd81} : s = 332;
	{8'd27,8'd82} : s = 453;
	{8'd27,8'd83} : s = 451;
	{8'd27,8'd84} : s = 498;
	{8'd27,8'd85} : s = 176;
	{8'd27,8'd86} : s = 330;
	{8'd27,8'd87} : s = 329;
	{8'd27,8'd88} : s = 440;
	{8'd27,8'd89} : s = 326;
	{8'd27,8'd90} : s = 436;
	{8'd27,8'd91} : s = 434;
	{8'd27,8'd92} : s = 497;
	{8'd27,8'd93} : s = 325;
	{8'd27,8'd94} : s = 433;
	{8'd27,8'd95} : s = 428;
	{8'd27,8'd96} : s = 492;
	{8'd27,8'd97} : s = 426;
	{8'd27,8'd98} : s = 490;
	{8'd27,8'd99} : s = 489;
	{8'd27,8'd100} : s = 508;
	{8'd27,8'd101} : s = 2;
	{8'd27,8'd102} : s = 48;
	{8'd27,8'd103} : s = 40;
	{8'd27,8'd104} : s = 168;
	{8'd27,8'd105} : s = 36;
	{8'd27,8'd106} : s = 164;
	{8'd27,8'd107} : s = 162;
	{8'd27,8'd108} : s = 323;
	{8'd27,8'd109} : s = 34;
	{8'd27,8'd110} : s = 161;
	{8'd27,8'd111} : s = 152;
	{8'd27,8'd112} : s = 312;
	{8'd27,8'd113} : s = 148;
	{8'd27,8'd114} : s = 308;
	{8'd27,8'd115} : s = 306;
	{8'd27,8'd116} : s = 425;
	{8'd27,8'd117} : s = 33;
	{8'd27,8'd118} : s = 146;
	{8'd27,8'd119} : s = 145;
	{8'd27,8'd120} : s = 305;
	{8'd27,8'd121} : s = 140;
	{8'd27,8'd122} : s = 300;
	{8'd27,8'd123} : s = 298;
	{8'd27,8'd124} : s = 422;
	{8'd27,8'd125} : s = 138;
	{8'd27,8'd126} : s = 297;
	{8'd27,8'd127} : s = 294;
	{8'd27,8'd128} : s = 421;
	{8'd27,8'd129} : s = 293;
	{8'd27,8'd130} : s = 419;
	{8'd27,8'd131} : s = 412;
	{8'd27,8'd132} : s = 486;
	{8'd27,8'd133} : s = 24;
	{8'd27,8'd134} : s = 137;
	{8'd27,8'd135} : s = 134;
	{8'd27,8'd136} : s = 291;
	{8'd27,8'd137} : s = 133;
	{8'd27,8'd138} : s = 284;
	{8'd27,8'd139} : s = 282;
	{8'd27,8'd140} : s = 410;
	{8'd27,8'd141} : s = 131;
	{8'd27,8'd142} : s = 281;
	{8'd27,8'd143} : s = 278;
	{8'd27,8'd144} : s = 409;
	{8'd27,8'd145} : s = 277;
	{8'd27,8'd146} : s = 406;
	{8'd27,8'd147} : s = 405;
	{8'd27,8'd148} : s = 485;
	{8'd27,8'd149} : s = 112;
	{8'd27,8'd150} : s = 275;
	{8'd27,8'd151} : s = 270;
	{8'd27,8'd152} : s = 403;
	{8'd27,8'd153} : s = 269;
	{8'd27,8'd154} : s = 398;
	{8'd27,8'd155} : s = 397;
	{8'd27,8'd156} : s = 483;
	{8'd27,8'd157} : s = 267;
	{8'd27,8'd158} : s = 395;
	{8'd27,8'd159} : s = 391;
	{8'd27,8'd160} : s = 476;
	{8'd27,8'd161} : s = 376;
	{8'd27,8'd162} : s = 474;
	{8'd27,8'd163} : s = 473;
	{8'd27,8'd164} : s = 506;
	{8'd27,8'd165} : s = 20;
	{8'd27,8'd166} : s = 104;
	{8'd27,8'd167} : s = 100;
	{8'd27,8'd168} : s = 263;
	{8'd27,8'd169} : s = 98;
	{8'd27,8'd170} : s = 240;
	{8'd27,8'd171} : s = 232;
	{8'd27,8'd172} : s = 372;
	{8'd27,8'd173} : s = 97;
	{8'd27,8'd174} : s = 228;
	{8'd27,8'd175} : s = 226;
	{8'd27,8'd176} : s = 370;
	{8'd27,8'd177} : s = 225;
	{8'd27,8'd178} : s = 369;
	{8'd27,8'd179} : s = 364;
	{8'd27,8'd180} : s = 470;
	{8'd27,8'd181} : s = 88;
	{8'd27,8'd182} : s = 216;
	{8'd27,8'd183} : s = 212;
	{8'd27,8'd184} : s = 362;
	{8'd27,8'd185} : s = 210;
	{8'd27,8'd186} : s = 361;
	{8'd27,8'd187} : s = 358;
	{8'd27,8'd188} : s = 469;
	{8'd27,8'd189} : s = 209;
	{8'd27,8'd190} : s = 357;
	{8'd27,8'd191} : s = 355;
	{8'd27,8'd192} : s = 467;
	{8'd27,8'd193} : s = 348;
	{8'd27,8'd194} : s = 462;
	{8'd27,8'd195} : s = 461;
	{8'd27,8'd196} : s = 505;
	{8'd27,8'd197} : s = 84;
	{8'd27,8'd198} : s = 204;
	{8'd27,8'd199} : s = 202;
	{8'd27,8'd200} : s = 346;
	{8'd27,8'd201} : s = 201;
	{8'd27,8'd202} : s = 345;
	{8'd27,8'd203} : s = 342;
	{8'd27,8'd204} : s = 459;
	{8'd27,8'd205} : s = 198;
	{8'd27,8'd206} : s = 341;
	{8'd27,8'd207} : s = 339;
	{8'd27,8'd208} : s = 455;
	{8'd27,8'd209} : s = 334;
	{8'd27,8'd210} : s = 444;
	{8'd27,8'd211} : s = 442;
	{8'd27,8'd212} : s = 502;
	{8'd27,8'd213} : s = 197;
	{8'd27,8'd214} : s = 333;
	{8'd27,8'd215} : s = 331;
	{8'd27,8'd216} : s = 441;
	{8'd27,8'd217} : s = 327;
	{8'd27,8'd218} : s = 438;
	{8'd27,8'd219} : s = 437;
	{8'd27,8'd220} : s = 501;
	{8'd27,8'd221} : s = 316;
	{8'd27,8'd222} : s = 435;
	{8'd27,8'd223} : s = 430;
	{8'd27,8'd224} : s = 499;
	{8'd27,8'd225} : s = 429;
	{8'd27,8'd226} : s = 494;
	{8'd27,8'd227} : s = 493;
	{8'd27,8'd228} : s = 510;
	{8'd27,8'd229} : s = 1;
	{8'd27,8'd230} : s = 18;
	{8'd27,8'd231} : s = 17;
	{8'd27,8'd232} : s = 82;
	{8'd27,8'd233} : s = 12;
	{8'd27,8'd234} : s = 81;
	{8'd27,8'd235} : s = 76;
	{8'd27,8'd236} : s = 195;
	{8'd27,8'd237} : s = 10;
	{8'd27,8'd238} : s = 74;
	{8'd27,8'd239} : s = 73;
	{8'd27,8'd240} : s = 184;
	{8'd27,8'd241} : s = 70;
	{8'd27,8'd242} : s = 180;
	{8'd27,8'd243} : s = 178;
	{8'd27,8'd244} : s = 314;
	{8'd27,8'd245} : s = 9;
	{8'd27,8'd246} : s = 69;
	{8'd27,8'd247} : s = 67;
	{8'd27,8'd248} : s = 177;
	{8'd27,8'd249} : s = 56;
	{8'd27,8'd250} : s = 172;
	{8'd27,8'd251} : s = 170;
	{8'd27,8'd252} : s = 313;
	{8'd27,8'd253} : s = 52;
	{8'd27,8'd254} : s = 169;
	{8'd27,8'd255} : s = 166;
	{8'd28,8'd0} : s = 328;
	{8'd28,8'd1} : s = 452;
	{8'd28,8'd2} : s = 450;
	{8'd28,8'd3} : s = 496;
	{8'd28,8'd4} : s = 16;
	{8'd28,8'd5} : s = 144;
	{8'd28,8'd6} : s = 136;
	{8'd28,8'd7} : s = 324;
	{8'd28,8'd8} : s = 132;
	{8'd28,8'd9} : s = 322;
	{8'd28,8'd10} : s = 321;
	{8'd28,8'd11} : s = 449;
	{8'd28,8'd12} : s = 130;
	{8'd28,8'd13} : s = 304;
	{8'd28,8'd14} : s = 296;
	{8'd28,8'd15} : s = 432;
	{8'd28,8'd16} : s = 292;
	{8'd28,8'd17} : s = 424;
	{8'd28,8'd18} : s = 420;
	{8'd28,8'd19} : s = 488;
	{8'd28,8'd20} : s = 129;
	{8'd28,8'd21} : s = 290;
	{8'd28,8'd22} : s = 289;
	{8'd28,8'd23} : s = 418;
	{8'd28,8'd24} : s = 280;
	{8'd28,8'd25} : s = 417;
	{8'd28,8'd26} : s = 408;
	{8'd28,8'd27} : s = 484;
	{8'd28,8'd28} : s = 276;
	{8'd28,8'd29} : s = 404;
	{8'd28,8'd30} : s = 402;
	{8'd28,8'd31} : s = 482;
	{8'd28,8'd32} : s = 401;
	{8'd28,8'd33} : s = 481;
	{8'd28,8'd34} : s = 472;
	{8'd28,8'd35} : s = 504;
	{8'd28,8'd36} : s = 4;
	{8'd28,8'd37} : s = 96;
	{8'd28,8'd38} : s = 80;
	{8'd28,8'd39} : s = 274;
	{8'd28,8'd40} : s = 72;
	{8'd28,8'd41} : s = 273;
	{8'd28,8'd42} : s = 268;
	{8'd28,8'd43} : s = 396;
	{8'd28,8'd44} : s = 68;
	{8'd28,8'd45} : s = 266;
	{8'd28,8'd46} : s = 265;
	{8'd28,8'd47} : s = 394;
	{8'd28,8'd48} : s = 262;
	{8'd28,8'd49} : s = 393;
	{8'd28,8'd50} : s = 390;
	{8'd28,8'd51} : s = 468;
	{8'd28,8'd52} : s = 66;
	{8'd28,8'd53} : s = 261;
	{8'd28,8'd54} : s = 259;
	{8'd28,8'd55} : s = 389;
	{8'd28,8'd56} : s = 224;
	{8'd28,8'd57} : s = 387;
	{8'd28,8'd58} : s = 368;
	{8'd28,8'd59} : s = 466;
	{8'd28,8'd60} : s = 208;
	{8'd28,8'd61} : s = 360;
	{8'd28,8'd62} : s = 356;
	{8'd28,8'd63} : s = 465;
	{8'd28,8'd64} : s = 354;
	{8'd28,8'd65} : s = 460;
	{8'd28,8'd66} : s = 458;
	{8'd28,8'd67} : s = 500;
	{8'd28,8'd68} : s = 65;
	{8'd28,8'd69} : s = 200;
	{8'd28,8'd70} : s = 196;
	{8'd28,8'd71} : s = 353;
	{8'd28,8'd72} : s = 194;
	{8'd28,8'd73} : s = 344;
	{8'd28,8'd74} : s = 340;
	{8'd28,8'd75} : s = 457;
	{8'd28,8'd76} : s = 193;
	{8'd28,8'd77} : s = 338;
	{8'd28,8'd78} : s = 337;
	{8'd28,8'd79} : s = 454;
	{8'd28,8'd80} : s = 332;
	{8'd28,8'd81} : s = 453;
	{8'd28,8'd82} : s = 451;
	{8'd28,8'd83} : s = 498;
	{8'd28,8'd84} : s = 176;
	{8'd28,8'd85} : s = 330;
	{8'd28,8'd86} : s = 329;
	{8'd28,8'd87} : s = 440;
	{8'd28,8'd88} : s = 326;
	{8'd28,8'd89} : s = 436;
	{8'd28,8'd90} : s = 434;
	{8'd28,8'd91} : s = 497;
	{8'd28,8'd92} : s = 325;
	{8'd28,8'd93} : s = 433;
	{8'd28,8'd94} : s = 428;
	{8'd28,8'd95} : s = 492;
	{8'd28,8'd96} : s = 426;
	{8'd28,8'd97} : s = 490;
	{8'd28,8'd98} : s = 489;
	{8'd28,8'd99} : s = 508;
	{8'd28,8'd100} : s = 2;
	{8'd28,8'd101} : s = 48;
	{8'd28,8'd102} : s = 40;
	{8'd28,8'd103} : s = 168;
	{8'd28,8'd104} : s = 36;
	{8'd28,8'd105} : s = 164;
	{8'd28,8'd106} : s = 162;
	{8'd28,8'd107} : s = 323;
	{8'd28,8'd108} : s = 34;
	{8'd28,8'd109} : s = 161;
	{8'd28,8'd110} : s = 152;
	{8'd28,8'd111} : s = 312;
	{8'd28,8'd112} : s = 148;
	{8'd28,8'd113} : s = 308;
	{8'd28,8'd114} : s = 306;
	{8'd28,8'd115} : s = 425;
	{8'd28,8'd116} : s = 33;
	{8'd28,8'd117} : s = 146;
	{8'd28,8'd118} : s = 145;
	{8'd28,8'd119} : s = 305;
	{8'd28,8'd120} : s = 140;
	{8'd28,8'd121} : s = 300;
	{8'd28,8'd122} : s = 298;
	{8'd28,8'd123} : s = 422;
	{8'd28,8'd124} : s = 138;
	{8'd28,8'd125} : s = 297;
	{8'd28,8'd126} : s = 294;
	{8'd28,8'd127} : s = 421;
	{8'd28,8'd128} : s = 293;
	{8'd28,8'd129} : s = 419;
	{8'd28,8'd130} : s = 412;
	{8'd28,8'd131} : s = 486;
	{8'd28,8'd132} : s = 24;
	{8'd28,8'd133} : s = 137;
	{8'd28,8'd134} : s = 134;
	{8'd28,8'd135} : s = 291;
	{8'd28,8'd136} : s = 133;
	{8'd28,8'd137} : s = 284;
	{8'd28,8'd138} : s = 282;
	{8'd28,8'd139} : s = 410;
	{8'd28,8'd140} : s = 131;
	{8'd28,8'd141} : s = 281;
	{8'd28,8'd142} : s = 278;
	{8'd28,8'd143} : s = 409;
	{8'd28,8'd144} : s = 277;
	{8'd28,8'd145} : s = 406;
	{8'd28,8'd146} : s = 405;
	{8'd28,8'd147} : s = 485;
	{8'd28,8'd148} : s = 112;
	{8'd28,8'd149} : s = 275;
	{8'd28,8'd150} : s = 270;
	{8'd28,8'd151} : s = 403;
	{8'd28,8'd152} : s = 269;
	{8'd28,8'd153} : s = 398;
	{8'd28,8'd154} : s = 397;
	{8'd28,8'd155} : s = 483;
	{8'd28,8'd156} : s = 267;
	{8'd28,8'd157} : s = 395;
	{8'd28,8'd158} : s = 391;
	{8'd28,8'd159} : s = 476;
	{8'd28,8'd160} : s = 376;
	{8'd28,8'd161} : s = 474;
	{8'd28,8'd162} : s = 473;
	{8'd28,8'd163} : s = 506;
	{8'd28,8'd164} : s = 20;
	{8'd28,8'd165} : s = 104;
	{8'd28,8'd166} : s = 100;
	{8'd28,8'd167} : s = 263;
	{8'd28,8'd168} : s = 98;
	{8'd28,8'd169} : s = 240;
	{8'd28,8'd170} : s = 232;
	{8'd28,8'd171} : s = 372;
	{8'd28,8'd172} : s = 97;
	{8'd28,8'd173} : s = 228;
	{8'd28,8'd174} : s = 226;
	{8'd28,8'd175} : s = 370;
	{8'd28,8'd176} : s = 225;
	{8'd28,8'd177} : s = 369;
	{8'd28,8'd178} : s = 364;
	{8'd28,8'd179} : s = 470;
	{8'd28,8'd180} : s = 88;
	{8'd28,8'd181} : s = 216;
	{8'd28,8'd182} : s = 212;
	{8'd28,8'd183} : s = 362;
	{8'd28,8'd184} : s = 210;
	{8'd28,8'd185} : s = 361;
	{8'd28,8'd186} : s = 358;
	{8'd28,8'd187} : s = 469;
	{8'd28,8'd188} : s = 209;
	{8'd28,8'd189} : s = 357;
	{8'd28,8'd190} : s = 355;
	{8'd28,8'd191} : s = 467;
	{8'd28,8'd192} : s = 348;
	{8'd28,8'd193} : s = 462;
	{8'd28,8'd194} : s = 461;
	{8'd28,8'd195} : s = 505;
	{8'd28,8'd196} : s = 84;
	{8'd28,8'd197} : s = 204;
	{8'd28,8'd198} : s = 202;
	{8'd28,8'd199} : s = 346;
	{8'd28,8'd200} : s = 201;
	{8'd28,8'd201} : s = 345;
	{8'd28,8'd202} : s = 342;
	{8'd28,8'd203} : s = 459;
	{8'd28,8'd204} : s = 198;
	{8'd28,8'd205} : s = 341;
	{8'd28,8'd206} : s = 339;
	{8'd28,8'd207} : s = 455;
	{8'd28,8'd208} : s = 334;
	{8'd28,8'd209} : s = 444;
	{8'd28,8'd210} : s = 442;
	{8'd28,8'd211} : s = 502;
	{8'd28,8'd212} : s = 197;
	{8'd28,8'd213} : s = 333;
	{8'd28,8'd214} : s = 331;
	{8'd28,8'd215} : s = 441;
	{8'd28,8'd216} : s = 327;
	{8'd28,8'd217} : s = 438;
	{8'd28,8'd218} : s = 437;
	{8'd28,8'd219} : s = 501;
	{8'd28,8'd220} : s = 316;
	{8'd28,8'd221} : s = 435;
	{8'd28,8'd222} : s = 430;
	{8'd28,8'd223} : s = 499;
	{8'd28,8'd224} : s = 429;
	{8'd28,8'd225} : s = 494;
	{8'd28,8'd226} : s = 493;
	{8'd28,8'd227} : s = 510;
	{8'd28,8'd228} : s = 1;
	{8'd28,8'd229} : s = 18;
	{8'd28,8'd230} : s = 17;
	{8'd28,8'd231} : s = 82;
	{8'd28,8'd232} : s = 12;
	{8'd28,8'd233} : s = 81;
	{8'd28,8'd234} : s = 76;
	{8'd28,8'd235} : s = 195;
	{8'd28,8'd236} : s = 10;
	{8'd28,8'd237} : s = 74;
	{8'd28,8'd238} : s = 73;
	{8'd28,8'd239} : s = 184;
	{8'd28,8'd240} : s = 70;
	{8'd28,8'd241} : s = 180;
	{8'd28,8'd242} : s = 178;
	{8'd28,8'd243} : s = 314;
	{8'd28,8'd244} : s = 9;
	{8'd28,8'd245} : s = 69;
	{8'd28,8'd246} : s = 67;
	{8'd28,8'd247} : s = 177;
	{8'd28,8'd248} : s = 56;
	{8'd28,8'd249} : s = 172;
	{8'd28,8'd250} : s = 170;
	{8'd28,8'd251} : s = 313;
	{8'd28,8'd252} : s = 52;
	{8'd28,8'd253} : s = 169;
	{8'd28,8'd254} : s = 166;
	{8'd28,8'd255} : s = 310;
	{8'd29,8'd0} : s = 452;
	{8'd29,8'd1} : s = 450;
	{8'd29,8'd2} : s = 496;
	{8'd29,8'd3} : s = 16;
	{8'd29,8'd4} : s = 144;
	{8'd29,8'd5} : s = 136;
	{8'd29,8'd6} : s = 324;
	{8'd29,8'd7} : s = 132;
	{8'd29,8'd8} : s = 322;
	{8'd29,8'd9} : s = 321;
	{8'd29,8'd10} : s = 449;
	{8'd29,8'd11} : s = 130;
	{8'd29,8'd12} : s = 304;
	{8'd29,8'd13} : s = 296;
	{8'd29,8'd14} : s = 432;
	{8'd29,8'd15} : s = 292;
	{8'd29,8'd16} : s = 424;
	{8'd29,8'd17} : s = 420;
	{8'd29,8'd18} : s = 488;
	{8'd29,8'd19} : s = 129;
	{8'd29,8'd20} : s = 290;
	{8'd29,8'd21} : s = 289;
	{8'd29,8'd22} : s = 418;
	{8'd29,8'd23} : s = 280;
	{8'd29,8'd24} : s = 417;
	{8'd29,8'd25} : s = 408;
	{8'd29,8'd26} : s = 484;
	{8'd29,8'd27} : s = 276;
	{8'd29,8'd28} : s = 404;
	{8'd29,8'd29} : s = 402;
	{8'd29,8'd30} : s = 482;
	{8'd29,8'd31} : s = 401;
	{8'd29,8'd32} : s = 481;
	{8'd29,8'd33} : s = 472;
	{8'd29,8'd34} : s = 504;
	{8'd29,8'd35} : s = 4;
	{8'd29,8'd36} : s = 96;
	{8'd29,8'd37} : s = 80;
	{8'd29,8'd38} : s = 274;
	{8'd29,8'd39} : s = 72;
	{8'd29,8'd40} : s = 273;
	{8'd29,8'd41} : s = 268;
	{8'd29,8'd42} : s = 396;
	{8'd29,8'd43} : s = 68;
	{8'd29,8'd44} : s = 266;
	{8'd29,8'd45} : s = 265;
	{8'd29,8'd46} : s = 394;
	{8'd29,8'd47} : s = 262;
	{8'd29,8'd48} : s = 393;
	{8'd29,8'd49} : s = 390;
	{8'd29,8'd50} : s = 468;
	{8'd29,8'd51} : s = 66;
	{8'd29,8'd52} : s = 261;
	{8'd29,8'd53} : s = 259;
	{8'd29,8'd54} : s = 389;
	{8'd29,8'd55} : s = 224;
	{8'd29,8'd56} : s = 387;
	{8'd29,8'd57} : s = 368;
	{8'd29,8'd58} : s = 466;
	{8'd29,8'd59} : s = 208;
	{8'd29,8'd60} : s = 360;
	{8'd29,8'd61} : s = 356;
	{8'd29,8'd62} : s = 465;
	{8'd29,8'd63} : s = 354;
	{8'd29,8'd64} : s = 460;
	{8'd29,8'd65} : s = 458;
	{8'd29,8'd66} : s = 500;
	{8'd29,8'd67} : s = 65;
	{8'd29,8'd68} : s = 200;
	{8'd29,8'd69} : s = 196;
	{8'd29,8'd70} : s = 353;
	{8'd29,8'd71} : s = 194;
	{8'd29,8'd72} : s = 344;
	{8'd29,8'd73} : s = 340;
	{8'd29,8'd74} : s = 457;
	{8'd29,8'd75} : s = 193;
	{8'd29,8'd76} : s = 338;
	{8'd29,8'd77} : s = 337;
	{8'd29,8'd78} : s = 454;
	{8'd29,8'd79} : s = 332;
	{8'd29,8'd80} : s = 453;
	{8'd29,8'd81} : s = 451;
	{8'd29,8'd82} : s = 498;
	{8'd29,8'd83} : s = 176;
	{8'd29,8'd84} : s = 330;
	{8'd29,8'd85} : s = 329;
	{8'd29,8'd86} : s = 440;
	{8'd29,8'd87} : s = 326;
	{8'd29,8'd88} : s = 436;
	{8'd29,8'd89} : s = 434;
	{8'd29,8'd90} : s = 497;
	{8'd29,8'd91} : s = 325;
	{8'd29,8'd92} : s = 433;
	{8'd29,8'd93} : s = 428;
	{8'd29,8'd94} : s = 492;
	{8'd29,8'd95} : s = 426;
	{8'd29,8'd96} : s = 490;
	{8'd29,8'd97} : s = 489;
	{8'd29,8'd98} : s = 508;
	{8'd29,8'd99} : s = 2;
	{8'd29,8'd100} : s = 48;
	{8'd29,8'd101} : s = 40;
	{8'd29,8'd102} : s = 168;
	{8'd29,8'd103} : s = 36;
	{8'd29,8'd104} : s = 164;
	{8'd29,8'd105} : s = 162;
	{8'd29,8'd106} : s = 323;
	{8'd29,8'd107} : s = 34;
	{8'd29,8'd108} : s = 161;
	{8'd29,8'd109} : s = 152;
	{8'd29,8'd110} : s = 312;
	{8'd29,8'd111} : s = 148;
	{8'd29,8'd112} : s = 308;
	{8'd29,8'd113} : s = 306;
	{8'd29,8'd114} : s = 425;
	{8'd29,8'd115} : s = 33;
	{8'd29,8'd116} : s = 146;
	{8'd29,8'd117} : s = 145;
	{8'd29,8'd118} : s = 305;
	{8'd29,8'd119} : s = 140;
	{8'd29,8'd120} : s = 300;
	{8'd29,8'd121} : s = 298;
	{8'd29,8'd122} : s = 422;
	{8'd29,8'd123} : s = 138;
	{8'd29,8'd124} : s = 297;
	{8'd29,8'd125} : s = 294;
	{8'd29,8'd126} : s = 421;
	{8'd29,8'd127} : s = 293;
	{8'd29,8'd128} : s = 419;
	{8'd29,8'd129} : s = 412;
	{8'd29,8'd130} : s = 486;
	{8'd29,8'd131} : s = 24;
	{8'd29,8'd132} : s = 137;
	{8'd29,8'd133} : s = 134;
	{8'd29,8'd134} : s = 291;
	{8'd29,8'd135} : s = 133;
	{8'd29,8'd136} : s = 284;
	{8'd29,8'd137} : s = 282;
	{8'd29,8'd138} : s = 410;
	{8'd29,8'd139} : s = 131;
	{8'd29,8'd140} : s = 281;
	{8'd29,8'd141} : s = 278;
	{8'd29,8'd142} : s = 409;
	{8'd29,8'd143} : s = 277;
	{8'd29,8'd144} : s = 406;
	{8'd29,8'd145} : s = 405;
	{8'd29,8'd146} : s = 485;
	{8'd29,8'd147} : s = 112;
	{8'd29,8'd148} : s = 275;
	{8'd29,8'd149} : s = 270;
	{8'd29,8'd150} : s = 403;
	{8'd29,8'd151} : s = 269;
	{8'd29,8'd152} : s = 398;
	{8'd29,8'd153} : s = 397;
	{8'd29,8'd154} : s = 483;
	{8'd29,8'd155} : s = 267;
	{8'd29,8'd156} : s = 395;
	{8'd29,8'd157} : s = 391;
	{8'd29,8'd158} : s = 476;
	{8'd29,8'd159} : s = 376;
	{8'd29,8'd160} : s = 474;
	{8'd29,8'd161} : s = 473;
	{8'd29,8'd162} : s = 506;
	{8'd29,8'd163} : s = 20;
	{8'd29,8'd164} : s = 104;
	{8'd29,8'd165} : s = 100;
	{8'd29,8'd166} : s = 263;
	{8'd29,8'd167} : s = 98;
	{8'd29,8'd168} : s = 240;
	{8'd29,8'd169} : s = 232;
	{8'd29,8'd170} : s = 372;
	{8'd29,8'd171} : s = 97;
	{8'd29,8'd172} : s = 228;
	{8'd29,8'd173} : s = 226;
	{8'd29,8'd174} : s = 370;
	{8'd29,8'd175} : s = 225;
	{8'd29,8'd176} : s = 369;
	{8'd29,8'd177} : s = 364;
	{8'd29,8'd178} : s = 470;
	{8'd29,8'd179} : s = 88;
	{8'd29,8'd180} : s = 216;
	{8'd29,8'd181} : s = 212;
	{8'd29,8'd182} : s = 362;
	{8'd29,8'd183} : s = 210;
	{8'd29,8'd184} : s = 361;
	{8'd29,8'd185} : s = 358;
	{8'd29,8'd186} : s = 469;
	{8'd29,8'd187} : s = 209;
	{8'd29,8'd188} : s = 357;
	{8'd29,8'd189} : s = 355;
	{8'd29,8'd190} : s = 467;
	{8'd29,8'd191} : s = 348;
	{8'd29,8'd192} : s = 462;
	{8'd29,8'd193} : s = 461;
	{8'd29,8'd194} : s = 505;
	{8'd29,8'd195} : s = 84;
	{8'd29,8'd196} : s = 204;
	{8'd29,8'd197} : s = 202;
	{8'd29,8'd198} : s = 346;
	{8'd29,8'd199} : s = 201;
	{8'd29,8'd200} : s = 345;
	{8'd29,8'd201} : s = 342;
	{8'd29,8'd202} : s = 459;
	{8'd29,8'd203} : s = 198;
	{8'd29,8'd204} : s = 341;
	{8'd29,8'd205} : s = 339;
	{8'd29,8'd206} : s = 455;
	{8'd29,8'd207} : s = 334;
	{8'd29,8'd208} : s = 444;
	{8'd29,8'd209} : s = 442;
	{8'd29,8'd210} : s = 502;
	{8'd29,8'd211} : s = 197;
	{8'd29,8'd212} : s = 333;
	{8'd29,8'd213} : s = 331;
	{8'd29,8'd214} : s = 441;
	{8'd29,8'd215} : s = 327;
	{8'd29,8'd216} : s = 438;
	{8'd29,8'd217} : s = 437;
	{8'd29,8'd218} : s = 501;
	{8'd29,8'd219} : s = 316;
	{8'd29,8'd220} : s = 435;
	{8'd29,8'd221} : s = 430;
	{8'd29,8'd222} : s = 499;
	{8'd29,8'd223} : s = 429;
	{8'd29,8'd224} : s = 494;
	{8'd29,8'd225} : s = 493;
	{8'd29,8'd226} : s = 510;
	{8'd29,8'd227} : s = 1;
	{8'd29,8'd228} : s = 18;
	{8'd29,8'd229} : s = 17;
	{8'd29,8'd230} : s = 82;
	{8'd29,8'd231} : s = 12;
	{8'd29,8'd232} : s = 81;
	{8'd29,8'd233} : s = 76;
	{8'd29,8'd234} : s = 195;
	{8'd29,8'd235} : s = 10;
	{8'd29,8'd236} : s = 74;
	{8'd29,8'd237} : s = 73;
	{8'd29,8'd238} : s = 184;
	{8'd29,8'd239} : s = 70;
	{8'd29,8'd240} : s = 180;
	{8'd29,8'd241} : s = 178;
	{8'd29,8'd242} : s = 314;
	{8'd29,8'd243} : s = 9;
	{8'd29,8'd244} : s = 69;
	{8'd29,8'd245} : s = 67;
	{8'd29,8'd246} : s = 177;
	{8'd29,8'd247} : s = 56;
	{8'd29,8'd248} : s = 172;
	{8'd29,8'd249} : s = 170;
	{8'd29,8'd250} : s = 313;
	{8'd29,8'd251} : s = 52;
	{8'd29,8'd252} : s = 169;
	{8'd29,8'd253} : s = 166;
	{8'd29,8'd254} : s = 310;
	{8'd29,8'd255} : s = 165;
	{8'd30,8'd0} : s = 450;
	{8'd30,8'd1} : s = 496;
	{8'd30,8'd2} : s = 16;
	{8'd30,8'd3} : s = 144;
	{8'd30,8'd4} : s = 136;
	{8'd30,8'd5} : s = 324;
	{8'd30,8'd6} : s = 132;
	{8'd30,8'd7} : s = 322;
	{8'd30,8'd8} : s = 321;
	{8'd30,8'd9} : s = 449;
	{8'd30,8'd10} : s = 130;
	{8'd30,8'd11} : s = 304;
	{8'd30,8'd12} : s = 296;
	{8'd30,8'd13} : s = 432;
	{8'd30,8'd14} : s = 292;
	{8'd30,8'd15} : s = 424;
	{8'd30,8'd16} : s = 420;
	{8'd30,8'd17} : s = 488;
	{8'd30,8'd18} : s = 129;
	{8'd30,8'd19} : s = 290;
	{8'd30,8'd20} : s = 289;
	{8'd30,8'd21} : s = 418;
	{8'd30,8'd22} : s = 280;
	{8'd30,8'd23} : s = 417;
	{8'd30,8'd24} : s = 408;
	{8'd30,8'd25} : s = 484;
	{8'd30,8'd26} : s = 276;
	{8'd30,8'd27} : s = 404;
	{8'd30,8'd28} : s = 402;
	{8'd30,8'd29} : s = 482;
	{8'd30,8'd30} : s = 401;
	{8'd30,8'd31} : s = 481;
	{8'd30,8'd32} : s = 472;
	{8'd30,8'd33} : s = 504;
	{8'd30,8'd34} : s = 4;
	{8'd30,8'd35} : s = 96;
	{8'd30,8'd36} : s = 80;
	{8'd30,8'd37} : s = 274;
	{8'd30,8'd38} : s = 72;
	{8'd30,8'd39} : s = 273;
	{8'd30,8'd40} : s = 268;
	{8'd30,8'd41} : s = 396;
	{8'd30,8'd42} : s = 68;
	{8'd30,8'd43} : s = 266;
	{8'd30,8'd44} : s = 265;
	{8'd30,8'd45} : s = 394;
	{8'd30,8'd46} : s = 262;
	{8'd30,8'd47} : s = 393;
	{8'd30,8'd48} : s = 390;
	{8'd30,8'd49} : s = 468;
	{8'd30,8'd50} : s = 66;
	{8'd30,8'd51} : s = 261;
	{8'd30,8'd52} : s = 259;
	{8'd30,8'd53} : s = 389;
	{8'd30,8'd54} : s = 224;
	{8'd30,8'd55} : s = 387;
	{8'd30,8'd56} : s = 368;
	{8'd30,8'd57} : s = 466;
	{8'd30,8'd58} : s = 208;
	{8'd30,8'd59} : s = 360;
	{8'd30,8'd60} : s = 356;
	{8'd30,8'd61} : s = 465;
	{8'd30,8'd62} : s = 354;
	{8'd30,8'd63} : s = 460;
	{8'd30,8'd64} : s = 458;
	{8'd30,8'd65} : s = 500;
	{8'd30,8'd66} : s = 65;
	{8'd30,8'd67} : s = 200;
	{8'd30,8'd68} : s = 196;
	{8'd30,8'd69} : s = 353;
	{8'd30,8'd70} : s = 194;
	{8'd30,8'd71} : s = 344;
	{8'd30,8'd72} : s = 340;
	{8'd30,8'd73} : s = 457;
	{8'd30,8'd74} : s = 193;
	{8'd30,8'd75} : s = 338;
	{8'd30,8'd76} : s = 337;
	{8'd30,8'd77} : s = 454;
	{8'd30,8'd78} : s = 332;
	{8'd30,8'd79} : s = 453;
	{8'd30,8'd80} : s = 451;
	{8'd30,8'd81} : s = 498;
	{8'd30,8'd82} : s = 176;
	{8'd30,8'd83} : s = 330;
	{8'd30,8'd84} : s = 329;
	{8'd30,8'd85} : s = 440;
	{8'd30,8'd86} : s = 326;
	{8'd30,8'd87} : s = 436;
	{8'd30,8'd88} : s = 434;
	{8'd30,8'd89} : s = 497;
	{8'd30,8'd90} : s = 325;
	{8'd30,8'd91} : s = 433;
	{8'd30,8'd92} : s = 428;
	{8'd30,8'd93} : s = 492;
	{8'd30,8'd94} : s = 426;
	{8'd30,8'd95} : s = 490;
	{8'd30,8'd96} : s = 489;
	{8'd30,8'd97} : s = 508;
	{8'd30,8'd98} : s = 2;
	{8'd30,8'd99} : s = 48;
	{8'd30,8'd100} : s = 40;
	{8'd30,8'd101} : s = 168;
	{8'd30,8'd102} : s = 36;
	{8'd30,8'd103} : s = 164;
	{8'd30,8'd104} : s = 162;
	{8'd30,8'd105} : s = 323;
	{8'd30,8'd106} : s = 34;
	{8'd30,8'd107} : s = 161;
	{8'd30,8'd108} : s = 152;
	{8'd30,8'd109} : s = 312;
	{8'd30,8'd110} : s = 148;
	{8'd30,8'd111} : s = 308;
	{8'd30,8'd112} : s = 306;
	{8'd30,8'd113} : s = 425;
	{8'd30,8'd114} : s = 33;
	{8'd30,8'd115} : s = 146;
	{8'd30,8'd116} : s = 145;
	{8'd30,8'd117} : s = 305;
	{8'd30,8'd118} : s = 140;
	{8'd30,8'd119} : s = 300;
	{8'd30,8'd120} : s = 298;
	{8'd30,8'd121} : s = 422;
	{8'd30,8'd122} : s = 138;
	{8'd30,8'd123} : s = 297;
	{8'd30,8'd124} : s = 294;
	{8'd30,8'd125} : s = 421;
	{8'd30,8'd126} : s = 293;
	{8'd30,8'd127} : s = 419;
	{8'd30,8'd128} : s = 412;
	{8'd30,8'd129} : s = 486;
	{8'd30,8'd130} : s = 24;
	{8'd30,8'd131} : s = 137;
	{8'd30,8'd132} : s = 134;
	{8'd30,8'd133} : s = 291;
	{8'd30,8'd134} : s = 133;
	{8'd30,8'd135} : s = 284;
	{8'd30,8'd136} : s = 282;
	{8'd30,8'd137} : s = 410;
	{8'd30,8'd138} : s = 131;
	{8'd30,8'd139} : s = 281;
	{8'd30,8'd140} : s = 278;
	{8'd30,8'd141} : s = 409;
	{8'd30,8'd142} : s = 277;
	{8'd30,8'd143} : s = 406;
	{8'd30,8'd144} : s = 405;
	{8'd30,8'd145} : s = 485;
	{8'd30,8'd146} : s = 112;
	{8'd30,8'd147} : s = 275;
	{8'd30,8'd148} : s = 270;
	{8'd30,8'd149} : s = 403;
	{8'd30,8'd150} : s = 269;
	{8'd30,8'd151} : s = 398;
	{8'd30,8'd152} : s = 397;
	{8'd30,8'd153} : s = 483;
	{8'd30,8'd154} : s = 267;
	{8'd30,8'd155} : s = 395;
	{8'd30,8'd156} : s = 391;
	{8'd30,8'd157} : s = 476;
	{8'd30,8'd158} : s = 376;
	{8'd30,8'd159} : s = 474;
	{8'd30,8'd160} : s = 473;
	{8'd30,8'd161} : s = 506;
	{8'd30,8'd162} : s = 20;
	{8'd30,8'd163} : s = 104;
	{8'd30,8'd164} : s = 100;
	{8'd30,8'd165} : s = 263;
	{8'd30,8'd166} : s = 98;
	{8'd30,8'd167} : s = 240;
	{8'd30,8'd168} : s = 232;
	{8'd30,8'd169} : s = 372;
	{8'd30,8'd170} : s = 97;
	{8'd30,8'd171} : s = 228;
	{8'd30,8'd172} : s = 226;
	{8'd30,8'd173} : s = 370;
	{8'd30,8'd174} : s = 225;
	{8'd30,8'd175} : s = 369;
	{8'd30,8'd176} : s = 364;
	{8'd30,8'd177} : s = 470;
	{8'd30,8'd178} : s = 88;
	{8'd30,8'd179} : s = 216;
	{8'd30,8'd180} : s = 212;
	{8'd30,8'd181} : s = 362;
	{8'd30,8'd182} : s = 210;
	{8'd30,8'd183} : s = 361;
	{8'd30,8'd184} : s = 358;
	{8'd30,8'd185} : s = 469;
	{8'd30,8'd186} : s = 209;
	{8'd30,8'd187} : s = 357;
	{8'd30,8'd188} : s = 355;
	{8'd30,8'd189} : s = 467;
	{8'd30,8'd190} : s = 348;
	{8'd30,8'd191} : s = 462;
	{8'd30,8'd192} : s = 461;
	{8'd30,8'd193} : s = 505;
	{8'd30,8'd194} : s = 84;
	{8'd30,8'd195} : s = 204;
	{8'd30,8'd196} : s = 202;
	{8'd30,8'd197} : s = 346;
	{8'd30,8'd198} : s = 201;
	{8'd30,8'd199} : s = 345;
	{8'd30,8'd200} : s = 342;
	{8'd30,8'd201} : s = 459;
	{8'd30,8'd202} : s = 198;
	{8'd30,8'd203} : s = 341;
	{8'd30,8'd204} : s = 339;
	{8'd30,8'd205} : s = 455;
	{8'd30,8'd206} : s = 334;
	{8'd30,8'd207} : s = 444;
	{8'd30,8'd208} : s = 442;
	{8'd30,8'd209} : s = 502;
	{8'd30,8'd210} : s = 197;
	{8'd30,8'd211} : s = 333;
	{8'd30,8'd212} : s = 331;
	{8'd30,8'd213} : s = 441;
	{8'd30,8'd214} : s = 327;
	{8'd30,8'd215} : s = 438;
	{8'd30,8'd216} : s = 437;
	{8'd30,8'd217} : s = 501;
	{8'd30,8'd218} : s = 316;
	{8'd30,8'd219} : s = 435;
	{8'd30,8'd220} : s = 430;
	{8'd30,8'd221} : s = 499;
	{8'd30,8'd222} : s = 429;
	{8'd30,8'd223} : s = 494;
	{8'd30,8'd224} : s = 493;
	{8'd30,8'd225} : s = 510;
	{8'd30,8'd226} : s = 1;
	{8'd30,8'd227} : s = 18;
	{8'd30,8'd228} : s = 17;
	{8'd30,8'd229} : s = 82;
	{8'd30,8'd230} : s = 12;
	{8'd30,8'd231} : s = 81;
	{8'd30,8'd232} : s = 76;
	{8'd30,8'd233} : s = 195;
	{8'd30,8'd234} : s = 10;
	{8'd30,8'd235} : s = 74;
	{8'd30,8'd236} : s = 73;
	{8'd30,8'd237} : s = 184;
	{8'd30,8'd238} : s = 70;
	{8'd30,8'd239} : s = 180;
	{8'd30,8'd240} : s = 178;
	{8'd30,8'd241} : s = 314;
	{8'd30,8'd242} : s = 9;
	{8'd30,8'd243} : s = 69;
	{8'd30,8'd244} : s = 67;
	{8'd30,8'd245} : s = 177;
	{8'd30,8'd246} : s = 56;
	{8'd30,8'd247} : s = 172;
	{8'd30,8'd248} : s = 170;
	{8'd30,8'd249} : s = 313;
	{8'd30,8'd250} : s = 52;
	{8'd30,8'd251} : s = 169;
	{8'd30,8'd252} : s = 166;
	{8'd30,8'd253} : s = 310;
	{8'd30,8'd254} : s = 165;
	{8'd30,8'd255} : s = 309;
	{8'd31,8'd0} : s = 496;
	{8'd31,8'd1} : s = 16;
	{8'd31,8'd2} : s = 144;
	{8'd31,8'd3} : s = 136;
	{8'd31,8'd4} : s = 324;
	{8'd31,8'd5} : s = 132;
	{8'd31,8'd6} : s = 322;
	{8'd31,8'd7} : s = 321;
	{8'd31,8'd8} : s = 449;
	{8'd31,8'd9} : s = 130;
	{8'd31,8'd10} : s = 304;
	{8'd31,8'd11} : s = 296;
	{8'd31,8'd12} : s = 432;
	{8'd31,8'd13} : s = 292;
	{8'd31,8'd14} : s = 424;
	{8'd31,8'd15} : s = 420;
	{8'd31,8'd16} : s = 488;
	{8'd31,8'd17} : s = 129;
	{8'd31,8'd18} : s = 290;
	{8'd31,8'd19} : s = 289;
	{8'd31,8'd20} : s = 418;
	{8'd31,8'd21} : s = 280;
	{8'd31,8'd22} : s = 417;
	{8'd31,8'd23} : s = 408;
	{8'd31,8'd24} : s = 484;
	{8'd31,8'd25} : s = 276;
	{8'd31,8'd26} : s = 404;
	{8'd31,8'd27} : s = 402;
	{8'd31,8'd28} : s = 482;
	{8'd31,8'd29} : s = 401;
	{8'd31,8'd30} : s = 481;
	{8'd31,8'd31} : s = 472;
	{8'd31,8'd32} : s = 504;
	{8'd31,8'd33} : s = 4;
	{8'd31,8'd34} : s = 96;
	{8'd31,8'd35} : s = 80;
	{8'd31,8'd36} : s = 274;
	{8'd31,8'd37} : s = 72;
	{8'd31,8'd38} : s = 273;
	{8'd31,8'd39} : s = 268;
	{8'd31,8'd40} : s = 396;
	{8'd31,8'd41} : s = 68;
	{8'd31,8'd42} : s = 266;
	{8'd31,8'd43} : s = 265;
	{8'd31,8'd44} : s = 394;
	{8'd31,8'd45} : s = 262;
	{8'd31,8'd46} : s = 393;
	{8'd31,8'd47} : s = 390;
	{8'd31,8'd48} : s = 468;
	{8'd31,8'd49} : s = 66;
	{8'd31,8'd50} : s = 261;
	{8'd31,8'd51} : s = 259;
	{8'd31,8'd52} : s = 389;
	{8'd31,8'd53} : s = 224;
	{8'd31,8'd54} : s = 387;
	{8'd31,8'd55} : s = 368;
	{8'd31,8'd56} : s = 466;
	{8'd31,8'd57} : s = 208;
	{8'd31,8'd58} : s = 360;
	{8'd31,8'd59} : s = 356;
	{8'd31,8'd60} : s = 465;
	{8'd31,8'd61} : s = 354;
	{8'd31,8'd62} : s = 460;
	{8'd31,8'd63} : s = 458;
	{8'd31,8'd64} : s = 500;
	{8'd31,8'd65} : s = 65;
	{8'd31,8'd66} : s = 200;
	{8'd31,8'd67} : s = 196;
	{8'd31,8'd68} : s = 353;
	{8'd31,8'd69} : s = 194;
	{8'd31,8'd70} : s = 344;
	{8'd31,8'd71} : s = 340;
	{8'd31,8'd72} : s = 457;
	{8'd31,8'd73} : s = 193;
	{8'd31,8'd74} : s = 338;
	{8'd31,8'd75} : s = 337;
	{8'd31,8'd76} : s = 454;
	{8'd31,8'd77} : s = 332;
	{8'd31,8'd78} : s = 453;
	{8'd31,8'd79} : s = 451;
	{8'd31,8'd80} : s = 498;
	{8'd31,8'd81} : s = 176;
	{8'd31,8'd82} : s = 330;
	{8'd31,8'd83} : s = 329;
	{8'd31,8'd84} : s = 440;
	{8'd31,8'd85} : s = 326;
	{8'd31,8'd86} : s = 436;
	{8'd31,8'd87} : s = 434;
	{8'd31,8'd88} : s = 497;
	{8'd31,8'd89} : s = 325;
	{8'd31,8'd90} : s = 433;
	{8'd31,8'd91} : s = 428;
	{8'd31,8'd92} : s = 492;
	{8'd31,8'd93} : s = 426;
	{8'd31,8'd94} : s = 490;
	{8'd31,8'd95} : s = 489;
	{8'd31,8'd96} : s = 508;
	{8'd31,8'd97} : s = 2;
	{8'd31,8'd98} : s = 48;
	{8'd31,8'd99} : s = 40;
	{8'd31,8'd100} : s = 168;
	{8'd31,8'd101} : s = 36;
	{8'd31,8'd102} : s = 164;
	{8'd31,8'd103} : s = 162;
	{8'd31,8'd104} : s = 323;
	{8'd31,8'd105} : s = 34;
	{8'd31,8'd106} : s = 161;
	{8'd31,8'd107} : s = 152;
	{8'd31,8'd108} : s = 312;
	{8'd31,8'd109} : s = 148;
	{8'd31,8'd110} : s = 308;
	{8'd31,8'd111} : s = 306;
	{8'd31,8'd112} : s = 425;
	{8'd31,8'd113} : s = 33;
	{8'd31,8'd114} : s = 146;
	{8'd31,8'd115} : s = 145;
	{8'd31,8'd116} : s = 305;
	{8'd31,8'd117} : s = 140;
	{8'd31,8'd118} : s = 300;
	{8'd31,8'd119} : s = 298;
	{8'd31,8'd120} : s = 422;
	{8'd31,8'd121} : s = 138;
	{8'd31,8'd122} : s = 297;
	{8'd31,8'd123} : s = 294;
	{8'd31,8'd124} : s = 421;
	{8'd31,8'd125} : s = 293;
	{8'd31,8'd126} : s = 419;
	{8'd31,8'd127} : s = 412;
	{8'd31,8'd128} : s = 486;
	{8'd31,8'd129} : s = 24;
	{8'd31,8'd130} : s = 137;
	{8'd31,8'd131} : s = 134;
	{8'd31,8'd132} : s = 291;
	{8'd31,8'd133} : s = 133;
	{8'd31,8'd134} : s = 284;
	{8'd31,8'd135} : s = 282;
	{8'd31,8'd136} : s = 410;
	{8'd31,8'd137} : s = 131;
	{8'd31,8'd138} : s = 281;
	{8'd31,8'd139} : s = 278;
	{8'd31,8'd140} : s = 409;
	{8'd31,8'd141} : s = 277;
	{8'd31,8'd142} : s = 406;
	{8'd31,8'd143} : s = 405;
	{8'd31,8'd144} : s = 485;
	{8'd31,8'd145} : s = 112;
	{8'd31,8'd146} : s = 275;
	{8'd31,8'd147} : s = 270;
	{8'd31,8'd148} : s = 403;
	{8'd31,8'd149} : s = 269;
	{8'd31,8'd150} : s = 398;
	{8'd31,8'd151} : s = 397;
	{8'd31,8'd152} : s = 483;
	{8'd31,8'd153} : s = 267;
	{8'd31,8'd154} : s = 395;
	{8'd31,8'd155} : s = 391;
	{8'd31,8'd156} : s = 476;
	{8'd31,8'd157} : s = 376;
	{8'd31,8'd158} : s = 474;
	{8'd31,8'd159} : s = 473;
	{8'd31,8'd160} : s = 506;
	{8'd31,8'd161} : s = 20;
	{8'd31,8'd162} : s = 104;
	{8'd31,8'd163} : s = 100;
	{8'd31,8'd164} : s = 263;
	{8'd31,8'd165} : s = 98;
	{8'd31,8'd166} : s = 240;
	{8'd31,8'd167} : s = 232;
	{8'd31,8'd168} : s = 372;
	{8'd31,8'd169} : s = 97;
	{8'd31,8'd170} : s = 228;
	{8'd31,8'd171} : s = 226;
	{8'd31,8'd172} : s = 370;
	{8'd31,8'd173} : s = 225;
	{8'd31,8'd174} : s = 369;
	{8'd31,8'd175} : s = 364;
	{8'd31,8'd176} : s = 470;
	{8'd31,8'd177} : s = 88;
	{8'd31,8'd178} : s = 216;
	{8'd31,8'd179} : s = 212;
	{8'd31,8'd180} : s = 362;
	{8'd31,8'd181} : s = 210;
	{8'd31,8'd182} : s = 361;
	{8'd31,8'd183} : s = 358;
	{8'd31,8'd184} : s = 469;
	{8'd31,8'd185} : s = 209;
	{8'd31,8'd186} : s = 357;
	{8'd31,8'd187} : s = 355;
	{8'd31,8'd188} : s = 467;
	{8'd31,8'd189} : s = 348;
	{8'd31,8'd190} : s = 462;
	{8'd31,8'd191} : s = 461;
	{8'd31,8'd192} : s = 505;
	{8'd31,8'd193} : s = 84;
	{8'd31,8'd194} : s = 204;
	{8'd31,8'd195} : s = 202;
	{8'd31,8'd196} : s = 346;
	{8'd31,8'd197} : s = 201;
	{8'd31,8'd198} : s = 345;
	{8'd31,8'd199} : s = 342;
	{8'd31,8'd200} : s = 459;
	{8'd31,8'd201} : s = 198;
	{8'd31,8'd202} : s = 341;
	{8'd31,8'd203} : s = 339;
	{8'd31,8'd204} : s = 455;
	{8'd31,8'd205} : s = 334;
	{8'd31,8'd206} : s = 444;
	{8'd31,8'd207} : s = 442;
	{8'd31,8'd208} : s = 502;
	{8'd31,8'd209} : s = 197;
	{8'd31,8'd210} : s = 333;
	{8'd31,8'd211} : s = 331;
	{8'd31,8'd212} : s = 441;
	{8'd31,8'd213} : s = 327;
	{8'd31,8'd214} : s = 438;
	{8'd31,8'd215} : s = 437;
	{8'd31,8'd216} : s = 501;
	{8'd31,8'd217} : s = 316;
	{8'd31,8'd218} : s = 435;
	{8'd31,8'd219} : s = 430;
	{8'd31,8'd220} : s = 499;
	{8'd31,8'd221} : s = 429;
	{8'd31,8'd222} : s = 494;
	{8'd31,8'd223} : s = 493;
	{8'd31,8'd224} : s = 510;
	{8'd31,8'd225} : s = 1;
	{8'd31,8'd226} : s = 18;
	{8'd31,8'd227} : s = 17;
	{8'd31,8'd228} : s = 82;
	{8'd31,8'd229} : s = 12;
	{8'd31,8'd230} : s = 81;
	{8'd31,8'd231} : s = 76;
	{8'd31,8'd232} : s = 195;
	{8'd31,8'd233} : s = 10;
	{8'd31,8'd234} : s = 74;
	{8'd31,8'd235} : s = 73;
	{8'd31,8'd236} : s = 184;
	{8'd31,8'd237} : s = 70;
	{8'd31,8'd238} : s = 180;
	{8'd31,8'd239} : s = 178;
	{8'd31,8'd240} : s = 314;
	{8'd31,8'd241} : s = 9;
	{8'd31,8'd242} : s = 69;
	{8'd31,8'd243} : s = 67;
	{8'd31,8'd244} : s = 177;
	{8'd31,8'd245} : s = 56;
	{8'd31,8'd246} : s = 172;
	{8'd31,8'd247} : s = 170;
	{8'd31,8'd248} : s = 313;
	{8'd31,8'd249} : s = 52;
	{8'd31,8'd250} : s = 169;
	{8'd31,8'd251} : s = 166;
	{8'd31,8'd252} : s = 310;
	{8'd31,8'd253} : s = 165;
	{8'd31,8'd254} : s = 309;
	{8'd31,8'd255} : s = 307;
	{8'd32,8'd0} : s = 16;
	{8'd32,8'd1} : s = 144;
	{8'd32,8'd2} : s = 136;
	{8'd32,8'd3} : s = 324;
	{8'd32,8'd4} : s = 132;
	{8'd32,8'd5} : s = 322;
	{8'd32,8'd6} : s = 321;
	{8'd32,8'd7} : s = 449;
	{8'd32,8'd8} : s = 130;
	{8'd32,8'd9} : s = 304;
	{8'd32,8'd10} : s = 296;
	{8'd32,8'd11} : s = 432;
	{8'd32,8'd12} : s = 292;
	{8'd32,8'd13} : s = 424;
	{8'd32,8'd14} : s = 420;
	{8'd32,8'd15} : s = 488;
	{8'd32,8'd16} : s = 129;
	{8'd32,8'd17} : s = 290;
	{8'd32,8'd18} : s = 289;
	{8'd32,8'd19} : s = 418;
	{8'd32,8'd20} : s = 280;
	{8'd32,8'd21} : s = 417;
	{8'd32,8'd22} : s = 408;
	{8'd32,8'd23} : s = 484;
	{8'd32,8'd24} : s = 276;
	{8'd32,8'd25} : s = 404;
	{8'd32,8'd26} : s = 402;
	{8'd32,8'd27} : s = 482;
	{8'd32,8'd28} : s = 401;
	{8'd32,8'd29} : s = 481;
	{8'd32,8'd30} : s = 472;
	{8'd32,8'd31} : s = 504;
	{8'd32,8'd32} : s = 4;
	{8'd32,8'd33} : s = 96;
	{8'd32,8'd34} : s = 80;
	{8'd32,8'd35} : s = 274;
	{8'd32,8'd36} : s = 72;
	{8'd32,8'd37} : s = 273;
	{8'd32,8'd38} : s = 268;
	{8'd32,8'd39} : s = 396;
	{8'd32,8'd40} : s = 68;
	{8'd32,8'd41} : s = 266;
	{8'd32,8'd42} : s = 265;
	{8'd32,8'd43} : s = 394;
	{8'd32,8'd44} : s = 262;
	{8'd32,8'd45} : s = 393;
	{8'd32,8'd46} : s = 390;
	{8'd32,8'd47} : s = 468;
	{8'd32,8'd48} : s = 66;
	{8'd32,8'd49} : s = 261;
	{8'd32,8'd50} : s = 259;
	{8'd32,8'd51} : s = 389;
	{8'd32,8'd52} : s = 224;
	{8'd32,8'd53} : s = 387;
	{8'd32,8'd54} : s = 368;
	{8'd32,8'd55} : s = 466;
	{8'd32,8'd56} : s = 208;
	{8'd32,8'd57} : s = 360;
	{8'd32,8'd58} : s = 356;
	{8'd32,8'd59} : s = 465;
	{8'd32,8'd60} : s = 354;
	{8'd32,8'd61} : s = 460;
	{8'd32,8'd62} : s = 458;
	{8'd32,8'd63} : s = 500;
	{8'd32,8'd64} : s = 65;
	{8'd32,8'd65} : s = 200;
	{8'd32,8'd66} : s = 196;
	{8'd32,8'd67} : s = 353;
	{8'd32,8'd68} : s = 194;
	{8'd32,8'd69} : s = 344;
	{8'd32,8'd70} : s = 340;
	{8'd32,8'd71} : s = 457;
	{8'd32,8'd72} : s = 193;
	{8'd32,8'd73} : s = 338;
	{8'd32,8'd74} : s = 337;
	{8'd32,8'd75} : s = 454;
	{8'd32,8'd76} : s = 332;
	{8'd32,8'd77} : s = 453;
	{8'd32,8'd78} : s = 451;
	{8'd32,8'd79} : s = 498;
	{8'd32,8'd80} : s = 176;
	{8'd32,8'd81} : s = 330;
	{8'd32,8'd82} : s = 329;
	{8'd32,8'd83} : s = 440;
	{8'd32,8'd84} : s = 326;
	{8'd32,8'd85} : s = 436;
	{8'd32,8'd86} : s = 434;
	{8'd32,8'd87} : s = 497;
	{8'd32,8'd88} : s = 325;
	{8'd32,8'd89} : s = 433;
	{8'd32,8'd90} : s = 428;
	{8'd32,8'd91} : s = 492;
	{8'd32,8'd92} : s = 426;
	{8'd32,8'd93} : s = 490;
	{8'd32,8'd94} : s = 489;
	{8'd32,8'd95} : s = 508;
	{8'd32,8'd96} : s = 2;
	{8'd32,8'd97} : s = 48;
	{8'd32,8'd98} : s = 40;
	{8'd32,8'd99} : s = 168;
	{8'd32,8'd100} : s = 36;
	{8'd32,8'd101} : s = 164;
	{8'd32,8'd102} : s = 162;
	{8'd32,8'd103} : s = 323;
	{8'd32,8'd104} : s = 34;
	{8'd32,8'd105} : s = 161;
	{8'd32,8'd106} : s = 152;
	{8'd32,8'd107} : s = 312;
	{8'd32,8'd108} : s = 148;
	{8'd32,8'd109} : s = 308;
	{8'd32,8'd110} : s = 306;
	{8'd32,8'd111} : s = 425;
	{8'd32,8'd112} : s = 33;
	{8'd32,8'd113} : s = 146;
	{8'd32,8'd114} : s = 145;
	{8'd32,8'd115} : s = 305;
	{8'd32,8'd116} : s = 140;
	{8'd32,8'd117} : s = 300;
	{8'd32,8'd118} : s = 298;
	{8'd32,8'd119} : s = 422;
	{8'd32,8'd120} : s = 138;
	{8'd32,8'd121} : s = 297;
	{8'd32,8'd122} : s = 294;
	{8'd32,8'd123} : s = 421;
	{8'd32,8'd124} : s = 293;
	{8'd32,8'd125} : s = 419;
	{8'd32,8'd126} : s = 412;
	{8'd32,8'd127} : s = 486;
	{8'd32,8'd128} : s = 24;
	{8'd32,8'd129} : s = 137;
	{8'd32,8'd130} : s = 134;
	{8'd32,8'd131} : s = 291;
	{8'd32,8'd132} : s = 133;
	{8'd32,8'd133} : s = 284;
	{8'd32,8'd134} : s = 282;
	{8'd32,8'd135} : s = 410;
	{8'd32,8'd136} : s = 131;
	{8'd32,8'd137} : s = 281;
	{8'd32,8'd138} : s = 278;
	{8'd32,8'd139} : s = 409;
	{8'd32,8'd140} : s = 277;
	{8'd32,8'd141} : s = 406;
	{8'd32,8'd142} : s = 405;
	{8'd32,8'd143} : s = 485;
	{8'd32,8'd144} : s = 112;
	{8'd32,8'd145} : s = 275;
	{8'd32,8'd146} : s = 270;
	{8'd32,8'd147} : s = 403;
	{8'd32,8'd148} : s = 269;
	{8'd32,8'd149} : s = 398;
	{8'd32,8'd150} : s = 397;
	{8'd32,8'd151} : s = 483;
	{8'd32,8'd152} : s = 267;
	{8'd32,8'd153} : s = 395;
	{8'd32,8'd154} : s = 391;
	{8'd32,8'd155} : s = 476;
	{8'd32,8'd156} : s = 376;
	{8'd32,8'd157} : s = 474;
	{8'd32,8'd158} : s = 473;
	{8'd32,8'd159} : s = 506;
	{8'd32,8'd160} : s = 20;
	{8'd32,8'd161} : s = 104;
	{8'd32,8'd162} : s = 100;
	{8'd32,8'd163} : s = 263;
	{8'd32,8'd164} : s = 98;
	{8'd32,8'd165} : s = 240;
	{8'd32,8'd166} : s = 232;
	{8'd32,8'd167} : s = 372;
	{8'd32,8'd168} : s = 97;
	{8'd32,8'd169} : s = 228;
	{8'd32,8'd170} : s = 226;
	{8'd32,8'd171} : s = 370;
	{8'd32,8'd172} : s = 225;
	{8'd32,8'd173} : s = 369;
	{8'd32,8'd174} : s = 364;
	{8'd32,8'd175} : s = 470;
	{8'd32,8'd176} : s = 88;
	{8'd32,8'd177} : s = 216;
	{8'd32,8'd178} : s = 212;
	{8'd32,8'd179} : s = 362;
	{8'd32,8'd180} : s = 210;
	{8'd32,8'd181} : s = 361;
	{8'd32,8'd182} : s = 358;
	{8'd32,8'd183} : s = 469;
	{8'd32,8'd184} : s = 209;
	{8'd32,8'd185} : s = 357;
	{8'd32,8'd186} : s = 355;
	{8'd32,8'd187} : s = 467;
	{8'd32,8'd188} : s = 348;
	{8'd32,8'd189} : s = 462;
	{8'd32,8'd190} : s = 461;
	{8'd32,8'd191} : s = 505;
	{8'd32,8'd192} : s = 84;
	{8'd32,8'd193} : s = 204;
	{8'd32,8'd194} : s = 202;
	{8'd32,8'd195} : s = 346;
	{8'd32,8'd196} : s = 201;
	{8'd32,8'd197} : s = 345;
	{8'd32,8'd198} : s = 342;
	{8'd32,8'd199} : s = 459;
	{8'd32,8'd200} : s = 198;
	{8'd32,8'd201} : s = 341;
	{8'd32,8'd202} : s = 339;
	{8'd32,8'd203} : s = 455;
	{8'd32,8'd204} : s = 334;
	{8'd32,8'd205} : s = 444;
	{8'd32,8'd206} : s = 442;
	{8'd32,8'd207} : s = 502;
	{8'd32,8'd208} : s = 197;
	{8'd32,8'd209} : s = 333;
	{8'd32,8'd210} : s = 331;
	{8'd32,8'd211} : s = 441;
	{8'd32,8'd212} : s = 327;
	{8'd32,8'd213} : s = 438;
	{8'd32,8'd214} : s = 437;
	{8'd32,8'd215} : s = 501;
	{8'd32,8'd216} : s = 316;
	{8'd32,8'd217} : s = 435;
	{8'd32,8'd218} : s = 430;
	{8'd32,8'd219} : s = 499;
	{8'd32,8'd220} : s = 429;
	{8'd32,8'd221} : s = 494;
	{8'd32,8'd222} : s = 493;
	{8'd32,8'd223} : s = 510;
	{8'd32,8'd224} : s = 1;
	{8'd32,8'd225} : s = 18;
	{8'd32,8'd226} : s = 17;
	{8'd32,8'd227} : s = 82;
	{8'd32,8'd228} : s = 12;
	{8'd32,8'd229} : s = 81;
	{8'd32,8'd230} : s = 76;
	{8'd32,8'd231} : s = 195;
	{8'd32,8'd232} : s = 10;
	{8'd32,8'd233} : s = 74;
	{8'd32,8'd234} : s = 73;
	{8'd32,8'd235} : s = 184;
	{8'd32,8'd236} : s = 70;
	{8'd32,8'd237} : s = 180;
	{8'd32,8'd238} : s = 178;
	{8'd32,8'd239} : s = 314;
	{8'd32,8'd240} : s = 9;
	{8'd32,8'd241} : s = 69;
	{8'd32,8'd242} : s = 67;
	{8'd32,8'd243} : s = 177;
	{8'd32,8'd244} : s = 56;
	{8'd32,8'd245} : s = 172;
	{8'd32,8'd246} : s = 170;
	{8'd32,8'd247} : s = 313;
	{8'd32,8'd248} : s = 52;
	{8'd32,8'd249} : s = 169;
	{8'd32,8'd250} : s = 166;
	{8'd32,8'd251} : s = 310;
	{8'd32,8'd252} : s = 165;
	{8'd32,8'd253} : s = 309;
	{8'd32,8'd254} : s = 307;
	{8'd32,8'd255} : s = 427;
	{8'd33,8'd0} : s = 144;
	{8'd33,8'd1} : s = 136;
	{8'd33,8'd2} : s = 324;
	{8'd33,8'd3} : s = 132;
	{8'd33,8'd4} : s = 322;
	{8'd33,8'd5} : s = 321;
	{8'd33,8'd6} : s = 449;
	{8'd33,8'd7} : s = 130;
	{8'd33,8'd8} : s = 304;
	{8'd33,8'd9} : s = 296;
	{8'd33,8'd10} : s = 432;
	{8'd33,8'd11} : s = 292;
	{8'd33,8'd12} : s = 424;
	{8'd33,8'd13} : s = 420;
	{8'd33,8'd14} : s = 488;
	{8'd33,8'd15} : s = 129;
	{8'd33,8'd16} : s = 290;
	{8'd33,8'd17} : s = 289;
	{8'd33,8'd18} : s = 418;
	{8'd33,8'd19} : s = 280;
	{8'd33,8'd20} : s = 417;
	{8'd33,8'd21} : s = 408;
	{8'd33,8'd22} : s = 484;
	{8'd33,8'd23} : s = 276;
	{8'd33,8'd24} : s = 404;
	{8'd33,8'd25} : s = 402;
	{8'd33,8'd26} : s = 482;
	{8'd33,8'd27} : s = 401;
	{8'd33,8'd28} : s = 481;
	{8'd33,8'd29} : s = 472;
	{8'd33,8'd30} : s = 504;
	{8'd33,8'd31} : s = 4;
	{8'd33,8'd32} : s = 96;
	{8'd33,8'd33} : s = 80;
	{8'd33,8'd34} : s = 274;
	{8'd33,8'd35} : s = 72;
	{8'd33,8'd36} : s = 273;
	{8'd33,8'd37} : s = 268;
	{8'd33,8'd38} : s = 396;
	{8'd33,8'd39} : s = 68;
	{8'd33,8'd40} : s = 266;
	{8'd33,8'd41} : s = 265;
	{8'd33,8'd42} : s = 394;
	{8'd33,8'd43} : s = 262;
	{8'd33,8'd44} : s = 393;
	{8'd33,8'd45} : s = 390;
	{8'd33,8'd46} : s = 468;
	{8'd33,8'd47} : s = 66;
	{8'd33,8'd48} : s = 261;
	{8'd33,8'd49} : s = 259;
	{8'd33,8'd50} : s = 389;
	{8'd33,8'd51} : s = 224;
	{8'd33,8'd52} : s = 387;
	{8'd33,8'd53} : s = 368;
	{8'd33,8'd54} : s = 466;
	{8'd33,8'd55} : s = 208;
	{8'd33,8'd56} : s = 360;
	{8'd33,8'd57} : s = 356;
	{8'd33,8'd58} : s = 465;
	{8'd33,8'd59} : s = 354;
	{8'd33,8'd60} : s = 460;
	{8'd33,8'd61} : s = 458;
	{8'd33,8'd62} : s = 500;
	{8'd33,8'd63} : s = 65;
	{8'd33,8'd64} : s = 200;
	{8'd33,8'd65} : s = 196;
	{8'd33,8'd66} : s = 353;
	{8'd33,8'd67} : s = 194;
	{8'd33,8'd68} : s = 344;
	{8'd33,8'd69} : s = 340;
	{8'd33,8'd70} : s = 457;
	{8'd33,8'd71} : s = 193;
	{8'd33,8'd72} : s = 338;
	{8'd33,8'd73} : s = 337;
	{8'd33,8'd74} : s = 454;
	{8'd33,8'd75} : s = 332;
	{8'd33,8'd76} : s = 453;
	{8'd33,8'd77} : s = 451;
	{8'd33,8'd78} : s = 498;
	{8'd33,8'd79} : s = 176;
	{8'd33,8'd80} : s = 330;
	{8'd33,8'd81} : s = 329;
	{8'd33,8'd82} : s = 440;
	{8'd33,8'd83} : s = 326;
	{8'd33,8'd84} : s = 436;
	{8'd33,8'd85} : s = 434;
	{8'd33,8'd86} : s = 497;
	{8'd33,8'd87} : s = 325;
	{8'd33,8'd88} : s = 433;
	{8'd33,8'd89} : s = 428;
	{8'd33,8'd90} : s = 492;
	{8'd33,8'd91} : s = 426;
	{8'd33,8'd92} : s = 490;
	{8'd33,8'd93} : s = 489;
	{8'd33,8'd94} : s = 508;
	{8'd33,8'd95} : s = 2;
	{8'd33,8'd96} : s = 48;
	{8'd33,8'd97} : s = 40;
	{8'd33,8'd98} : s = 168;
	{8'd33,8'd99} : s = 36;
	{8'd33,8'd100} : s = 164;
	{8'd33,8'd101} : s = 162;
	{8'd33,8'd102} : s = 323;
	{8'd33,8'd103} : s = 34;
	{8'd33,8'd104} : s = 161;
	{8'd33,8'd105} : s = 152;
	{8'd33,8'd106} : s = 312;
	{8'd33,8'd107} : s = 148;
	{8'd33,8'd108} : s = 308;
	{8'd33,8'd109} : s = 306;
	{8'd33,8'd110} : s = 425;
	{8'd33,8'd111} : s = 33;
	{8'd33,8'd112} : s = 146;
	{8'd33,8'd113} : s = 145;
	{8'd33,8'd114} : s = 305;
	{8'd33,8'd115} : s = 140;
	{8'd33,8'd116} : s = 300;
	{8'd33,8'd117} : s = 298;
	{8'd33,8'd118} : s = 422;
	{8'd33,8'd119} : s = 138;
	{8'd33,8'd120} : s = 297;
	{8'd33,8'd121} : s = 294;
	{8'd33,8'd122} : s = 421;
	{8'd33,8'd123} : s = 293;
	{8'd33,8'd124} : s = 419;
	{8'd33,8'd125} : s = 412;
	{8'd33,8'd126} : s = 486;
	{8'd33,8'd127} : s = 24;
	{8'd33,8'd128} : s = 137;
	{8'd33,8'd129} : s = 134;
	{8'd33,8'd130} : s = 291;
	{8'd33,8'd131} : s = 133;
	{8'd33,8'd132} : s = 284;
	{8'd33,8'd133} : s = 282;
	{8'd33,8'd134} : s = 410;
	{8'd33,8'd135} : s = 131;
	{8'd33,8'd136} : s = 281;
	{8'd33,8'd137} : s = 278;
	{8'd33,8'd138} : s = 409;
	{8'd33,8'd139} : s = 277;
	{8'd33,8'd140} : s = 406;
	{8'd33,8'd141} : s = 405;
	{8'd33,8'd142} : s = 485;
	{8'd33,8'd143} : s = 112;
	{8'd33,8'd144} : s = 275;
	{8'd33,8'd145} : s = 270;
	{8'd33,8'd146} : s = 403;
	{8'd33,8'd147} : s = 269;
	{8'd33,8'd148} : s = 398;
	{8'd33,8'd149} : s = 397;
	{8'd33,8'd150} : s = 483;
	{8'd33,8'd151} : s = 267;
	{8'd33,8'd152} : s = 395;
	{8'd33,8'd153} : s = 391;
	{8'd33,8'd154} : s = 476;
	{8'd33,8'd155} : s = 376;
	{8'd33,8'd156} : s = 474;
	{8'd33,8'd157} : s = 473;
	{8'd33,8'd158} : s = 506;
	{8'd33,8'd159} : s = 20;
	{8'd33,8'd160} : s = 104;
	{8'd33,8'd161} : s = 100;
	{8'd33,8'd162} : s = 263;
	{8'd33,8'd163} : s = 98;
	{8'd33,8'd164} : s = 240;
	{8'd33,8'd165} : s = 232;
	{8'd33,8'd166} : s = 372;
	{8'd33,8'd167} : s = 97;
	{8'd33,8'd168} : s = 228;
	{8'd33,8'd169} : s = 226;
	{8'd33,8'd170} : s = 370;
	{8'd33,8'd171} : s = 225;
	{8'd33,8'd172} : s = 369;
	{8'd33,8'd173} : s = 364;
	{8'd33,8'd174} : s = 470;
	{8'd33,8'd175} : s = 88;
	{8'd33,8'd176} : s = 216;
	{8'd33,8'd177} : s = 212;
	{8'd33,8'd178} : s = 362;
	{8'd33,8'd179} : s = 210;
	{8'd33,8'd180} : s = 361;
	{8'd33,8'd181} : s = 358;
	{8'd33,8'd182} : s = 469;
	{8'd33,8'd183} : s = 209;
	{8'd33,8'd184} : s = 357;
	{8'd33,8'd185} : s = 355;
	{8'd33,8'd186} : s = 467;
	{8'd33,8'd187} : s = 348;
	{8'd33,8'd188} : s = 462;
	{8'd33,8'd189} : s = 461;
	{8'd33,8'd190} : s = 505;
	{8'd33,8'd191} : s = 84;
	{8'd33,8'd192} : s = 204;
	{8'd33,8'd193} : s = 202;
	{8'd33,8'd194} : s = 346;
	{8'd33,8'd195} : s = 201;
	{8'd33,8'd196} : s = 345;
	{8'd33,8'd197} : s = 342;
	{8'd33,8'd198} : s = 459;
	{8'd33,8'd199} : s = 198;
	{8'd33,8'd200} : s = 341;
	{8'd33,8'd201} : s = 339;
	{8'd33,8'd202} : s = 455;
	{8'd33,8'd203} : s = 334;
	{8'd33,8'd204} : s = 444;
	{8'd33,8'd205} : s = 442;
	{8'd33,8'd206} : s = 502;
	{8'd33,8'd207} : s = 197;
	{8'd33,8'd208} : s = 333;
	{8'd33,8'd209} : s = 331;
	{8'd33,8'd210} : s = 441;
	{8'd33,8'd211} : s = 327;
	{8'd33,8'd212} : s = 438;
	{8'd33,8'd213} : s = 437;
	{8'd33,8'd214} : s = 501;
	{8'd33,8'd215} : s = 316;
	{8'd33,8'd216} : s = 435;
	{8'd33,8'd217} : s = 430;
	{8'd33,8'd218} : s = 499;
	{8'd33,8'd219} : s = 429;
	{8'd33,8'd220} : s = 494;
	{8'd33,8'd221} : s = 493;
	{8'd33,8'd222} : s = 510;
	{8'd33,8'd223} : s = 1;
	{8'd33,8'd224} : s = 18;
	{8'd33,8'd225} : s = 17;
	{8'd33,8'd226} : s = 82;
	{8'd33,8'd227} : s = 12;
	{8'd33,8'd228} : s = 81;
	{8'd33,8'd229} : s = 76;
	{8'd33,8'd230} : s = 195;
	{8'd33,8'd231} : s = 10;
	{8'd33,8'd232} : s = 74;
	{8'd33,8'd233} : s = 73;
	{8'd33,8'd234} : s = 184;
	{8'd33,8'd235} : s = 70;
	{8'd33,8'd236} : s = 180;
	{8'd33,8'd237} : s = 178;
	{8'd33,8'd238} : s = 314;
	{8'd33,8'd239} : s = 9;
	{8'd33,8'd240} : s = 69;
	{8'd33,8'd241} : s = 67;
	{8'd33,8'd242} : s = 177;
	{8'd33,8'd243} : s = 56;
	{8'd33,8'd244} : s = 172;
	{8'd33,8'd245} : s = 170;
	{8'd33,8'd246} : s = 313;
	{8'd33,8'd247} : s = 52;
	{8'd33,8'd248} : s = 169;
	{8'd33,8'd249} : s = 166;
	{8'd33,8'd250} : s = 310;
	{8'd33,8'd251} : s = 165;
	{8'd33,8'd252} : s = 309;
	{8'd33,8'd253} : s = 307;
	{8'd33,8'd254} : s = 427;
	{8'd33,8'd255} : s = 6;
	{8'd34,8'd0} : s = 136;
	{8'd34,8'd1} : s = 324;
	{8'd34,8'd2} : s = 132;
	{8'd34,8'd3} : s = 322;
	{8'd34,8'd4} : s = 321;
	{8'd34,8'd5} : s = 449;
	{8'd34,8'd6} : s = 130;
	{8'd34,8'd7} : s = 304;
	{8'd34,8'd8} : s = 296;
	{8'd34,8'd9} : s = 432;
	{8'd34,8'd10} : s = 292;
	{8'd34,8'd11} : s = 424;
	{8'd34,8'd12} : s = 420;
	{8'd34,8'd13} : s = 488;
	{8'd34,8'd14} : s = 129;
	{8'd34,8'd15} : s = 290;
	{8'd34,8'd16} : s = 289;
	{8'd34,8'd17} : s = 418;
	{8'd34,8'd18} : s = 280;
	{8'd34,8'd19} : s = 417;
	{8'd34,8'd20} : s = 408;
	{8'd34,8'd21} : s = 484;
	{8'd34,8'd22} : s = 276;
	{8'd34,8'd23} : s = 404;
	{8'd34,8'd24} : s = 402;
	{8'd34,8'd25} : s = 482;
	{8'd34,8'd26} : s = 401;
	{8'd34,8'd27} : s = 481;
	{8'd34,8'd28} : s = 472;
	{8'd34,8'd29} : s = 504;
	{8'd34,8'd30} : s = 4;
	{8'd34,8'd31} : s = 96;
	{8'd34,8'd32} : s = 80;
	{8'd34,8'd33} : s = 274;
	{8'd34,8'd34} : s = 72;
	{8'd34,8'd35} : s = 273;
	{8'd34,8'd36} : s = 268;
	{8'd34,8'd37} : s = 396;
	{8'd34,8'd38} : s = 68;
	{8'd34,8'd39} : s = 266;
	{8'd34,8'd40} : s = 265;
	{8'd34,8'd41} : s = 394;
	{8'd34,8'd42} : s = 262;
	{8'd34,8'd43} : s = 393;
	{8'd34,8'd44} : s = 390;
	{8'd34,8'd45} : s = 468;
	{8'd34,8'd46} : s = 66;
	{8'd34,8'd47} : s = 261;
	{8'd34,8'd48} : s = 259;
	{8'd34,8'd49} : s = 389;
	{8'd34,8'd50} : s = 224;
	{8'd34,8'd51} : s = 387;
	{8'd34,8'd52} : s = 368;
	{8'd34,8'd53} : s = 466;
	{8'd34,8'd54} : s = 208;
	{8'd34,8'd55} : s = 360;
	{8'd34,8'd56} : s = 356;
	{8'd34,8'd57} : s = 465;
	{8'd34,8'd58} : s = 354;
	{8'd34,8'd59} : s = 460;
	{8'd34,8'd60} : s = 458;
	{8'd34,8'd61} : s = 500;
	{8'd34,8'd62} : s = 65;
	{8'd34,8'd63} : s = 200;
	{8'd34,8'd64} : s = 196;
	{8'd34,8'd65} : s = 353;
	{8'd34,8'd66} : s = 194;
	{8'd34,8'd67} : s = 344;
	{8'd34,8'd68} : s = 340;
	{8'd34,8'd69} : s = 457;
	{8'd34,8'd70} : s = 193;
	{8'd34,8'd71} : s = 338;
	{8'd34,8'd72} : s = 337;
	{8'd34,8'd73} : s = 454;
	{8'd34,8'd74} : s = 332;
	{8'd34,8'd75} : s = 453;
	{8'd34,8'd76} : s = 451;
	{8'd34,8'd77} : s = 498;
	{8'd34,8'd78} : s = 176;
	{8'd34,8'd79} : s = 330;
	{8'd34,8'd80} : s = 329;
	{8'd34,8'd81} : s = 440;
	{8'd34,8'd82} : s = 326;
	{8'd34,8'd83} : s = 436;
	{8'd34,8'd84} : s = 434;
	{8'd34,8'd85} : s = 497;
	{8'd34,8'd86} : s = 325;
	{8'd34,8'd87} : s = 433;
	{8'd34,8'd88} : s = 428;
	{8'd34,8'd89} : s = 492;
	{8'd34,8'd90} : s = 426;
	{8'd34,8'd91} : s = 490;
	{8'd34,8'd92} : s = 489;
	{8'd34,8'd93} : s = 508;
	{8'd34,8'd94} : s = 2;
	{8'd34,8'd95} : s = 48;
	{8'd34,8'd96} : s = 40;
	{8'd34,8'd97} : s = 168;
	{8'd34,8'd98} : s = 36;
	{8'd34,8'd99} : s = 164;
	{8'd34,8'd100} : s = 162;
	{8'd34,8'd101} : s = 323;
	{8'd34,8'd102} : s = 34;
	{8'd34,8'd103} : s = 161;
	{8'd34,8'd104} : s = 152;
	{8'd34,8'd105} : s = 312;
	{8'd34,8'd106} : s = 148;
	{8'd34,8'd107} : s = 308;
	{8'd34,8'd108} : s = 306;
	{8'd34,8'd109} : s = 425;
	{8'd34,8'd110} : s = 33;
	{8'd34,8'd111} : s = 146;
	{8'd34,8'd112} : s = 145;
	{8'd34,8'd113} : s = 305;
	{8'd34,8'd114} : s = 140;
	{8'd34,8'd115} : s = 300;
	{8'd34,8'd116} : s = 298;
	{8'd34,8'd117} : s = 422;
	{8'd34,8'd118} : s = 138;
	{8'd34,8'd119} : s = 297;
	{8'd34,8'd120} : s = 294;
	{8'd34,8'd121} : s = 421;
	{8'd34,8'd122} : s = 293;
	{8'd34,8'd123} : s = 419;
	{8'd34,8'd124} : s = 412;
	{8'd34,8'd125} : s = 486;
	{8'd34,8'd126} : s = 24;
	{8'd34,8'd127} : s = 137;
	{8'd34,8'd128} : s = 134;
	{8'd34,8'd129} : s = 291;
	{8'd34,8'd130} : s = 133;
	{8'd34,8'd131} : s = 284;
	{8'd34,8'd132} : s = 282;
	{8'd34,8'd133} : s = 410;
	{8'd34,8'd134} : s = 131;
	{8'd34,8'd135} : s = 281;
	{8'd34,8'd136} : s = 278;
	{8'd34,8'd137} : s = 409;
	{8'd34,8'd138} : s = 277;
	{8'd34,8'd139} : s = 406;
	{8'd34,8'd140} : s = 405;
	{8'd34,8'd141} : s = 485;
	{8'd34,8'd142} : s = 112;
	{8'd34,8'd143} : s = 275;
	{8'd34,8'd144} : s = 270;
	{8'd34,8'd145} : s = 403;
	{8'd34,8'd146} : s = 269;
	{8'd34,8'd147} : s = 398;
	{8'd34,8'd148} : s = 397;
	{8'd34,8'd149} : s = 483;
	{8'd34,8'd150} : s = 267;
	{8'd34,8'd151} : s = 395;
	{8'd34,8'd152} : s = 391;
	{8'd34,8'd153} : s = 476;
	{8'd34,8'd154} : s = 376;
	{8'd34,8'd155} : s = 474;
	{8'd34,8'd156} : s = 473;
	{8'd34,8'd157} : s = 506;
	{8'd34,8'd158} : s = 20;
	{8'd34,8'd159} : s = 104;
	{8'd34,8'd160} : s = 100;
	{8'd34,8'd161} : s = 263;
	{8'd34,8'd162} : s = 98;
	{8'd34,8'd163} : s = 240;
	{8'd34,8'd164} : s = 232;
	{8'd34,8'd165} : s = 372;
	{8'd34,8'd166} : s = 97;
	{8'd34,8'd167} : s = 228;
	{8'd34,8'd168} : s = 226;
	{8'd34,8'd169} : s = 370;
	{8'd34,8'd170} : s = 225;
	{8'd34,8'd171} : s = 369;
	{8'd34,8'd172} : s = 364;
	{8'd34,8'd173} : s = 470;
	{8'd34,8'd174} : s = 88;
	{8'd34,8'd175} : s = 216;
	{8'd34,8'd176} : s = 212;
	{8'd34,8'd177} : s = 362;
	{8'd34,8'd178} : s = 210;
	{8'd34,8'd179} : s = 361;
	{8'd34,8'd180} : s = 358;
	{8'd34,8'd181} : s = 469;
	{8'd34,8'd182} : s = 209;
	{8'd34,8'd183} : s = 357;
	{8'd34,8'd184} : s = 355;
	{8'd34,8'd185} : s = 467;
	{8'd34,8'd186} : s = 348;
	{8'd34,8'd187} : s = 462;
	{8'd34,8'd188} : s = 461;
	{8'd34,8'd189} : s = 505;
	{8'd34,8'd190} : s = 84;
	{8'd34,8'd191} : s = 204;
	{8'd34,8'd192} : s = 202;
	{8'd34,8'd193} : s = 346;
	{8'd34,8'd194} : s = 201;
	{8'd34,8'd195} : s = 345;
	{8'd34,8'd196} : s = 342;
	{8'd34,8'd197} : s = 459;
	{8'd34,8'd198} : s = 198;
	{8'd34,8'd199} : s = 341;
	{8'd34,8'd200} : s = 339;
	{8'd34,8'd201} : s = 455;
	{8'd34,8'd202} : s = 334;
	{8'd34,8'd203} : s = 444;
	{8'd34,8'd204} : s = 442;
	{8'd34,8'd205} : s = 502;
	{8'd34,8'd206} : s = 197;
	{8'd34,8'd207} : s = 333;
	{8'd34,8'd208} : s = 331;
	{8'd34,8'd209} : s = 441;
	{8'd34,8'd210} : s = 327;
	{8'd34,8'd211} : s = 438;
	{8'd34,8'd212} : s = 437;
	{8'd34,8'd213} : s = 501;
	{8'd34,8'd214} : s = 316;
	{8'd34,8'd215} : s = 435;
	{8'd34,8'd216} : s = 430;
	{8'd34,8'd217} : s = 499;
	{8'd34,8'd218} : s = 429;
	{8'd34,8'd219} : s = 494;
	{8'd34,8'd220} : s = 493;
	{8'd34,8'd221} : s = 510;
	{8'd34,8'd222} : s = 1;
	{8'd34,8'd223} : s = 18;
	{8'd34,8'd224} : s = 17;
	{8'd34,8'd225} : s = 82;
	{8'd34,8'd226} : s = 12;
	{8'd34,8'd227} : s = 81;
	{8'd34,8'd228} : s = 76;
	{8'd34,8'd229} : s = 195;
	{8'd34,8'd230} : s = 10;
	{8'd34,8'd231} : s = 74;
	{8'd34,8'd232} : s = 73;
	{8'd34,8'd233} : s = 184;
	{8'd34,8'd234} : s = 70;
	{8'd34,8'd235} : s = 180;
	{8'd34,8'd236} : s = 178;
	{8'd34,8'd237} : s = 314;
	{8'd34,8'd238} : s = 9;
	{8'd34,8'd239} : s = 69;
	{8'd34,8'd240} : s = 67;
	{8'd34,8'd241} : s = 177;
	{8'd34,8'd242} : s = 56;
	{8'd34,8'd243} : s = 172;
	{8'd34,8'd244} : s = 170;
	{8'd34,8'd245} : s = 313;
	{8'd34,8'd246} : s = 52;
	{8'd34,8'd247} : s = 169;
	{8'd34,8'd248} : s = 166;
	{8'd34,8'd249} : s = 310;
	{8'd34,8'd250} : s = 165;
	{8'd34,8'd251} : s = 309;
	{8'd34,8'd252} : s = 307;
	{8'd34,8'd253} : s = 427;
	{8'd34,8'd254} : s = 6;
	{8'd34,8'd255} : s = 50;
	{8'd35,8'd0} : s = 324;
	{8'd35,8'd1} : s = 132;
	{8'd35,8'd2} : s = 322;
	{8'd35,8'd3} : s = 321;
	{8'd35,8'd4} : s = 449;
	{8'd35,8'd5} : s = 130;
	{8'd35,8'd6} : s = 304;
	{8'd35,8'd7} : s = 296;
	{8'd35,8'd8} : s = 432;
	{8'd35,8'd9} : s = 292;
	{8'd35,8'd10} : s = 424;
	{8'd35,8'd11} : s = 420;
	{8'd35,8'd12} : s = 488;
	{8'd35,8'd13} : s = 129;
	{8'd35,8'd14} : s = 290;
	{8'd35,8'd15} : s = 289;
	{8'd35,8'd16} : s = 418;
	{8'd35,8'd17} : s = 280;
	{8'd35,8'd18} : s = 417;
	{8'd35,8'd19} : s = 408;
	{8'd35,8'd20} : s = 484;
	{8'd35,8'd21} : s = 276;
	{8'd35,8'd22} : s = 404;
	{8'd35,8'd23} : s = 402;
	{8'd35,8'd24} : s = 482;
	{8'd35,8'd25} : s = 401;
	{8'd35,8'd26} : s = 481;
	{8'd35,8'd27} : s = 472;
	{8'd35,8'd28} : s = 504;
	{8'd35,8'd29} : s = 4;
	{8'd35,8'd30} : s = 96;
	{8'd35,8'd31} : s = 80;
	{8'd35,8'd32} : s = 274;
	{8'd35,8'd33} : s = 72;
	{8'd35,8'd34} : s = 273;
	{8'd35,8'd35} : s = 268;
	{8'd35,8'd36} : s = 396;
	{8'd35,8'd37} : s = 68;
	{8'd35,8'd38} : s = 266;
	{8'd35,8'd39} : s = 265;
	{8'd35,8'd40} : s = 394;
	{8'd35,8'd41} : s = 262;
	{8'd35,8'd42} : s = 393;
	{8'd35,8'd43} : s = 390;
	{8'd35,8'd44} : s = 468;
	{8'd35,8'd45} : s = 66;
	{8'd35,8'd46} : s = 261;
	{8'd35,8'd47} : s = 259;
	{8'd35,8'd48} : s = 389;
	{8'd35,8'd49} : s = 224;
	{8'd35,8'd50} : s = 387;
	{8'd35,8'd51} : s = 368;
	{8'd35,8'd52} : s = 466;
	{8'd35,8'd53} : s = 208;
	{8'd35,8'd54} : s = 360;
	{8'd35,8'd55} : s = 356;
	{8'd35,8'd56} : s = 465;
	{8'd35,8'd57} : s = 354;
	{8'd35,8'd58} : s = 460;
	{8'd35,8'd59} : s = 458;
	{8'd35,8'd60} : s = 500;
	{8'd35,8'd61} : s = 65;
	{8'd35,8'd62} : s = 200;
	{8'd35,8'd63} : s = 196;
	{8'd35,8'd64} : s = 353;
	{8'd35,8'd65} : s = 194;
	{8'd35,8'd66} : s = 344;
	{8'd35,8'd67} : s = 340;
	{8'd35,8'd68} : s = 457;
	{8'd35,8'd69} : s = 193;
	{8'd35,8'd70} : s = 338;
	{8'd35,8'd71} : s = 337;
	{8'd35,8'd72} : s = 454;
	{8'd35,8'd73} : s = 332;
	{8'd35,8'd74} : s = 453;
	{8'd35,8'd75} : s = 451;
	{8'd35,8'd76} : s = 498;
	{8'd35,8'd77} : s = 176;
	{8'd35,8'd78} : s = 330;
	{8'd35,8'd79} : s = 329;
	{8'd35,8'd80} : s = 440;
	{8'd35,8'd81} : s = 326;
	{8'd35,8'd82} : s = 436;
	{8'd35,8'd83} : s = 434;
	{8'd35,8'd84} : s = 497;
	{8'd35,8'd85} : s = 325;
	{8'd35,8'd86} : s = 433;
	{8'd35,8'd87} : s = 428;
	{8'd35,8'd88} : s = 492;
	{8'd35,8'd89} : s = 426;
	{8'd35,8'd90} : s = 490;
	{8'd35,8'd91} : s = 489;
	{8'd35,8'd92} : s = 508;
	{8'd35,8'd93} : s = 2;
	{8'd35,8'd94} : s = 48;
	{8'd35,8'd95} : s = 40;
	{8'd35,8'd96} : s = 168;
	{8'd35,8'd97} : s = 36;
	{8'd35,8'd98} : s = 164;
	{8'd35,8'd99} : s = 162;
	{8'd35,8'd100} : s = 323;
	{8'd35,8'd101} : s = 34;
	{8'd35,8'd102} : s = 161;
	{8'd35,8'd103} : s = 152;
	{8'd35,8'd104} : s = 312;
	{8'd35,8'd105} : s = 148;
	{8'd35,8'd106} : s = 308;
	{8'd35,8'd107} : s = 306;
	{8'd35,8'd108} : s = 425;
	{8'd35,8'd109} : s = 33;
	{8'd35,8'd110} : s = 146;
	{8'd35,8'd111} : s = 145;
	{8'd35,8'd112} : s = 305;
	{8'd35,8'd113} : s = 140;
	{8'd35,8'd114} : s = 300;
	{8'd35,8'd115} : s = 298;
	{8'd35,8'd116} : s = 422;
	{8'd35,8'd117} : s = 138;
	{8'd35,8'd118} : s = 297;
	{8'd35,8'd119} : s = 294;
	{8'd35,8'd120} : s = 421;
	{8'd35,8'd121} : s = 293;
	{8'd35,8'd122} : s = 419;
	{8'd35,8'd123} : s = 412;
	{8'd35,8'd124} : s = 486;
	{8'd35,8'd125} : s = 24;
	{8'd35,8'd126} : s = 137;
	{8'd35,8'd127} : s = 134;
	{8'd35,8'd128} : s = 291;
	{8'd35,8'd129} : s = 133;
	{8'd35,8'd130} : s = 284;
	{8'd35,8'd131} : s = 282;
	{8'd35,8'd132} : s = 410;
	{8'd35,8'd133} : s = 131;
	{8'd35,8'd134} : s = 281;
	{8'd35,8'd135} : s = 278;
	{8'd35,8'd136} : s = 409;
	{8'd35,8'd137} : s = 277;
	{8'd35,8'd138} : s = 406;
	{8'd35,8'd139} : s = 405;
	{8'd35,8'd140} : s = 485;
	{8'd35,8'd141} : s = 112;
	{8'd35,8'd142} : s = 275;
	{8'd35,8'd143} : s = 270;
	{8'd35,8'd144} : s = 403;
	{8'd35,8'd145} : s = 269;
	{8'd35,8'd146} : s = 398;
	{8'd35,8'd147} : s = 397;
	{8'd35,8'd148} : s = 483;
	{8'd35,8'd149} : s = 267;
	{8'd35,8'd150} : s = 395;
	{8'd35,8'd151} : s = 391;
	{8'd35,8'd152} : s = 476;
	{8'd35,8'd153} : s = 376;
	{8'd35,8'd154} : s = 474;
	{8'd35,8'd155} : s = 473;
	{8'd35,8'd156} : s = 506;
	{8'd35,8'd157} : s = 20;
	{8'd35,8'd158} : s = 104;
	{8'd35,8'd159} : s = 100;
	{8'd35,8'd160} : s = 263;
	{8'd35,8'd161} : s = 98;
	{8'd35,8'd162} : s = 240;
	{8'd35,8'd163} : s = 232;
	{8'd35,8'd164} : s = 372;
	{8'd35,8'd165} : s = 97;
	{8'd35,8'd166} : s = 228;
	{8'd35,8'd167} : s = 226;
	{8'd35,8'd168} : s = 370;
	{8'd35,8'd169} : s = 225;
	{8'd35,8'd170} : s = 369;
	{8'd35,8'd171} : s = 364;
	{8'd35,8'd172} : s = 470;
	{8'd35,8'd173} : s = 88;
	{8'd35,8'd174} : s = 216;
	{8'd35,8'd175} : s = 212;
	{8'd35,8'd176} : s = 362;
	{8'd35,8'd177} : s = 210;
	{8'd35,8'd178} : s = 361;
	{8'd35,8'd179} : s = 358;
	{8'd35,8'd180} : s = 469;
	{8'd35,8'd181} : s = 209;
	{8'd35,8'd182} : s = 357;
	{8'd35,8'd183} : s = 355;
	{8'd35,8'd184} : s = 467;
	{8'd35,8'd185} : s = 348;
	{8'd35,8'd186} : s = 462;
	{8'd35,8'd187} : s = 461;
	{8'd35,8'd188} : s = 505;
	{8'd35,8'd189} : s = 84;
	{8'd35,8'd190} : s = 204;
	{8'd35,8'd191} : s = 202;
	{8'd35,8'd192} : s = 346;
	{8'd35,8'd193} : s = 201;
	{8'd35,8'd194} : s = 345;
	{8'd35,8'd195} : s = 342;
	{8'd35,8'd196} : s = 459;
	{8'd35,8'd197} : s = 198;
	{8'd35,8'd198} : s = 341;
	{8'd35,8'd199} : s = 339;
	{8'd35,8'd200} : s = 455;
	{8'd35,8'd201} : s = 334;
	{8'd35,8'd202} : s = 444;
	{8'd35,8'd203} : s = 442;
	{8'd35,8'd204} : s = 502;
	{8'd35,8'd205} : s = 197;
	{8'd35,8'd206} : s = 333;
	{8'd35,8'd207} : s = 331;
	{8'd35,8'd208} : s = 441;
	{8'd35,8'd209} : s = 327;
	{8'd35,8'd210} : s = 438;
	{8'd35,8'd211} : s = 437;
	{8'd35,8'd212} : s = 501;
	{8'd35,8'd213} : s = 316;
	{8'd35,8'd214} : s = 435;
	{8'd35,8'd215} : s = 430;
	{8'd35,8'd216} : s = 499;
	{8'd35,8'd217} : s = 429;
	{8'd35,8'd218} : s = 494;
	{8'd35,8'd219} : s = 493;
	{8'd35,8'd220} : s = 510;
	{8'd35,8'd221} : s = 1;
	{8'd35,8'd222} : s = 18;
	{8'd35,8'd223} : s = 17;
	{8'd35,8'd224} : s = 82;
	{8'd35,8'd225} : s = 12;
	{8'd35,8'd226} : s = 81;
	{8'd35,8'd227} : s = 76;
	{8'd35,8'd228} : s = 195;
	{8'd35,8'd229} : s = 10;
	{8'd35,8'd230} : s = 74;
	{8'd35,8'd231} : s = 73;
	{8'd35,8'd232} : s = 184;
	{8'd35,8'd233} : s = 70;
	{8'd35,8'd234} : s = 180;
	{8'd35,8'd235} : s = 178;
	{8'd35,8'd236} : s = 314;
	{8'd35,8'd237} : s = 9;
	{8'd35,8'd238} : s = 69;
	{8'd35,8'd239} : s = 67;
	{8'd35,8'd240} : s = 177;
	{8'd35,8'd241} : s = 56;
	{8'd35,8'd242} : s = 172;
	{8'd35,8'd243} : s = 170;
	{8'd35,8'd244} : s = 313;
	{8'd35,8'd245} : s = 52;
	{8'd35,8'd246} : s = 169;
	{8'd35,8'd247} : s = 166;
	{8'd35,8'd248} : s = 310;
	{8'd35,8'd249} : s = 165;
	{8'd35,8'd250} : s = 309;
	{8'd35,8'd251} : s = 307;
	{8'd35,8'd252} : s = 427;
	{8'd35,8'd253} : s = 6;
	{8'd35,8'd254} : s = 50;
	{8'd35,8'd255} : s = 49;
	{8'd36,8'd0} : s = 132;
	{8'd36,8'd1} : s = 322;
	{8'd36,8'd2} : s = 321;
	{8'd36,8'd3} : s = 449;
	{8'd36,8'd4} : s = 130;
	{8'd36,8'd5} : s = 304;
	{8'd36,8'd6} : s = 296;
	{8'd36,8'd7} : s = 432;
	{8'd36,8'd8} : s = 292;
	{8'd36,8'd9} : s = 424;
	{8'd36,8'd10} : s = 420;
	{8'd36,8'd11} : s = 488;
	{8'd36,8'd12} : s = 129;
	{8'd36,8'd13} : s = 290;
	{8'd36,8'd14} : s = 289;
	{8'd36,8'd15} : s = 418;
	{8'd36,8'd16} : s = 280;
	{8'd36,8'd17} : s = 417;
	{8'd36,8'd18} : s = 408;
	{8'd36,8'd19} : s = 484;
	{8'd36,8'd20} : s = 276;
	{8'd36,8'd21} : s = 404;
	{8'd36,8'd22} : s = 402;
	{8'd36,8'd23} : s = 482;
	{8'd36,8'd24} : s = 401;
	{8'd36,8'd25} : s = 481;
	{8'd36,8'd26} : s = 472;
	{8'd36,8'd27} : s = 504;
	{8'd36,8'd28} : s = 4;
	{8'd36,8'd29} : s = 96;
	{8'd36,8'd30} : s = 80;
	{8'd36,8'd31} : s = 274;
	{8'd36,8'd32} : s = 72;
	{8'd36,8'd33} : s = 273;
	{8'd36,8'd34} : s = 268;
	{8'd36,8'd35} : s = 396;
	{8'd36,8'd36} : s = 68;
	{8'd36,8'd37} : s = 266;
	{8'd36,8'd38} : s = 265;
	{8'd36,8'd39} : s = 394;
	{8'd36,8'd40} : s = 262;
	{8'd36,8'd41} : s = 393;
	{8'd36,8'd42} : s = 390;
	{8'd36,8'd43} : s = 468;
	{8'd36,8'd44} : s = 66;
	{8'd36,8'd45} : s = 261;
	{8'd36,8'd46} : s = 259;
	{8'd36,8'd47} : s = 389;
	{8'd36,8'd48} : s = 224;
	{8'd36,8'd49} : s = 387;
	{8'd36,8'd50} : s = 368;
	{8'd36,8'd51} : s = 466;
	{8'd36,8'd52} : s = 208;
	{8'd36,8'd53} : s = 360;
	{8'd36,8'd54} : s = 356;
	{8'd36,8'd55} : s = 465;
	{8'd36,8'd56} : s = 354;
	{8'd36,8'd57} : s = 460;
	{8'd36,8'd58} : s = 458;
	{8'd36,8'd59} : s = 500;
	{8'd36,8'd60} : s = 65;
	{8'd36,8'd61} : s = 200;
	{8'd36,8'd62} : s = 196;
	{8'd36,8'd63} : s = 353;
	{8'd36,8'd64} : s = 194;
	{8'd36,8'd65} : s = 344;
	{8'd36,8'd66} : s = 340;
	{8'd36,8'd67} : s = 457;
	{8'd36,8'd68} : s = 193;
	{8'd36,8'd69} : s = 338;
	{8'd36,8'd70} : s = 337;
	{8'd36,8'd71} : s = 454;
	{8'd36,8'd72} : s = 332;
	{8'd36,8'd73} : s = 453;
	{8'd36,8'd74} : s = 451;
	{8'd36,8'd75} : s = 498;
	{8'd36,8'd76} : s = 176;
	{8'd36,8'd77} : s = 330;
	{8'd36,8'd78} : s = 329;
	{8'd36,8'd79} : s = 440;
	{8'd36,8'd80} : s = 326;
	{8'd36,8'd81} : s = 436;
	{8'd36,8'd82} : s = 434;
	{8'd36,8'd83} : s = 497;
	{8'd36,8'd84} : s = 325;
	{8'd36,8'd85} : s = 433;
	{8'd36,8'd86} : s = 428;
	{8'd36,8'd87} : s = 492;
	{8'd36,8'd88} : s = 426;
	{8'd36,8'd89} : s = 490;
	{8'd36,8'd90} : s = 489;
	{8'd36,8'd91} : s = 508;
	{8'd36,8'd92} : s = 2;
	{8'd36,8'd93} : s = 48;
	{8'd36,8'd94} : s = 40;
	{8'd36,8'd95} : s = 168;
	{8'd36,8'd96} : s = 36;
	{8'd36,8'd97} : s = 164;
	{8'd36,8'd98} : s = 162;
	{8'd36,8'd99} : s = 323;
	{8'd36,8'd100} : s = 34;
	{8'd36,8'd101} : s = 161;
	{8'd36,8'd102} : s = 152;
	{8'd36,8'd103} : s = 312;
	{8'd36,8'd104} : s = 148;
	{8'd36,8'd105} : s = 308;
	{8'd36,8'd106} : s = 306;
	{8'd36,8'd107} : s = 425;
	{8'd36,8'd108} : s = 33;
	{8'd36,8'd109} : s = 146;
	{8'd36,8'd110} : s = 145;
	{8'd36,8'd111} : s = 305;
	{8'd36,8'd112} : s = 140;
	{8'd36,8'd113} : s = 300;
	{8'd36,8'd114} : s = 298;
	{8'd36,8'd115} : s = 422;
	{8'd36,8'd116} : s = 138;
	{8'd36,8'd117} : s = 297;
	{8'd36,8'd118} : s = 294;
	{8'd36,8'd119} : s = 421;
	{8'd36,8'd120} : s = 293;
	{8'd36,8'd121} : s = 419;
	{8'd36,8'd122} : s = 412;
	{8'd36,8'd123} : s = 486;
	{8'd36,8'd124} : s = 24;
	{8'd36,8'd125} : s = 137;
	{8'd36,8'd126} : s = 134;
	{8'd36,8'd127} : s = 291;
	{8'd36,8'd128} : s = 133;
	{8'd36,8'd129} : s = 284;
	{8'd36,8'd130} : s = 282;
	{8'd36,8'd131} : s = 410;
	{8'd36,8'd132} : s = 131;
	{8'd36,8'd133} : s = 281;
	{8'd36,8'd134} : s = 278;
	{8'd36,8'd135} : s = 409;
	{8'd36,8'd136} : s = 277;
	{8'd36,8'd137} : s = 406;
	{8'd36,8'd138} : s = 405;
	{8'd36,8'd139} : s = 485;
	{8'd36,8'd140} : s = 112;
	{8'd36,8'd141} : s = 275;
	{8'd36,8'd142} : s = 270;
	{8'd36,8'd143} : s = 403;
	{8'd36,8'd144} : s = 269;
	{8'd36,8'd145} : s = 398;
	{8'd36,8'd146} : s = 397;
	{8'd36,8'd147} : s = 483;
	{8'd36,8'd148} : s = 267;
	{8'd36,8'd149} : s = 395;
	{8'd36,8'd150} : s = 391;
	{8'd36,8'd151} : s = 476;
	{8'd36,8'd152} : s = 376;
	{8'd36,8'd153} : s = 474;
	{8'd36,8'd154} : s = 473;
	{8'd36,8'd155} : s = 506;
	{8'd36,8'd156} : s = 20;
	{8'd36,8'd157} : s = 104;
	{8'd36,8'd158} : s = 100;
	{8'd36,8'd159} : s = 263;
	{8'd36,8'd160} : s = 98;
	{8'd36,8'd161} : s = 240;
	{8'd36,8'd162} : s = 232;
	{8'd36,8'd163} : s = 372;
	{8'd36,8'd164} : s = 97;
	{8'd36,8'd165} : s = 228;
	{8'd36,8'd166} : s = 226;
	{8'd36,8'd167} : s = 370;
	{8'd36,8'd168} : s = 225;
	{8'd36,8'd169} : s = 369;
	{8'd36,8'd170} : s = 364;
	{8'd36,8'd171} : s = 470;
	{8'd36,8'd172} : s = 88;
	{8'd36,8'd173} : s = 216;
	{8'd36,8'd174} : s = 212;
	{8'd36,8'd175} : s = 362;
	{8'd36,8'd176} : s = 210;
	{8'd36,8'd177} : s = 361;
	{8'd36,8'd178} : s = 358;
	{8'd36,8'd179} : s = 469;
	{8'd36,8'd180} : s = 209;
	{8'd36,8'd181} : s = 357;
	{8'd36,8'd182} : s = 355;
	{8'd36,8'd183} : s = 467;
	{8'd36,8'd184} : s = 348;
	{8'd36,8'd185} : s = 462;
	{8'd36,8'd186} : s = 461;
	{8'd36,8'd187} : s = 505;
	{8'd36,8'd188} : s = 84;
	{8'd36,8'd189} : s = 204;
	{8'd36,8'd190} : s = 202;
	{8'd36,8'd191} : s = 346;
	{8'd36,8'd192} : s = 201;
	{8'd36,8'd193} : s = 345;
	{8'd36,8'd194} : s = 342;
	{8'd36,8'd195} : s = 459;
	{8'd36,8'd196} : s = 198;
	{8'd36,8'd197} : s = 341;
	{8'd36,8'd198} : s = 339;
	{8'd36,8'd199} : s = 455;
	{8'd36,8'd200} : s = 334;
	{8'd36,8'd201} : s = 444;
	{8'd36,8'd202} : s = 442;
	{8'd36,8'd203} : s = 502;
	{8'd36,8'd204} : s = 197;
	{8'd36,8'd205} : s = 333;
	{8'd36,8'd206} : s = 331;
	{8'd36,8'd207} : s = 441;
	{8'd36,8'd208} : s = 327;
	{8'd36,8'd209} : s = 438;
	{8'd36,8'd210} : s = 437;
	{8'd36,8'd211} : s = 501;
	{8'd36,8'd212} : s = 316;
	{8'd36,8'd213} : s = 435;
	{8'd36,8'd214} : s = 430;
	{8'd36,8'd215} : s = 499;
	{8'd36,8'd216} : s = 429;
	{8'd36,8'd217} : s = 494;
	{8'd36,8'd218} : s = 493;
	{8'd36,8'd219} : s = 510;
	{8'd36,8'd220} : s = 1;
	{8'd36,8'd221} : s = 18;
	{8'd36,8'd222} : s = 17;
	{8'd36,8'd223} : s = 82;
	{8'd36,8'd224} : s = 12;
	{8'd36,8'd225} : s = 81;
	{8'd36,8'd226} : s = 76;
	{8'd36,8'd227} : s = 195;
	{8'd36,8'd228} : s = 10;
	{8'd36,8'd229} : s = 74;
	{8'd36,8'd230} : s = 73;
	{8'd36,8'd231} : s = 184;
	{8'd36,8'd232} : s = 70;
	{8'd36,8'd233} : s = 180;
	{8'd36,8'd234} : s = 178;
	{8'd36,8'd235} : s = 314;
	{8'd36,8'd236} : s = 9;
	{8'd36,8'd237} : s = 69;
	{8'd36,8'd238} : s = 67;
	{8'd36,8'd239} : s = 177;
	{8'd36,8'd240} : s = 56;
	{8'd36,8'd241} : s = 172;
	{8'd36,8'd242} : s = 170;
	{8'd36,8'd243} : s = 313;
	{8'd36,8'd244} : s = 52;
	{8'd36,8'd245} : s = 169;
	{8'd36,8'd246} : s = 166;
	{8'd36,8'd247} : s = 310;
	{8'd36,8'd248} : s = 165;
	{8'd36,8'd249} : s = 309;
	{8'd36,8'd250} : s = 307;
	{8'd36,8'd251} : s = 427;
	{8'd36,8'd252} : s = 6;
	{8'd36,8'd253} : s = 50;
	{8'd36,8'd254} : s = 49;
	{8'd36,8'd255} : s = 163;
	{8'd37,8'd0} : s = 322;
	{8'd37,8'd1} : s = 321;
	{8'd37,8'd2} : s = 449;
	{8'd37,8'd3} : s = 130;
	{8'd37,8'd4} : s = 304;
	{8'd37,8'd5} : s = 296;
	{8'd37,8'd6} : s = 432;
	{8'd37,8'd7} : s = 292;
	{8'd37,8'd8} : s = 424;
	{8'd37,8'd9} : s = 420;
	{8'd37,8'd10} : s = 488;
	{8'd37,8'd11} : s = 129;
	{8'd37,8'd12} : s = 290;
	{8'd37,8'd13} : s = 289;
	{8'd37,8'd14} : s = 418;
	{8'd37,8'd15} : s = 280;
	{8'd37,8'd16} : s = 417;
	{8'd37,8'd17} : s = 408;
	{8'd37,8'd18} : s = 484;
	{8'd37,8'd19} : s = 276;
	{8'd37,8'd20} : s = 404;
	{8'd37,8'd21} : s = 402;
	{8'd37,8'd22} : s = 482;
	{8'd37,8'd23} : s = 401;
	{8'd37,8'd24} : s = 481;
	{8'd37,8'd25} : s = 472;
	{8'd37,8'd26} : s = 504;
	{8'd37,8'd27} : s = 4;
	{8'd37,8'd28} : s = 96;
	{8'd37,8'd29} : s = 80;
	{8'd37,8'd30} : s = 274;
	{8'd37,8'd31} : s = 72;
	{8'd37,8'd32} : s = 273;
	{8'd37,8'd33} : s = 268;
	{8'd37,8'd34} : s = 396;
	{8'd37,8'd35} : s = 68;
	{8'd37,8'd36} : s = 266;
	{8'd37,8'd37} : s = 265;
	{8'd37,8'd38} : s = 394;
	{8'd37,8'd39} : s = 262;
	{8'd37,8'd40} : s = 393;
	{8'd37,8'd41} : s = 390;
	{8'd37,8'd42} : s = 468;
	{8'd37,8'd43} : s = 66;
	{8'd37,8'd44} : s = 261;
	{8'd37,8'd45} : s = 259;
	{8'd37,8'd46} : s = 389;
	{8'd37,8'd47} : s = 224;
	{8'd37,8'd48} : s = 387;
	{8'd37,8'd49} : s = 368;
	{8'd37,8'd50} : s = 466;
	{8'd37,8'd51} : s = 208;
	{8'd37,8'd52} : s = 360;
	{8'd37,8'd53} : s = 356;
	{8'd37,8'd54} : s = 465;
	{8'd37,8'd55} : s = 354;
	{8'd37,8'd56} : s = 460;
	{8'd37,8'd57} : s = 458;
	{8'd37,8'd58} : s = 500;
	{8'd37,8'd59} : s = 65;
	{8'd37,8'd60} : s = 200;
	{8'd37,8'd61} : s = 196;
	{8'd37,8'd62} : s = 353;
	{8'd37,8'd63} : s = 194;
	{8'd37,8'd64} : s = 344;
	{8'd37,8'd65} : s = 340;
	{8'd37,8'd66} : s = 457;
	{8'd37,8'd67} : s = 193;
	{8'd37,8'd68} : s = 338;
	{8'd37,8'd69} : s = 337;
	{8'd37,8'd70} : s = 454;
	{8'd37,8'd71} : s = 332;
	{8'd37,8'd72} : s = 453;
	{8'd37,8'd73} : s = 451;
	{8'd37,8'd74} : s = 498;
	{8'd37,8'd75} : s = 176;
	{8'd37,8'd76} : s = 330;
	{8'd37,8'd77} : s = 329;
	{8'd37,8'd78} : s = 440;
	{8'd37,8'd79} : s = 326;
	{8'd37,8'd80} : s = 436;
	{8'd37,8'd81} : s = 434;
	{8'd37,8'd82} : s = 497;
	{8'd37,8'd83} : s = 325;
	{8'd37,8'd84} : s = 433;
	{8'd37,8'd85} : s = 428;
	{8'd37,8'd86} : s = 492;
	{8'd37,8'd87} : s = 426;
	{8'd37,8'd88} : s = 490;
	{8'd37,8'd89} : s = 489;
	{8'd37,8'd90} : s = 508;
	{8'd37,8'd91} : s = 2;
	{8'd37,8'd92} : s = 48;
	{8'd37,8'd93} : s = 40;
	{8'd37,8'd94} : s = 168;
	{8'd37,8'd95} : s = 36;
	{8'd37,8'd96} : s = 164;
	{8'd37,8'd97} : s = 162;
	{8'd37,8'd98} : s = 323;
	{8'd37,8'd99} : s = 34;
	{8'd37,8'd100} : s = 161;
	{8'd37,8'd101} : s = 152;
	{8'd37,8'd102} : s = 312;
	{8'd37,8'd103} : s = 148;
	{8'd37,8'd104} : s = 308;
	{8'd37,8'd105} : s = 306;
	{8'd37,8'd106} : s = 425;
	{8'd37,8'd107} : s = 33;
	{8'd37,8'd108} : s = 146;
	{8'd37,8'd109} : s = 145;
	{8'd37,8'd110} : s = 305;
	{8'd37,8'd111} : s = 140;
	{8'd37,8'd112} : s = 300;
	{8'd37,8'd113} : s = 298;
	{8'd37,8'd114} : s = 422;
	{8'd37,8'd115} : s = 138;
	{8'd37,8'd116} : s = 297;
	{8'd37,8'd117} : s = 294;
	{8'd37,8'd118} : s = 421;
	{8'd37,8'd119} : s = 293;
	{8'd37,8'd120} : s = 419;
	{8'd37,8'd121} : s = 412;
	{8'd37,8'd122} : s = 486;
	{8'd37,8'd123} : s = 24;
	{8'd37,8'd124} : s = 137;
	{8'd37,8'd125} : s = 134;
	{8'd37,8'd126} : s = 291;
	{8'd37,8'd127} : s = 133;
	{8'd37,8'd128} : s = 284;
	{8'd37,8'd129} : s = 282;
	{8'd37,8'd130} : s = 410;
	{8'd37,8'd131} : s = 131;
	{8'd37,8'd132} : s = 281;
	{8'd37,8'd133} : s = 278;
	{8'd37,8'd134} : s = 409;
	{8'd37,8'd135} : s = 277;
	{8'd37,8'd136} : s = 406;
	{8'd37,8'd137} : s = 405;
	{8'd37,8'd138} : s = 485;
	{8'd37,8'd139} : s = 112;
	{8'd37,8'd140} : s = 275;
	{8'd37,8'd141} : s = 270;
	{8'd37,8'd142} : s = 403;
	{8'd37,8'd143} : s = 269;
	{8'd37,8'd144} : s = 398;
	{8'd37,8'd145} : s = 397;
	{8'd37,8'd146} : s = 483;
	{8'd37,8'd147} : s = 267;
	{8'd37,8'd148} : s = 395;
	{8'd37,8'd149} : s = 391;
	{8'd37,8'd150} : s = 476;
	{8'd37,8'd151} : s = 376;
	{8'd37,8'd152} : s = 474;
	{8'd37,8'd153} : s = 473;
	{8'd37,8'd154} : s = 506;
	{8'd37,8'd155} : s = 20;
	{8'd37,8'd156} : s = 104;
	{8'd37,8'd157} : s = 100;
	{8'd37,8'd158} : s = 263;
	{8'd37,8'd159} : s = 98;
	{8'd37,8'd160} : s = 240;
	{8'd37,8'd161} : s = 232;
	{8'd37,8'd162} : s = 372;
	{8'd37,8'd163} : s = 97;
	{8'd37,8'd164} : s = 228;
	{8'd37,8'd165} : s = 226;
	{8'd37,8'd166} : s = 370;
	{8'd37,8'd167} : s = 225;
	{8'd37,8'd168} : s = 369;
	{8'd37,8'd169} : s = 364;
	{8'd37,8'd170} : s = 470;
	{8'd37,8'd171} : s = 88;
	{8'd37,8'd172} : s = 216;
	{8'd37,8'd173} : s = 212;
	{8'd37,8'd174} : s = 362;
	{8'd37,8'd175} : s = 210;
	{8'd37,8'd176} : s = 361;
	{8'd37,8'd177} : s = 358;
	{8'd37,8'd178} : s = 469;
	{8'd37,8'd179} : s = 209;
	{8'd37,8'd180} : s = 357;
	{8'd37,8'd181} : s = 355;
	{8'd37,8'd182} : s = 467;
	{8'd37,8'd183} : s = 348;
	{8'd37,8'd184} : s = 462;
	{8'd37,8'd185} : s = 461;
	{8'd37,8'd186} : s = 505;
	{8'd37,8'd187} : s = 84;
	{8'd37,8'd188} : s = 204;
	{8'd37,8'd189} : s = 202;
	{8'd37,8'd190} : s = 346;
	{8'd37,8'd191} : s = 201;
	{8'd37,8'd192} : s = 345;
	{8'd37,8'd193} : s = 342;
	{8'd37,8'd194} : s = 459;
	{8'd37,8'd195} : s = 198;
	{8'd37,8'd196} : s = 341;
	{8'd37,8'd197} : s = 339;
	{8'd37,8'd198} : s = 455;
	{8'd37,8'd199} : s = 334;
	{8'd37,8'd200} : s = 444;
	{8'd37,8'd201} : s = 442;
	{8'd37,8'd202} : s = 502;
	{8'd37,8'd203} : s = 197;
	{8'd37,8'd204} : s = 333;
	{8'd37,8'd205} : s = 331;
	{8'd37,8'd206} : s = 441;
	{8'd37,8'd207} : s = 327;
	{8'd37,8'd208} : s = 438;
	{8'd37,8'd209} : s = 437;
	{8'd37,8'd210} : s = 501;
	{8'd37,8'd211} : s = 316;
	{8'd37,8'd212} : s = 435;
	{8'd37,8'd213} : s = 430;
	{8'd37,8'd214} : s = 499;
	{8'd37,8'd215} : s = 429;
	{8'd37,8'd216} : s = 494;
	{8'd37,8'd217} : s = 493;
	{8'd37,8'd218} : s = 510;
	{8'd37,8'd219} : s = 1;
	{8'd37,8'd220} : s = 18;
	{8'd37,8'd221} : s = 17;
	{8'd37,8'd222} : s = 82;
	{8'd37,8'd223} : s = 12;
	{8'd37,8'd224} : s = 81;
	{8'd37,8'd225} : s = 76;
	{8'd37,8'd226} : s = 195;
	{8'd37,8'd227} : s = 10;
	{8'd37,8'd228} : s = 74;
	{8'd37,8'd229} : s = 73;
	{8'd37,8'd230} : s = 184;
	{8'd37,8'd231} : s = 70;
	{8'd37,8'd232} : s = 180;
	{8'd37,8'd233} : s = 178;
	{8'd37,8'd234} : s = 314;
	{8'd37,8'd235} : s = 9;
	{8'd37,8'd236} : s = 69;
	{8'd37,8'd237} : s = 67;
	{8'd37,8'd238} : s = 177;
	{8'd37,8'd239} : s = 56;
	{8'd37,8'd240} : s = 172;
	{8'd37,8'd241} : s = 170;
	{8'd37,8'd242} : s = 313;
	{8'd37,8'd243} : s = 52;
	{8'd37,8'd244} : s = 169;
	{8'd37,8'd245} : s = 166;
	{8'd37,8'd246} : s = 310;
	{8'd37,8'd247} : s = 165;
	{8'd37,8'd248} : s = 309;
	{8'd37,8'd249} : s = 307;
	{8'd37,8'd250} : s = 427;
	{8'd37,8'd251} : s = 6;
	{8'd37,8'd252} : s = 50;
	{8'd37,8'd253} : s = 49;
	{8'd37,8'd254} : s = 163;
	{8'd37,8'd255} : s = 44;
	{8'd38,8'd0} : s = 321;
	{8'd38,8'd1} : s = 449;
	{8'd38,8'd2} : s = 130;
	{8'd38,8'd3} : s = 304;
	{8'd38,8'd4} : s = 296;
	{8'd38,8'd5} : s = 432;
	{8'd38,8'd6} : s = 292;
	{8'd38,8'd7} : s = 424;
	{8'd38,8'd8} : s = 420;
	{8'd38,8'd9} : s = 488;
	{8'd38,8'd10} : s = 129;
	{8'd38,8'd11} : s = 290;
	{8'd38,8'd12} : s = 289;
	{8'd38,8'd13} : s = 418;
	{8'd38,8'd14} : s = 280;
	{8'd38,8'd15} : s = 417;
	{8'd38,8'd16} : s = 408;
	{8'd38,8'd17} : s = 484;
	{8'd38,8'd18} : s = 276;
	{8'd38,8'd19} : s = 404;
	{8'd38,8'd20} : s = 402;
	{8'd38,8'd21} : s = 482;
	{8'd38,8'd22} : s = 401;
	{8'd38,8'd23} : s = 481;
	{8'd38,8'd24} : s = 472;
	{8'd38,8'd25} : s = 504;
	{8'd38,8'd26} : s = 4;
	{8'd38,8'd27} : s = 96;
	{8'd38,8'd28} : s = 80;
	{8'd38,8'd29} : s = 274;
	{8'd38,8'd30} : s = 72;
	{8'd38,8'd31} : s = 273;
	{8'd38,8'd32} : s = 268;
	{8'd38,8'd33} : s = 396;
	{8'd38,8'd34} : s = 68;
	{8'd38,8'd35} : s = 266;
	{8'd38,8'd36} : s = 265;
	{8'd38,8'd37} : s = 394;
	{8'd38,8'd38} : s = 262;
	{8'd38,8'd39} : s = 393;
	{8'd38,8'd40} : s = 390;
	{8'd38,8'd41} : s = 468;
	{8'd38,8'd42} : s = 66;
	{8'd38,8'd43} : s = 261;
	{8'd38,8'd44} : s = 259;
	{8'd38,8'd45} : s = 389;
	{8'd38,8'd46} : s = 224;
	{8'd38,8'd47} : s = 387;
	{8'd38,8'd48} : s = 368;
	{8'd38,8'd49} : s = 466;
	{8'd38,8'd50} : s = 208;
	{8'd38,8'd51} : s = 360;
	{8'd38,8'd52} : s = 356;
	{8'd38,8'd53} : s = 465;
	{8'd38,8'd54} : s = 354;
	{8'd38,8'd55} : s = 460;
	{8'd38,8'd56} : s = 458;
	{8'd38,8'd57} : s = 500;
	{8'd38,8'd58} : s = 65;
	{8'd38,8'd59} : s = 200;
	{8'd38,8'd60} : s = 196;
	{8'd38,8'd61} : s = 353;
	{8'd38,8'd62} : s = 194;
	{8'd38,8'd63} : s = 344;
	{8'd38,8'd64} : s = 340;
	{8'd38,8'd65} : s = 457;
	{8'd38,8'd66} : s = 193;
	{8'd38,8'd67} : s = 338;
	{8'd38,8'd68} : s = 337;
	{8'd38,8'd69} : s = 454;
	{8'd38,8'd70} : s = 332;
	{8'd38,8'd71} : s = 453;
	{8'd38,8'd72} : s = 451;
	{8'd38,8'd73} : s = 498;
	{8'd38,8'd74} : s = 176;
	{8'd38,8'd75} : s = 330;
	{8'd38,8'd76} : s = 329;
	{8'd38,8'd77} : s = 440;
	{8'd38,8'd78} : s = 326;
	{8'd38,8'd79} : s = 436;
	{8'd38,8'd80} : s = 434;
	{8'd38,8'd81} : s = 497;
	{8'd38,8'd82} : s = 325;
	{8'd38,8'd83} : s = 433;
	{8'd38,8'd84} : s = 428;
	{8'd38,8'd85} : s = 492;
	{8'd38,8'd86} : s = 426;
	{8'd38,8'd87} : s = 490;
	{8'd38,8'd88} : s = 489;
	{8'd38,8'd89} : s = 508;
	{8'd38,8'd90} : s = 2;
	{8'd38,8'd91} : s = 48;
	{8'd38,8'd92} : s = 40;
	{8'd38,8'd93} : s = 168;
	{8'd38,8'd94} : s = 36;
	{8'd38,8'd95} : s = 164;
	{8'd38,8'd96} : s = 162;
	{8'd38,8'd97} : s = 323;
	{8'd38,8'd98} : s = 34;
	{8'd38,8'd99} : s = 161;
	{8'd38,8'd100} : s = 152;
	{8'd38,8'd101} : s = 312;
	{8'd38,8'd102} : s = 148;
	{8'd38,8'd103} : s = 308;
	{8'd38,8'd104} : s = 306;
	{8'd38,8'd105} : s = 425;
	{8'd38,8'd106} : s = 33;
	{8'd38,8'd107} : s = 146;
	{8'd38,8'd108} : s = 145;
	{8'd38,8'd109} : s = 305;
	{8'd38,8'd110} : s = 140;
	{8'd38,8'd111} : s = 300;
	{8'd38,8'd112} : s = 298;
	{8'd38,8'd113} : s = 422;
	{8'd38,8'd114} : s = 138;
	{8'd38,8'd115} : s = 297;
	{8'd38,8'd116} : s = 294;
	{8'd38,8'd117} : s = 421;
	{8'd38,8'd118} : s = 293;
	{8'd38,8'd119} : s = 419;
	{8'd38,8'd120} : s = 412;
	{8'd38,8'd121} : s = 486;
	{8'd38,8'd122} : s = 24;
	{8'd38,8'd123} : s = 137;
	{8'd38,8'd124} : s = 134;
	{8'd38,8'd125} : s = 291;
	{8'd38,8'd126} : s = 133;
	{8'd38,8'd127} : s = 284;
	{8'd38,8'd128} : s = 282;
	{8'd38,8'd129} : s = 410;
	{8'd38,8'd130} : s = 131;
	{8'd38,8'd131} : s = 281;
	{8'd38,8'd132} : s = 278;
	{8'd38,8'd133} : s = 409;
	{8'd38,8'd134} : s = 277;
	{8'd38,8'd135} : s = 406;
	{8'd38,8'd136} : s = 405;
	{8'd38,8'd137} : s = 485;
	{8'd38,8'd138} : s = 112;
	{8'd38,8'd139} : s = 275;
	{8'd38,8'd140} : s = 270;
	{8'd38,8'd141} : s = 403;
	{8'd38,8'd142} : s = 269;
	{8'd38,8'd143} : s = 398;
	{8'd38,8'd144} : s = 397;
	{8'd38,8'd145} : s = 483;
	{8'd38,8'd146} : s = 267;
	{8'd38,8'd147} : s = 395;
	{8'd38,8'd148} : s = 391;
	{8'd38,8'd149} : s = 476;
	{8'd38,8'd150} : s = 376;
	{8'd38,8'd151} : s = 474;
	{8'd38,8'd152} : s = 473;
	{8'd38,8'd153} : s = 506;
	{8'd38,8'd154} : s = 20;
	{8'd38,8'd155} : s = 104;
	{8'd38,8'd156} : s = 100;
	{8'd38,8'd157} : s = 263;
	{8'd38,8'd158} : s = 98;
	{8'd38,8'd159} : s = 240;
	{8'd38,8'd160} : s = 232;
	{8'd38,8'd161} : s = 372;
	{8'd38,8'd162} : s = 97;
	{8'd38,8'd163} : s = 228;
	{8'd38,8'd164} : s = 226;
	{8'd38,8'd165} : s = 370;
	{8'd38,8'd166} : s = 225;
	{8'd38,8'd167} : s = 369;
	{8'd38,8'd168} : s = 364;
	{8'd38,8'd169} : s = 470;
	{8'd38,8'd170} : s = 88;
	{8'd38,8'd171} : s = 216;
	{8'd38,8'd172} : s = 212;
	{8'd38,8'd173} : s = 362;
	{8'd38,8'd174} : s = 210;
	{8'd38,8'd175} : s = 361;
	{8'd38,8'd176} : s = 358;
	{8'd38,8'd177} : s = 469;
	{8'd38,8'd178} : s = 209;
	{8'd38,8'd179} : s = 357;
	{8'd38,8'd180} : s = 355;
	{8'd38,8'd181} : s = 467;
	{8'd38,8'd182} : s = 348;
	{8'd38,8'd183} : s = 462;
	{8'd38,8'd184} : s = 461;
	{8'd38,8'd185} : s = 505;
	{8'd38,8'd186} : s = 84;
	{8'd38,8'd187} : s = 204;
	{8'd38,8'd188} : s = 202;
	{8'd38,8'd189} : s = 346;
	{8'd38,8'd190} : s = 201;
	{8'd38,8'd191} : s = 345;
	{8'd38,8'd192} : s = 342;
	{8'd38,8'd193} : s = 459;
	{8'd38,8'd194} : s = 198;
	{8'd38,8'd195} : s = 341;
	{8'd38,8'd196} : s = 339;
	{8'd38,8'd197} : s = 455;
	{8'd38,8'd198} : s = 334;
	{8'd38,8'd199} : s = 444;
	{8'd38,8'd200} : s = 442;
	{8'd38,8'd201} : s = 502;
	{8'd38,8'd202} : s = 197;
	{8'd38,8'd203} : s = 333;
	{8'd38,8'd204} : s = 331;
	{8'd38,8'd205} : s = 441;
	{8'd38,8'd206} : s = 327;
	{8'd38,8'd207} : s = 438;
	{8'd38,8'd208} : s = 437;
	{8'd38,8'd209} : s = 501;
	{8'd38,8'd210} : s = 316;
	{8'd38,8'd211} : s = 435;
	{8'd38,8'd212} : s = 430;
	{8'd38,8'd213} : s = 499;
	{8'd38,8'd214} : s = 429;
	{8'd38,8'd215} : s = 494;
	{8'd38,8'd216} : s = 493;
	{8'd38,8'd217} : s = 510;
	{8'd38,8'd218} : s = 1;
	{8'd38,8'd219} : s = 18;
	{8'd38,8'd220} : s = 17;
	{8'd38,8'd221} : s = 82;
	{8'd38,8'd222} : s = 12;
	{8'd38,8'd223} : s = 81;
	{8'd38,8'd224} : s = 76;
	{8'd38,8'd225} : s = 195;
	{8'd38,8'd226} : s = 10;
	{8'd38,8'd227} : s = 74;
	{8'd38,8'd228} : s = 73;
	{8'd38,8'd229} : s = 184;
	{8'd38,8'd230} : s = 70;
	{8'd38,8'd231} : s = 180;
	{8'd38,8'd232} : s = 178;
	{8'd38,8'd233} : s = 314;
	{8'd38,8'd234} : s = 9;
	{8'd38,8'd235} : s = 69;
	{8'd38,8'd236} : s = 67;
	{8'd38,8'd237} : s = 177;
	{8'd38,8'd238} : s = 56;
	{8'd38,8'd239} : s = 172;
	{8'd38,8'd240} : s = 170;
	{8'd38,8'd241} : s = 313;
	{8'd38,8'd242} : s = 52;
	{8'd38,8'd243} : s = 169;
	{8'd38,8'd244} : s = 166;
	{8'd38,8'd245} : s = 310;
	{8'd38,8'd246} : s = 165;
	{8'd38,8'd247} : s = 309;
	{8'd38,8'd248} : s = 307;
	{8'd38,8'd249} : s = 427;
	{8'd38,8'd250} : s = 6;
	{8'd38,8'd251} : s = 50;
	{8'd38,8'd252} : s = 49;
	{8'd38,8'd253} : s = 163;
	{8'd38,8'd254} : s = 44;
	{8'd38,8'd255} : s = 156;
	{8'd39,8'd0} : s = 449;
	{8'd39,8'd1} : s = 130;
	{8'd39,8'd2} : s = 304;
	{8'd39,8'd3} : s = 296;
	{8'd39,8'd4} : s = 432;
	{8'd39,8'd5} : s = 292;
	{8'd39,8'd6} : s = 424;
	{8'd39,8'd7} : s = 420;
	{8'd39,8'd8} : s = 488;
	{8'd39,8'd9} : s = 129;
	{8'd39,8'd10} : s = 290;
	{8'd39,8'd11} : s = 289;
	{8'd39,8'd12} : s = 418;
	{8'd39,8'd13} : s = 280;
	{8'd39,8'd14} : s = 417;
	{8'd39,8'd15} : s = 408;
	{8'd39,8'd16} : s = 484;
	{8'd39,8'd17} : s = 276;
	{8'd39,8'd18} : s = 404;
	{8'd39,8'd19} : s = 402;
	{8'd39,8'd20} : s = 482;
	{8'd39,8'd21} : s = 401;
	{8'd39,8'd22} : s = 481;
	{8'd39,8'd23} : s = 472;
	{8'd39,8'd24} : s = 504;
	{8'd39,8'd25} : s = 4;
	{8'd39,8'd26} : s = 96;
	{8'd39,8'd27} : s = 80;
	{8'd39,8'd28} : s = 274;
	{8'd39,8'd29} : s = 72;
	{8'd39,8'd30} : s = 273;
	{8'd39,8'd31} : s = 268;
	{8'd39,8'd32} : s = 396;
	{8'd39,8'd33} : s = 68;
	{8'd39,8'd34} : s = 266;
	{8'd39,8'd35} : s = 265;
	{8'd39,8'd36} : s = 394;
	{8'd39,8'd37} : s = 262;
	{8'd39,8'd38} : s = 393;
	{8'd39,8'd39} : s = 390;
	{8'd39,8'd40} : s = 468;
	{8'd39,8'd41} : s = 66;
	{8'd39,8'd42} : s = 261;
	{8'd39,8'd43} : s = 259;
	{8'd39,8'd44} : s = 389;
	{8'd39,8'd45} : s = 224;
	{8'd39,8'd46} : s = 387;
	{8'd39,8'd47} : s = 368;
	{8'd39,8'd48} : s = 466;
	{8'd39,8'd49} : s = 208;
	{8'd39,8'd50} : s = 360;
	{8'd39,8'd51} : s = 356;
	{8'd39,8'd52} : s = 465;
	{8'd39,8'd53} : s = 354;
	{8'd39,8'd54} : s = 460;
	{8'd39,8'd55} : s = 458;
	{8'd39,8'd56} : s = 500;
	{8'd39,8'd57} : s = 65;
	{8'd39,8'd58} : s = 200;
	{8'd39,8'd59} : s = 196;
	{8'd39,8'd60} : s = 353;
	{8'd39,8'd61} : s = 194;
	{8'd39,8'd62} : s = 344;
	{8'd39,8'd63} : s = 340;
	{8'd39,8'd64} : s = 457;
	{8'd39,8'd65} : s = 193;
	{8'd39,8'd66} : s = 338;
	{8'd39,8'd67} : s = 337;
	{8'd39,8'd68} : s = 454;
	{8'd39,8'd69} : s = 332;
	{8'd39,8'd70} : s = 453;
	{8'd39,8'd71} : s = 451;
	{8'd39,8'd72} : s = 498;
	{8'd39,8'd73} : s = 176;
	{8'd39,8'd74} : s = 330;
	{8'd39,8'd75} : s = 329;
	{8'd39,8'd76} : s = 440;
	{8'd39,8'd77} : s = 326;
	{8'd39,8'd78} : s = 436;
	{8'd39,8'd79} : s = 434;
	{8'd39,8'd80} : s = 497;
	{8'd39,8'd81} : s = 325;
	{8'd39,8'd82} : s = 433;
	{8'd39,8'd83} : s = 428;
	{8'd39,8'd84} : s = 492;
	{8'd39,8'd85} : s = 426;
	{8'd39,8'd86} : s = 490;
	{8'd39,8'd87} : s = 489;
	{8'd39,8'd88} : s = 508;
	{8'd39,8'd89} : s = 2;
	{8'd39,8'd90} : s = 48;
	{8'd39,8'd91} : s = 40;
	{8'd39,8'd92} : s = 168;
	{8'd39,8'd93} : s = 36;
	{8'd39,8'd94} : s = 164;
	{8'd39,8'd95} : s = 162;
	{8'd39,8'd96} : s = 323;
	{8'd39,8'd97} : s = 34;
	{8'd39,8'd98} : s = 161;
	{8'd39,8'd99} : s = 152;
	{8'd39,8'd100} : s = 312;
	{8'd39,8'd101} : s = 148;
	{8'd39,8'd102} : s = 308;
	{8'd39,8'd103} : s = 306;
	{8'd39,8'd104} : s = 425;
	{8'd39,8'd105} : s = 33;
	{8'd39,8'd106} : s = 146;
	{8'd39,8'd107} : s = 145;
	{8'd39,8'd108} : s = 305;
	{8'd39,8'd109} : s = 140;
	{8'd39,8'd110} : s = 300;
	{8'd39,8'd111} : s = 298;
	{8'd39,8'd112} : s = 422;
	{8'd39,8'd113} : s = 138;
	{8'd39,8'd114} : s = 297;
	{8'd39,8'd115} : s = 294;
	{8'd39,8'd116} : s = 421;
	{8'd39,8'd117} : s = 293;
	{8'd39,8'd118} : s = 419;
	{8'd39,8'd119} : s = 412;
	{8'd39,8'd120} : s = 486;
	{8'd39,8'd121} : s = 24;
	{8'd39,8'd122} : s = 137;
	{8'd39,8'd123} : s = 134;
	{8'd39,8'd124} : s = 291;
	{8'd39,8'd125} : s = 133;
	{8'd39,8'd126} : s = 284;
	{8'd39,8'd127} : s = 282;
	{8'd39,8'd128} : s = 410;
	{8'd39,8'd129} : s = 131;
	{8'd39,8'd130} : s = 281;
	{8'd39,8'd131} : s = 278;
	{8'd39,8'd132} : s = 409;
	{8'd39,8'd133} : s = 277;
	{8'd39,8'd134} : s = 406;
	{8'd39,8'd135} : s = 405;
	{8'd39,8'd136} : s = 485;
	{8'd39,8'd137} : s = 112;
	{8'd39,8'd138} : s = 275;
	{8'd39,8'd139} : s = 270;
	{8'd39,8'd140} : s = 403;
	{8'd39,8'd141} : s = 269;
	{8'd39,8'd142} : s = 398;
	{8'd39,8'd143} : s = 397;
	{8'd39,8'd144} : s = 483;
	{8'd39,8'd145} : s = 267;
	{8'd39,8'd146} : s = 395;
	{8'd39,8'd147} : s = 391;
	{8'd39,8'd148} : s = 476;
	{8'd39,8'd149} : s = 376;
	{8'd39,8'd150} : s = 474;
	{8'd39,8'd151} : s = 473;
	{8'd39,8'd152} : s = 506;
	{8'd39,8'd153} : s = 20;
	{8'd39,8'd154} : s = 104;
	{8'd39,8'd155} : s = 100;
	{8'd39,8'd156} : s = 263;
	{8'd39,8'd157} : s = 98;
	{8'd39,8'd158} : s = 240;
	{8'd39,8'd159} : s = 232;
	{8'd39,8'd160} : s = 372;
	{8'd39,8'd161} : s = 97;
	{8'd39,8'd162} : s = 228;
	{8'd39,8'd163} : s = 226;
	{8'd39,8'd164} : s = 370;
	{8'd39,8'd165} : s = 225;
	{8'd39,8'd166} : s = 369;
	{8'd39,8'd167} : s = 364;
	{8'd39,8'd168} : s = 470;
	{8'd39,8'd169} : s = 88;
	{8'd39,8'd170} : s = 216;
	{8'd39,8'd171} : s = 212;
	{8'd39,8'd172} : s = 362;
	{8'd39,8'd173} : s = 210;
	{8'd39,8'd174} : s = 361;
	{8'd39,8'd175} : s = 358;
	{8'd39,8'd176} : s = 469;
	{8'd39,8'd177} : s = 209;
	{8'd39,8'd178} : s = 357;
	{8'd39,8'd179} : s = 355;
	{8'd39,8'd180} : s = 467;
	{8'd39,8'd181} : s = 348;
	{8'd39,8'd182} : s = 462;
	{8'd39,8'd183} : s = 461;
	{8'd39,8'd184} : s = 505;
	{8'd39,8'd185} : s = 84;
	{8'd39,8'd186} : s = 204;
	{8'd39,8'd187} : s = 202;
	{8'd39,8'd188} : s = 346;
	{8'd39,8'd189} : s = 201;
	{8'd39,8'd190} : s = 345;
	{8'd39,8'd191} : s = 342;
	{8'd39,8'd192} : s = 459;
	{8'd39,8'd193} : s = 198;
	{8'd39,8'd194} : s = 341;
	{8'd39,8'd195} : s = 339;
	{8'd39,8'd196} : s = 455;
	{8'd39,8'd197} : s = 334;
	{8'd39,8'd198} : s = 444;
	{8'd39,8'd199} : s = 442;
	{8'd39,8'd200} : s = 502;
	{8'd39,8'd201} : s = 197;
	{8'd39,8'd202} : s = 333;
	{8'd39,8'd203} : s = 331;
	{8'd39,8'd204} : s = 441;
	{8'd39,8'd205} : s = 327;
	{8'd39,8'd206} : s = 438;
	{8'd39,8'd207} : s = 437;
	{8'd39,8'd208} : s = 501;
	{8'd39,8'd209} : s = 316;
	{8'd39,8'd210} : s = 435;
	{8'd39,8'd211} : s = 430;
	{8'd39,8'd212} : s = 499;
	{8'd39,8'd213} : s = 429;
	{8'd39,8'd214} : s = 494;
	{8'd39,8'd215} : s = 493;
	{8'd39,8'd216} : s = 510;
	{8'd39,8'd217} : s = 1;
	{8'd39,8'd218} : s = 18;
	{8'd39,8'd219} : s = 17;
	{8'd39,8'd220} : s = 82;
	{8'd39,8'd221} : s = 12;
	{8'd39,8'd222} : s = 81;
	{8'd39,8'd223} : s = 76;
	{8'd39,8'd224} : s = 195;
	{8'd39,8'd225} : s = 10;
	{8'd39,8'd226} : s = 74;
	{8'd39,8'd227} : s = 73;
	{8'd39,8'd228} : s = 184;
	{8'd39,8'd229} : s = 70;
	{8'd39,8'd230} : s = 180;
	{8'd39,8'd231} : s = 178;
	{8'd39,8'd232} : s = 314;
	{8'd39,8'd233} : s = 9;
	{8'd39,8'd234} : s = 69;
	{8'd39,8'd235} : s = 67;
	{8'd39,8'd236} : s = 177;
	{8'd39,8'd237} : s = 56;
	{8'd39,8'd238} : s = 172;
	{8'd39,8'd239} : s = 170;
	{8'd39,8'd240} : s = 313;
	{8'd39,8'd241} : s = 52;
	{8'd39,8'd242} : s = 169;
	{8'd39,8'd243} : s = 166;
	{8'd39,8'd244} : s = 310;
	{8'd39,8'd245} : s = 165;
	{8'd39,8'd246} : s = 309;
	{8'd39,8'd247} : s = 307;
	{8'd39,8'd248} : s = 427;
	{8'd39,8'd249} : s = 6;
	{8'd39,8'd250} : s = 50;
	{8'd39,8'd251} : s = 49;
	{8'd39,8'd252} : s = 163;
	{8'd39,8'd253} : s = 44;
	{8'd39,8'd254} : s = 156;
	{8'd39,8'd255} : s = 154;
	{8'd40,8'd0} : s = 130;
	{8'd40,8'd1} : s = 304;
	{8'd40,8'd2} : s = 296;
	{8'd40,8'd3} : s = 432;
	{8'd40,8'd4} : s = 292;
	{8'd40,8'd5} : s = 424;
	{8'd40,8'd6} : s = 420;
	{8'd40,8'd7} : s = 488;
	{8'd40,8'd8} : s = 129;
	{8'd40,8'd9} : s = 290;
	{8'd40,8'd10} : s = 289;
	{8'd40,8'd11} : s = 418;
	{8'd40,8'd12} : s = 280;
	{8'd40,8'd13} : s = 417;
	{8'd40,8'd14} : s = 408;
	{8'd40,8'd15} : s = 484;
	{8'd40,8'd16} : s = 276;
	{8'd40,8'd17} : s = 404;
	{8'd40,8'd18} : s = 402;
	{8'd40,8'd19} : s = 482;
	{8'd40,8'd20} : s = 401;
	{8'd40,8'd21} : s = 481;
	{8'd40,8'd22} : s = 472;
	{8'd40,8'd23} : s = 504;
	{8'd40,8'd24} : s = 4;
	{8'd40,8'd25} : s = 96;
	{8'd40,8'd26} : s = 80;
	{8'd40,8'd27} : s = 274;
	{8'd40,8'd28} : s = 72;
	{8'd40,8'd29} : s = 273;
	{8'd40,8'd30} : s = 268;
	{8'd40,8'd31} : s = 396;
	{8'd40,8'd32} : s = 68;
	{8'd40,8'd33} : s = 266;
	{8'd40,8'd34} : s = 265;
	{8'd40,8'd35} : s = 394;
	{8'd40,8'd36} : s = 262;
	{8'd40,8'd37} : s = 393;
	{8'd40,8'd38} : s = 390;
	{8'd40,8'd39} : s = 468;
	{8'd40,8'd40} : s = 66;
	{8'd40,8'd41} : s = 261;
	{8'd40,8'd42} : s = 259;
	{8'd40,8'd43} : s = 389;
	{8'd40,8'd44} : s = 224;
	{8'd40,8'd45} : s = 387;
	{8'd40,8'd46} : s = 368;
	{8'd40,8'd47} : s = 466;
	{8'd40,8'd48} : s = 208;
	{8'd40,8'd49} : s = 360;
	{8'd40,8'd50} : s = 356;
	{8'd40,8'd51} : s = 465;
	{8'd40,8'd52} : s = 354;
	{8'd40,8'd53} : s = 460;
	{8'd40,8'd54} : s = 458;
	{8'd40,8'd55} : s = 500;
	{8'd40,8'd56} : s = 65;
	{8'd40,8'd57} : s = 200;
	{8'd40,8'd58} : s = 196;
	{8'd40,8'd59} : s = 353;
	{8'd40,8'd60} : s = 194;
	{8'd40,8'd61} : s = 344;
	{8'd40,8'd62} : s = 340;
	{8'd40,8'd63} : s = 457;
	{8'd40,8'd64} : s = 193;
	{8'd40,8'd65} : s = 338;
	{8'd40,8'd66} : s = 337;
	{8'd40,8'd67} : s = 454;
	{8'd40,8'd68} : s = 332;
	{8'd40,8'd69} : s = 453;
	{8'd40,8'd70} : s = 451;
	{8'd40,8'd71} : s = 498;
	{8'd40,8'd72} : s = 176;
	{8'd40,8'd73} : s = 330;
	{8'd40,8'd74} : s = 329;
	{8'd40,8'd75} : s = 440;
	{8'd40,8'd76} : s = 326;
	{8'd40,8'd77} : s = 436;
	{8'd40,8'd78} : s = 434;
	{8'd40,8'd79} : s = 497;
	{8'd40,8'd80} : s = 325;
	{8'd40,8'd81} : s = 433;
	{8'd40,8'd82} : s = 428;
	{8'd40,8'd83} : s = 492;
	{8'd40,8'd84} : s = 426;
	{8'd40,8'd85} : s = 490;
	{8'd40,8'd86} : s = 489;
	{8'd40,8'd87} : s = 508;
	{8'd40,8'd88} : s = 2;
	{8'd40,8'd89} : s = 48;
	{8'd40,8'd90} : s = 40;
	{8'd40,8'd91} : s = 168;
	{8'd40,8'd92} : s = 36;
	{8'd40,8'd93} : s = 164;
	{8'd40,8'd94} : s = 162;
	{8'd40,8'd95} : s = 323;
	{8'd40,8'd96} : s = 34;
	{8'd40,8'd97} : s = 161;
	{8'd40,8'd98} : s = 152;
	{8'd40,8'd99} : s = 312;
	{8'd40,8'd100} : s = 148;
	{8'd40,8'd101} : s = 308;
	{8'd40,8'd102} : s = 306;
	{8'd40,8'd103} : s = 425;
	{8'd40,8'd104} : s = 33;
	{8'd40,8'd105} : s = 146;
	{8'd40,8'd106} : s = 145;
	{8'd40,8'd107} : s = 305;
	{8'd40,8'd108} : s = 140;
	{8'd40,8'd109} : s = 300;
	{8'd40,8'd110} : s = 298;
	{8'd40,8'd111} : s = 422;
	{8'd40,8'd112} : s = 138;
	{8'd40,8'd113} : s = 297;
	{8'd40,8'd114} : s = 294;
	{8'd40,8'd115} : s = 421;
	{8'd40,8'd116} : s = 293;
	{8'd40,8'd117} : s = 419;
	{8'd40,8'd118} : s = 412;
	{8'd40,8'd119} : s = 486;
	{8'd40,8'd120} : s = 24;
	{8'd40,8'd121} : s = 137;
	{8'd40,8'd122} : s = 134;
	{8'd40,8'd123} : s = 291;
	{8'd40,8'd124} : s = 133;
	{8'd40,8'd125} : s = 284;
	{8'd40,8'd126} : s = 282;
	{8'd40,8'd127} : s = 410;
	{8'd40,8'd128} : s = 131;
	{8'd40,8'd129} : s = 281;
	{8'd40,8'd130} : s = 278;
	{8'd40,8'd131} : s = 409;
	{8'd40,8'd132} : s = 277;
	{8'd40,8'd133} : s = 406;
	{8'd40,8'd134} : s = 405;
	{8'd40,8'd135} : s = 485;
	{8'd40,8'd136} : s = 112;
	{8'd40,8'd137} : s = 275;
	{8'd40,8'd138} : s = 270;
	{8'd40,8'd139} : s = 403;
	{8'd40,8'd140} : s = 269;
	{8'd40,8'd141} : s = 398;
	{8'd40,8'd142} : s = 397;
	{8'd40,8'd143} : s = 483;
	{8'd40,8'd144} : s = 267;
	{8'd40,8'd145} : s = 395;
	{8'd40,8'd146} : s = 391;
	{8'd40,8'd147} : s = 476;
	{8'd40,8'd148} : s = 376;
	{8'd40,8'd149} : s = 474;
	{8'd40,8'd150} : s = 473;
	{8'd40,8'd151} : s = 506;
	{8'd40,8'd152} : s = 20;
	{8'd40,8'd153} : s = 104;
	{8'd40,8'd154} : s = 100;
	{8'd40,8'd155} : s = 263;
	{8'd40,8'd156} : s = 98;
	{8'd40,8'd157} : s = 240;
	{8'd40,8'd158} : s = 232;
	{8'd40,8'd159} : s = 372;
	{8'd40,8'd160} : s = 97;
	{8'd40,8'd161} : s = 228;
	{8'd40,8'd162} : s = 226;
	{8'd40,8'd163} : s = 370;
	{8'd40,8'd164} : s = 225;
	{8'd40,8'd165} : s = 369;
	{8'd40,8'd166} : s = 364;
	{8'd40,8'd167} : s = 470;
	{8'd40,8'd168} : s = 88;
	{8'd40,8'd169} : s = 216;
	{8'd40,8'd170} : s = 212;
	{8'd40,8'd171} : s = 362;
	{8'd40,8'd172} : s = 210;
	{8'd40,8'd173} : s = 361;
	{8'd40,8'd174} : s = 358;
	{8'd40,8'd175} : s = 469;
	{8'd40,8'd176} : s = 209;
	{8'd40,8'd177} : s = 357;
	{8'd40,8'd178} : s = 355;
	{8'd40,8'd179} : s = 467;
	{8'd40,8'd180} : s = 348;
	{8'd40,8'd181} : s = 462;
	{8'd40,8'd182} : s = 461;
	{8'd40,8'd183} : s = 505;
	{8'd40,8'd184} : s = 84;
	{8'd40,8'd185} : s = 204;
	{8'd40,8'd186} : s = 202;
	{8'd40,8'd187} : s = 346;
	{8'd40,8'd188} : s = 201;
	{8'd40,8'd189} : s = 345;
	{8'd40,8'd190} : s = 342;
	{8'd40,8'd191} : s = 459;
	{8'd40,8'd192} : s = 198;
	{8'd40,8'd193} : s = 341;
	{8'd40,8'd194} : s = 339;
	{8'd40,8'd195} : s = 455;
	{8'd40,8'd196} : s = 334;
	{8'd40,8'd197} : s = 444;
	{8'd40,8'd198} : s = 442;
	{8'd40,8'd199} : s = 502;
	{8'd40,8'd200} : s = 197;
	{8'd40,8'd201} : s = 333;
	{8'd40,8'd202} : s = 331;
	{8'd40,8'd203} : s = 441;
	{8'd40,8'd204} : s = 327;
	{8'd40,8'd205} : s = 438;
	{8'd40,8'd206} : s = 437;
	{8'd40,8'd207} : s = 501;
	{8'd40,8'd208} : s = 316;
	{8'd40,8'd209} : s = 435;
	{8'd40,8'd210} : s = 430;
	{8'd40,8'd211} : s = 499;
	{8'd40,8'd212} : s = 429;
	{8'd40,8'd213} : s = 494;
	{8'd40,8'd214} : s = 493;
	{8'd40,8'd215} : s = 510;
	{8'd40,8'd216} : s = 1;
	{8'd40,8'd217} : s = 18;
	{8'd40,8'd218} : s = 17;
	{8'd40,8'd219} : s = 82;
	{8'd40,8'd220} : s = 12;
	{8'd40,8'd221} : s = 81;
	{8'd40,8'd222} : s = 76;
	{8'd40,8'd223} : s = 195;
	{8'd40,8'd224} : s = 10;
	{8'd40,8'd225} : s = 74;
	{8'd40,8'd226} : s = 73;
	{8'd40,8'd227} : s = 184;
	{8'd40,8'd228} : s = 70;
	{8'd40,8'd229} : s = 180;
	{8'd40,8'd230} : s = 178;
	{8'd40,8'd231} : s = 314;
	{8'd40,8'd232} : s = 9;
	{8'd40,8'd233} : s = 69;
	{8'd40,8'd234} : s = 67;
	{8'd40,8'd235} : s = 177;
	{8'd40,8'd236} : s = 56;
	{8'd40,8'd237} : s = 172;
	{8'd40,8'd238} : s = 170;
	{8'd40,8'd239} : s = 313;
	{8'd40,8'd240} : s = 52;
	{8'd40,8'd241} : s = 169;
	{8'd40,8'd242} : s = 166;
	{8'd40,8'd243} : s = 310;
	{8'd40,8'd244} : s = 165;
	{8'd40,8'd245} : s = 309;
	{8'd40,8'd246} : s = 307;
	{8'd40,8'd247} : s = 427;
	{8'd40,8'd248} : s = 6;
	{8'd40,8'd249} : s = 50;
	{8'd40,8'd250} : s = 49;
	{8'd40,8'd251} : s = 163;
	{8'd40,8'd252} : s = 44;
	{8'd40,8'd253} : s = 156;
	{8'd40,8'd254} : s = 154;
	{8'd40,8'd255} : s = 302;
	{8'd41,8'd0} : s = 304;
	{8'd41,8'd1} : s = 296;
	{8'd41,8'd2} : s = 432;
	{8'd41,8'd3} : s = 292;
	{8'd41,8'd4} : s = 424;
	{8'd41,8'd5} : s = 420;
	{8'd41,8'd6} : s = 488;
	{8'd41,8'd7} : s = 129;
	{8'd41,8'd8} : s = 290;
	{8'd41,8'd9} : s = 289;
	{8'd41,8'd10} : s = 418;
	{8'd41,8'd11} : s = 280;
	{8'd41,8'd12} : s = 417;
	{8'd41,8'd13} : s = 408;
	{8'd41,8'd14} : s = 484;
	{8'd41,8'd15} : s = 276;
	{8'd41,8'd16} : s = 404;
	{8'd41,8'd17} : s = 402;
	{8'd41,8'd18} : s = 482;
	{8'd41,8'd19} : s = 401;
	{8'd41,8'd20} : s = 481;
	{8'd41,8'd21} : s = 472;
	{8'd41,8'd22} : s = 504;
	{8'd41,8'd23} : s = 4;
	{8'd41,8'd24} : s = 96;
	{8'd41,8'd25} : s = 80;
	{8'd41,8'd26} : s = 274;
	{8'd41,8'd27} : s = 72;
	{8'd41,8'd28} : s = 273;
	{8'd41,8'd29} : s = 268;
	{8'd41,8'd30} : s = 396;
	{8'd41,8'd31} : s = 68;
	{8'd41,8'd32} : s = 266;
	{8'd41,8'd33} : s = 265;
	{8'd41,8'd34} : s = 394;
	{8'd41,8'd35} : s = 262;
	{8'd41,8'd36} : s = 393;
	{8'd41,8'd37} : s = 390;
	{8'd41,8'd38} : s = 468;
	{8'd41,8'd39} : s = 66;
	{8'd41,8'd40} : s = 261;
	{8'd41,8'd41} : s = 259;
	{8'd41,8'd42} : s = 389;
	{8'd41,8'd43} : s = 224;
	{8'd41,8'd44} : s = 387;
	{8'd41,8'd45} : s = 368;
	{8'd41,8'd46} : s = 466;
	{8'd41,8'd47} : s = 208;
	{8'd41,8'd48} : s = 360;
	{8'd41,8'd49} : s = 356;
	{8'd41,8'd50} : s = 465;
	{8'd41,8'd51} : s = 354;
	{8'd41,8'd52} : s = 460;
	{8'd41,8'd53} : s = 458;
	{8'd41,8'd54} : s = 500;
	{8'd41,8'd55} : s = 65;
	{8'd41,8'd56} : s = 200;
	{8'd41,8'd57} : s = 196;
	{8'd41,8'd58} : s = 353;
	{8'd41,8'd59} : s = 194;
	{8'd41,8'd60} : s = 344;
	{8'd41,8'd61} : s = 340;
	{8'd41,8'd62} : s = 457;
	{8'd41,8'd63} : s = 193;
	{8'd41,8'd64} : s = 338;
	{8'd41,8'd65} : s = 337;
	{8'd41,8'd66} : s = 454;
	{8'd41,8'd67} : s = 332;
	{8'd41,8'd68} : s = 453;
	{8'd41,8'd69} : s = 451;
	{8'd41,8'd70} : s = 498;
	{8'd41,8'd71} : s = 176;
	{8'd41,8'd72} : s = 330;
	{8'd41,8'd73} : s = 329;
	{8'd41,8'd74} : s = 440;
	{8'd41,8'd75} : s = 326;
	{8'd41,8'd76} : s = 436;
	{8'd41,8'd77} : s = 434;
	{8'd41,8'd78} : s = 497;
	{8'd41,8'd79} : s = 325;
	{8'd41,8'd80} : s = 433;
	{8'd41,8'd81} : s = 428;
	{8'd41,8'd82} : s = 492;
	{8'd41,8'd83} : s = 426;
	{8'd41,8'd84} : s = 490;
	{8'd41,8'd85} : s = 489;
	{8'd41,8'd86} : s = 508;
	{8'd41,8'd87} : s = 2;
	{8'd41,8'd88} : s = 48;
	{8'd41,8'd89} : s = 40;
	{8'd41,8'd90} : s = 168;
	{8'd41,8'd91} : s = 36;
	{8'd41,8'd92} : s = 164;
	{8'd41,8'd93} : s = 162;
	{8'd41,8'd94} : s = 323;
	{8'd41,8'd95} : s = 34;
	{8'd41,8'd96} : s = 161;
	{8'd41,8'd97} : s = 152;
	{8'd41,8'd98} : s = 312;
	{8'd41,8'd99} : s = 148;
	{8'd41,8'd100} : s = 308;
	{8'd41,8'd101} : s = 306;
	{8'd41,8'd102} : s = 425;
	{8'd41,8'd103} : s = 33;
	{8'd41,8'd104} : s = 146;
	{8'd41,8'd105} : s = 145;
	{8'd41,8'd106} : s = 305;
	{8'd41,8'd107} : s = 140;
	{8'd41,8'd108} : s = 300;
	{8'd41,8'd109} : s = 298;
	{8'd41,8'd110} : s = 422;
	{8'd41,8'd111} : s = 138;
	{8'd41,8'd112} : s = 297;
	{8'd41,8'd113} : s = 294;
	{8'd41,8'd114} : s = 421;
	{8'd41,8'd115} : s = 293;
	{8'd41,8'd116} : s = 419;
	{8'd41,8'd117} : s = 412;
	{8'd41,8'd118} : s = 486;
	{8'd41,8'd119} : s = 24;
	{8'd41,8'd120} : s = 137;
	{8'd41,8'd121} : s = 134;
	{8'd41,8'd122} : s = 291;
	{8'd41,8'd123} : s = 133;
	{8'd41,8'd124} : s = 284;
	{8'd41,8'd125} : s = 282;
	{8'd41,8'd126} : s = 410;
	{8'd41,8'd127} : s = 131;
	{8'd41,8'd128} : s = 281;
	{8'd41,8'd129} : s = 278;
	{8'd41,8'd130} : s = 409;
	{8'd41,8'd131} : s = 277;
	{8'd41,8'd132} : s = 406;
	{8'd41,8'd133} : s = 405;
	{8'd41,8'd134} : s = 485;
	{8'd41,8'd135} : s = 112;
	{8'd41,8'd136} : s = 275;
	{8'd41,8'd137} : s = 270;
	{8'd41,8'd138} : s = 403;
	{8'd41,8'd139} : s = 269;
	{8'd41,8'd140} : s = 398;
	{8'd41,8'd141} : s = 397;
	{8'd41,8'd142} : s = 483;
	{8'd41,8'd143} : s = 267;
	{8'd41,8'd144} : s = 395;
	{8'd41,8'd145} : s = 391;
	{8'd41,8'd146} : s = 476;
	{8'd41,8'd147} : s = 376;
	{8'd41,8'd148} : s = 474;
	{8'd41,8'd149} : s = 473;
	{8'd41,8'd150} : s = 506;
	{8'd41,8'd151} : s = 20;
	{8'd41,8'd152} : s = 104;
	{8'd41,8'd153} : s = 100;
	{8'd41,8'd154} : s = 263;
	{8'd41,8'd155} : s = 98;
	{8'd41,8'd156} : s = 240;
	{8'd41,8'd157} : s = 232;
	{8'd41,8'd158} : s = 372;
	{8'd41,8'd159} : s = 97;
	{8'd41,8'd160} : s = 228;
	{8'd41,8'd161} : s = 226;
	{8'd41,8'd162} : s = 370;
	{8'd41,8'd163} : s = 225;
	{8'd41,8'd164} : s = 369;
	{8'd41,8'd165} : s = 364;
	{8'd41,8'd166} : s = 470;
	{8'd41,8'd167} : s = 88;
	{8'd41,8'd168} : s = 216;
	{8'd41,8'd169} : s = 212;
	{8'd41,8'd170} : s = 362;
	{8'd41,8'd171} : s = 210;
	{8'd41,8'd172} : s = 361;
	{8'd41,8'd173} : s = 358;
	{8'd41,8'd174} : s = 469;
	{8'd41,8'd175} : s = 209;
	{8'd41,8'd176} : s = 357;
	{8'd41,8'd177} : s = 355;
	{8'd41,8'd178} : s = 467;
	{8'd41,8'd179} : s = 348;
	{8'd41,8'd180} : s = 462;
	{8'd41,8'd181} : s = 461;
	{8'd41,8'd182} : s = 505;
	{8'd41,8'd183} : s = 84;
	{8'd41,8'd184} : s = 204;
	{8'd41,8'd185} : s = 202;
	{8'd41,8'd186} : s = 346;
	{8'd41,8'd187} : s = 201;
	{8'd41,8'd188} : s = 345;
	{8'd41,8'd189} : s = 342;
	{8'd41,8'd190} : s = 459;
	{8'd41,8'd191} : s = 198;
	{8'd41,8'd192} : s = 341;
	{8'd41,8'd193} : s = 339;
	{8'd41,8'd194} : s = 455;
	{8'd41,8'd195} : s = 334;
	{8'd41,8'd196} : s = 444;
	{8'd41,8'd197} : s = 442;
	{8'd41,8'd198} : s = 502;
	{8'd41,8'd199} : s = 197;
	{8'd41,8'd200} : s = 333;
	{8'd41,8'd201} : s = 331;
	{8'd41,8'd202} : s = 441;
	{8'd41,8'd203} : s = 327;
	{8'd41,8'd204} : s = 438;
	{8'd41,8'd205} : s = 437;
	{8'd41,8'd206} : s = 501;
	{8'd41,8'd207} : s = 316;
	{8'd41,8'd208} : s = 435;
	{8'd41,8'd209} : s = 430;
	{8'd41,8'd210} : s = 499;
	{8'd41,8'd211} : s = 429;
	{8'd41,8'd212} : s = 494;
	{8'd41,8'd213} : s = 493;
	{8'd41,8'd214} : s = 510;
	{8'd41,8'd215} : s = 1;
	{8'd41,8'd216} : s = 18;
	{8'd41,8'd217} : s = 17;
	{8'd41,8'd218} : s = 82;
	{8'd41,8'd219} : s = 12;
	{8'd41,8'd220} : s = 81;
	{8'd41,8'd221} : s = 76;
	{8'd41,8'd222} : s = 195;
	{8'd41,8'd223} : s = 10;
	{8'd41,8'd224} : s = 74;
	{8'd41,8'd225} : s = 73;
	{8'd41,8'd226} : s = 184;
	{8'd41,8'd227} : s = 70;
	{8'd41,8'd228} : s = 180;
	{8'd41,8'd229} : s = 178;
	{8'd41,8'd230} : s = 314;
	{8'd41,8'd231} : s = 9;
	{8'd41,8'd232} : s = 69;
	{8'd41,8'd233} : s = 67;
	{8'd41,8'd234} : s = 177;
	{8'd41,8'd235} : s = 56;
	{8'd41,8'd236} : s = 172;
	{8'd41,8'd237} : s = 170;
	{8'd41,8'd238} : s = 313;
	{8'd41,8'd239} : s = 52;
	{8'd41,8'd240} : s = 169;
	{8'd41,8'd241} : s = 166;
	{8'd41,8'd242} : s = 310;
	{8'd41,8'd243} : s = 165;
	{8'd41,8'd244} : s = 309;
	{8'd41,8'd245} : s = 307;
	{8'd41,8'd246} : s = 427;
	{8'd41,8'd247} : s = 6;
	{8'd41,8'd248} : s = 50;
	{8'd41,8'd249} : s = 49;
	{8'd41,8'd250} : s = 163;
	{8'd41,8'd251} : s = 44;
	{8'd41,8'd252} : s = 156;
	{8'd41,8'd253} : s = 154;
	{8'd41,8'd254} : s = 302;
	{8'd41,8'd255} : s = 42;
	{8'd42,8'd0} : s = 296;
	{8'd42,8'd1} : s = 432;
	{8'd42,8'd2} : s = 292;
	{8'd42,8'd3} : s = 424;
	{8'd42,8'd4} : s = 420;
	{8'd42,8'd5} : s = 488;
	{8'd42,8'd6} : s = 129;
	{8'd42,8'd7} : s = 290;
	{8'd42,8'd8} : s = 289;
	{8'd42,8'd9} : s = 418;
	{8'd42,8'd10} : s = 280;
	{8'd42,8'd11} : s = 417;
	{8'd42,8'd12} : s = 408;
	{8'd42,8'd13} : s = 484;
	{8'd42,8'd14} : s = 276;
	{8'd42,8'd15} : s = 404;
	{8'd42,8'd16} : s = 402;
	{8'd42,8'd17} : s = 482;
	{8'd42,8'd18} : s = 401;
	{8'd42,8'd19} : s = 481;
	{8'd42,8'd20} : s = 472;
	{8'd42,8'd21} : s = 504;
	{8'd42,8'd22} : s = 4;
	{8'd42,8'd23} : s = 96;
	{8'd42,8'd24} : s = 80;
	{8'd42,8'd25} : s = 274;
	{8'd42,8'd26} : s = 72;
	{8'd42,8'd27} : s = 273;
	{8'd42,8'd28} : s = 268;
	{8'd42,8'd29} : s = 396;
	{8'd42,8'd30} : s = 68;
	{8'd42,8'd31} : s = 266;
	{8'd42,8'd32} : s = 265;
	{8'd42,8'd33} : s = 394;
	{8'd42,8'd34} : s = 262;
	{8'd42,8'd35} : s = 393;
	{8'd42,8'd36} : s = 390;
	{8'd42,8'd37} : s = 468;
	{8'd42,8'd38} : s = 66;
	{8'd42,8'd39} : s = 261;
	{8'd42,8'd40} : s = 259;
	{8'd42,8'd41} : s = 389;
	{8'd42,8'd42} : s = 224;
	{8'd42,8'd43} : s = 387;
	{8'd42,8'd44} : s = 368;
	{8'd42,8'd45} : s = 466;
	{8'd42,8'd46} : s = 208;
	{8'd42,8'd47} : s = 360;
	{8'd42,8'd48} : s = 356;
	{8'd42,8'd49} : s = 465;
	{8'd42,8'd50} : s = 354;
	{8'd42,8'd51} : s = 460;
	{8'd42,8'd52} : s = 458;
	{8'd42,8'd53} : s = 500;
	{8'd42,8'd54} : s = 65;
	{8'd42,8'd55} : s = 200;
	{8'd42,8'd56} : s = 196;
	{8'd42,8'd57} : s = 353;
	{8'd42,8'd58} : s = 194;
	{8'd42,8'd59} : s = 344;
	{8'd42,8'd60} : s = 340;
	{8'd42,8'd61} : s = 457;
	{8'd42,8'd62} : s = 193;
	{8'd42,8'd63} : s = 338;
	{8'd42,8'd64} : s = 337;
	{8'd42,8'd65} : s = 454;
	{8'd42,8'd66} : s = 332;
	{8'd42,8'd67} : s = 453;
	{8'd42,8'd68} : s = 451;
	{8'd42,8'd69} : s = 498;
	{8'd42,8'd70} : s = 176;
	{8'd42,8'd71} : s = 330;
	{8'd42,8'd72} : s = 329;
	{8'd42,8'd73} : s = 440;
	{8'd42,8'd74} : s = 326;
	{8'd42,8'd75} : s = 436;
	{8'd42,8'd76} : s = 434;
	{8'd42,8'd77} : s = 497;
	{8'd42,8'd78} : s = 325;
	{8'd42,8'd79} : s = 433;
	{8'd42,8'd80} : s = 428;
	{8'd42,8'd81} : s = 492;
	{8'd42,8'd82} : s = 426;
	{8'd42,8'd83} : s = 490;
	{8'd42,8'd84} : s = 489;
	{8'd42,8'd85} : s = 508;
	{8'd42,8'd86} : s = 2;
	{8'd42,8'd87} : s = 48;
	{8'd42,8'd88} : s = 40;
	{8'd42,8'd89} : s = 168;
	{8'd42,8'd90} : s = 36;
	{8'd42,8'd91} : s = 164;
	{8'd42,8'd92} : s = 162;
	{8'd42,8'd93} : s = 323;
	{8'd42,8'd94} : s = 34;
	{8'd42,8'd95} : s = 161;
	{8'd42,8'd96} : s = 152;
	{8'd42,8'd97} : s = 312;
	{8'd42,8'd98} : s = 148;
	{8'd42,8'd99} : s = 308;
	{8'd42,8'd100} : s = 306;
	{8'd42,8'd101} : s = 425;
	{8'd42,8'd102} : s = 33;
	{8'd42,8'd103} : s = 146;
	{8'd42,8'd104} : s = 145;
	{8'd42,8'd105} : s = 305;
	{8'd42,8'd106} : s = 140;
	{8'd42,8'd107} : s = 300;
	{8'd42,8'd108} : s = 298;
	{8'd42,8'd109} : s = 422;
	{8'd42,8'd110} : s = 138;
	{8'd42,8'd111} : s = 297;
	{8'd42,8'd112} : s = 294;
	{8'd42,8'd113} : s = 421;
	{8'd42,8'd114} : s = 293;
	{8'd42,8'd115} : s = 419;
	{8'd42,8'd116} : s = 412;
	{8'd42,8'd117} : s = 486;
	{8'd42,8'd118} : s = 24;
	{8'd42,8'd119} : s = 137;
	{8'd42,8'd120} : s = 134;
	{8'd42,8'd121} : s = 291;
	{8'd42,8'd122} : s = 133;
	{8'd42,8'd123} : s = 284;
	{8'd42,8'd124} : s = 282;
	{8'd42,8'd125} : s = 410;
	{8'd42,8'd126} : s = 131;
	{8'd42,8'd127} : s = 281;
	{8'd42,8'd128} : s = 278;
	{8'd42,8'd129} : s = 409;
	{8'd42,8'd130} : s = 277;
	{8'd42,8'd131} : s = 406;
	{8'd42,8'd132} : s = 405;
	{8'd42,8'd133} : s = 485;
	{8'd42,8'd134} : s = 112;
	{8'd42,8'd135} : s = 275;
	{8'd42,8'd136} : s = 270;
	{8'd42,8'd137} : s = 403;
	{8'd42,8'd138} : s = 269;
	{8'd42,8'd139} : s = 398;
	{8'd42,8'd140} : s = 397;
	{8'd42,8'd141} : s = 483;
	{8'd42,8'd142} : s = 267;
	{8'd42,8'd143} : s = 395;
	{8'd42,8'd144} : s = 391;
	{8'd42,8'd145} : s = 476;
	{8'd42,8'd146} : s = 376;
	{8'd42,8'd147} : s = 474;
	{8'd42,8'd148} : s = 473;
	{8'd42,8'd149} : s = 506;
	{8'd42,8'd150} : s = 20;
	{8'd42,8'd151} : s = 104;
	{8'd42,8'd152} : s = 100;
	{8'd42,8'd153} : s = 263;
	{8'd42,8'd154} : s = 98;
	{8'd42,8'd155} : s = 240;
	{8'd42,8'd156} : s = 232;
	{8'd42,8'd157} : s = 372;
	{8'd42,8'd158} : s = 97;
	{8'd42,8'd159} : s = 228;
	{8'd42,8'd160} : s = 226;
	{8'd42,8'd161} : s = 370;
	{8'd42,8'd162} : s = 225;
	{8'd42,8'd163} : s = 369;
	{8'd42,8'd164} : s = 364;
	{8'd42,8'd165} : s = 470;
	{8'd42,8'd166} : s = 88;
	{8'd42,8'd167} : s = 216;
	{8'd42,8'd168} : s = 212;
	{8'd42,8'd169} : s = 362;
	{8'd42,8'd170} : s = 210;
	{8'd42,8'd171} : s = 361;
	{8'd42,8'd172} : s = 358;
	{8'd42,8'd173} : s = 469;
	{8'd42,8'd174} : s = 209;
	{8'd42,8'd175} : s = 357;
	{8'd42,8'd176} : s = 355;
	{8'd42,8'd177} : s = 467;
	{8'd42,8'd178} : s = 348;
	{8'd42,8'd179} : s = 462;
	{8'd42,8'd180} : s = 461;
	{8'd42,8'd181} : s = 505;
	{8'd42,8'd182} : s = 84;
	{8'd42,8'd183} : s = 204;
	{8'd42,8'd184} : s = 202;
	{8'd42,8'd185} : s = 346;
	{8'd42,8'd186} : s = 201;
	{8'd42,8'd187} : s = 345;
	{8'd42,8'd188} : s = 342;
	{8'd42,8'd189} : s = 459;
	{8'd42,8'd190} : s = 198;
	{8'd42,8'd191} : s = 341;
	{8'd42,8'd192} : s = 339;
	{8'd42,8'd193} : s = 455;
	{8'd42,8'd194} : s = 334;
	{8'd42,8'd195} : s = 444;
	{8'd42,8'd196} : s = 442;
	{8'd42,8'd197} : s = 502;
	{8'd42,8'd198} : s = 197;
	{8'd42,8'd199} : s = 333;
	{8'd42,8'd200} : s = 331;
	{8'd42,8'd201} : s = 441;
	{8'd42,8'd202} : s = 327;
	{8'd42,8'd203} : s = 438;
	{8'd42,8'd204} : s = 437;
	{8'd42,8'd205} : s = 501;
	{8'd42,8'd206} : s = 316;
	{8'd42,8'd207} : s = 435;
	{8'd42,8'd208} : s = 430;
	{8'd42,8'd209} : s = 499;
	{8'd42,8'd210} : s = 429;
	{8'd42,8'd211} : s = 494;
	{8'd42,8'd212} : s = 493;
	{8'd42,8'd213} : s = 510;
	{8'd42,8'd214} : s = 1;
	{8'd42,8'd215} : s = 18;
	{8'd42,8'd216} : s = 17;
	{8'd42,8'd217} : s = 82;
	{8'd42,8'd218} : s = 12;
	{8'd42,8'd219} : s = 81;
	{8'd42,8'd220} : s = 76;
	{8'd42,8'd221} : s = 195;
	{8'd42,8'd222} : s = 10;
	{8'd42,8'd223} : s = 74;
	{8'd42,8'd224} : s = 73;
	{8'd42,8'd225} : s = 184;
	{8'd42,8'd226} : s = 70;
	{8'd42,8'd227} : s = 180;
	{8'd42,8'd228} : s = 178;
	{8'd42,8'd229} : s = 314;
	{8'd42,8'd230} : s = 9;
	{8'd42,8'd231} : s = 69;
	{8'd42,8'd232} : s = 67;
	{8'd42,8'd233} : s = 177;
	{8'd42,8'd234} : s = 56;
	{8'd42,8'd235} : s = 172;
	{8'd42,8'd236} : s = 170;
	{8'd42,8'd237} : s = 313;
	{8'd42,8'd238} : s = 52;
	{8'd42,8'd239} : s = 169;
	{8'd42,8'd240} : s = 166;
	{8'd42,8'd241} : s = 310;
	{8'd42,8'd242} : s = 165;
	{8'd42,8'd243} : s = 309;
	{8'd42,8'd244} : s = 307;
	{8'd42,8'd245} : s = 427;
	{8'd42,8'd246} : s = 6;
	{8'd42,8'd247} : s = 50;
	{8'd42,8'd248} : s = 49;
	{8'd42,8'd249} : s = 163;
	{8'd42,8'd250} : s = 44;
	{8'd42,8'd251} : s = 156;
	{8'd42,8'd252} : s = 154;
	{8'd42,8'd253} : s = 302;
	{8'd42,8'd254} : s = 42;
	{8'd42,8'd255} : s = 153;
	{8'd43,8'd0} : s = 432;
	{8'd43,8'd1} : s = 292;
	{8'd43,8'd2} : s = 424;
	{8'd43,8'd3} : s = 420;
	{8'd43,8'd4} : s = 488;
	{8'd43,8'd5} : s = 129;
	{8'd43,8'd6} : s = 290;
	{8'd43,8'd7} : s = 289;
	{8'd43,8'd8} : s = 418;
	{8'd43,8'd9} : s = 280;
	{8'd43,8'd10} : s = 417;
	{8'd43,8'd11} : s = 408;
	{8'd43,8'd12} : s = 484;
	{8'd43,8'd13} : s = 276;
	{8'd43,8'd14} : s = 404;
	{8'd43,8'd15} : s = 402;
	{8'd43,8'd16} : s = 482;
	{8'd43,8'd17} : s = 401;
	{8'd43,8'd18} : s = 481;
	{8'd43,8'd19} : s = 472;
	{8'd43,8'd20} : s = 504;
	{8'd43,8'd21} : s = 4;
	{8'd43,8'd22} : s = 96;
	{8'd43,8'd23} : s = 80;
	{8'd43,8'd24} : s = 274;
	{8'd43,8'd25} : s = 72;
	{8'd43,8'd26} : s = 273;
	{8'd43,8'd27} : s = 268;
	{8'd43,8'd28} : s = 396;
	{8'd43,8'd29} : s = 68;
	{8'd43,8'd30} : s = 266;
	{8'd43,8'd31} : s = 265;
	{8'd43,8'd32} : s = 394;
	{8'd43,8'd33} : s = 262;
	{8'd43,8'd34} : s = 393;
	{8'd43,8'd35} : s = 390;
	{8'd43,8'd36} : s = 468;
	{8'd43,8'd37} : s = 66;
	{8'd43,8'd38} : s = 261;
	{8'd43,8'd39} : s = 259;
	{8'd43,8'd40} : s = 389;
	{8'd43,8'd41} : s = 224;
	{8'd43,8'd42} : s = 387;
	{8'd43,8'd43} : s = 368;
	{8'd43,8'd44} : s = 466;
	{8'd43,8'd45} : s = 208;
	{8'd43,8'd46} : s = 360;
	{8'd43,8'd47} : s = 356;
	{8'd43,8'd48} : s = 465;
	{8'd43,8'd49} : s = 354;
	{8'd43,8'd50} : s = 460;
	{8'd43,8'd51} : s = 458;
	{8'd43,8'd52} : s = 500;
	{8'd43,8'd53} : s = 65;
	{8'd43,8'd54} : s = 200;
	{8'd43,8'd55} : s = 196;
	{8'd43,8'd56} : s = 353;
	{8'd43,8'd57} : s = 194;
	{8'd43,8'd58} : s = 344;
	{8'd43,8'd59} : s = 340;
	{8'd43,8'd60} : s = 457;
	{8'd43,8'd61} : s = 193;
	{8'd43,8'd62} : s = 338;
	{8'd43,8'd63} : s = 337;
	{8'd43,8'd64} : s = 454;
	{8'd43,8'd65} : s = 332;
	{8'd43,8'd66} : s = 453;
	{8'd43,8'd67} : s = 451;
	{8'd43,8'd68} : s = 498;
	{8'd43,8'd69} : s = 176;
	{8'd43,8'd70} : s = 330;
	{8'd43,8'd71} : s = 329;
	{8'd43,8'd72} : s = 440;
	{8'd43,8'd73} : s = 326;
	{8'd43,8'd74} : s = 436;
	{8'd43,8'd75} : s = 434;
	{8'd43,8'd76} : s = 497;
	{8'd43,8'd77} : s = 325;
	{8'd43,8'd78} : s = 433;
	{8'd43,8'd79} : s = 428;
	{8'd43,8'd80} : s = 492;
	{8'd43,8'd81} : s = 426;
	{8'd43,8'd82} : s = 490;
	{8'd43,8'd83} : s = 489;
	{8'd43,8'd84} : s = 508;
	{8'd43,8'd85} : s = 2;
	{8'd43,8'd86} : s = 48;
	{8'd43,8'd87} : s = 40;
	{8'd43,8'd88} : s = 168;
	{8'd43,8'd89} : s = 36;
	{8'd43,8'd90} : s = 164;
	{8'd43,8'd91} : s = 162;
	{8'd43,8'd92} : s = 323;
	{8'd43,8'd93} : s = 34;
	{8'd43,8'd94} : s = 161;
	{8'd43,8'd95} : s = 152;
	{8'd43,8'd96} : s = 312;
	{8'd43,8'd97} : s = 148;
	{8'd43,8'd98} : s = 308;
	{8'd43,8'd99} : s = 306;
	{8'd43,8'd100} : s = 425;
	{8'd43,8'd101} : s = 33;
	{8'd43,8'd102} : s = 146;
	{8'd43,8'd103} : s = 145;
	{8'd43,8'd104} : s = 305;
	{8'd43,8'd105} : s = 140;
	{8'd43,8'd106} : s = 300;
	{8'd43,8'd107} : s = 298;
	{8'd43,8'd108} : s = 422;
	{8'd43,8'd109} : s = 138;
	{8'd43,8'd110} : s = 297;
	{8'd43,8'd111} : s = 294;
	{8'd43,8'd112} : s = 421;
	{8'd43,8'd113} : s = 293;
	{8'd43,8'd114} : s = 419;
	{8'd43,8'd115} : s = 412;
	{8'd43,8'd116} : s = 486;
	{8'd43,8'd117} : s = 24;
	{8'd43,8'd118} : s = 137;
	{8'd43,8'd119} : s = 134;
	{8'd43,8'd120} : s = 291;
	{8'd43,8'd121} : s = 133;
	{8'd43,8'd122} : s = 284;
	{8'd43,8'd123} : s = 282;
	{8'd43,8'd124} : s = 410;
	{8'd43,8'd125} : s = 131;
	{8'd43,8'd126} : s = 281;
	{8'd43,8'd127} : s = 278;
	{8'd43,8'd128} : s = 409;
	{8'd43,8'd129} : s = 277;
	{8'd43,8'd130} : s = 406;
	{8'd43,8'd131} : s = 405;
	{8'd43,8'd132} : s = 485;
	{8'd43,8'd133} : s = 112;
	{8'd43,8'd134} : s = 275;
	{8'd43,8'd135} : s = 270;
	{8'd43,8'd136} : s = 403;
	{8'd43,8'd137} : s = 269;
	{8'd43,8'd138} : s = 398;
	{8'd43,8'd139} : s = 397;
	{8'd43,8'd140} : s = 483;
	{8'd43,8'd141} : s = 267;
	{8'd43,8'd142} : s = 395;
	{8'd43,8'd143} : s = 391;
	{8'd43,8'd144} : s = 476;
	{8'd43,8'd145} : s = 376;
	{8'd43,8'd146} : s = 474;
	{8'd43,8'd147} : s = 473;
	{8'd43,8'd148} : s = 506;
	{8'd43,8'd149} : s = 20;
	{8'd43,8'd150} : s = 104;
	{8'd43,8'd151} : s = 100;
	{8'd43,8'd152} : s = 263;
	{8'd43,8'd153} : s = 98;
	{8'd43,8'd154} : s = 240;
	{8'd43,8'd155} : s = 232;
	{8'd43,8'd156} : s = 372;
	{8'd43,8'd157} : s = 97;
	{8'd43,8'd158} : s = 228;
	{8'd43,8'd159} : s = 226;
	{8'd43,8'd160} : s = 370;
	{8'd43,8'd161} : s = 225;
	{8'd43,8'd162} : s = 369;
	{8'd43,8'd163} : s = 364;
	{8'd43,8'd164} : s = 470;
	{8'd43,8'd165} : s = 88;
	{8'd43,8'd166} : s = 216;
	{8'd43,8'd167} : s = 212;
	{8'd43,8'd168} : s = 362;
	{8'd43,8'd169} : s = 210;
	{8'd43,8'd170} : s = 361;
	{8'd43,8'd171} : s = 358;
	{8'd43,8'd172} : s = 469;
	{8'd43,8'd173} : s = 209;
	{8'd43,8'd174} : s = 357;
	{8'd43,8'd175} : s = 355;
	{8'd43,8'd176} : s = 467;
	{8'd43,8'd177} : s = 348;
	{8'd43,8'd178} : s = 462;
	{8'd43,8'd179} : s = 461;
	{8'd43,8'd180} : s = 505;
	{8'd43,8'd181} : s = 84;
	{8'd43,8'd182} : s = 204;
	{8'd43,8'd183} : s = 202;
	{8'd43,8'd184} : s = 346;
	{8'd43,8'd185} : s = 201;
	{8'd43,8'd186} : s = 345;
	{8'd43,8'd187} : s = 342;
	{8'd43,8'd188} : s = 459;
	{8'd43,8'd189} : s = 198;
	{8'd43,8'd190} : s = 341;
	{8'd43,8'd191} : s = 339;
	{8'd43,8'd192} : s = 455;
	{8'd43,8'd193} : s = 334;
	{8'd43,8'd194} : s = 444;
	{8'd43,8'd195} : s = 442;
	{8'd43,8'd196} : s = 502;
	{8'd43,8'd197} : s = 197;
	{8'd43,8'd198} : s = 333;
	{8'd43,8'd199} : s = 331;
	{8'd43,8'd200} : s = 441;
	{8'd43,8'd201} : s = 327;
	{8'd43,8'd202} : s = 438;
	{8'd43,8'd203} : s = 437;
	{8'd43,8'd204} : s = 501;
	{8'd43,8'd205} : s = 316;
	{8'd43,8'd206} : s = 435;
	{8'd43,8'd207} : s = 430;
	{8'd43,8'd208} : s = 499;
	{8'd43,8'd209} : s = 429;
	{8'd43,8'd210} : s = 494;
	{8'd43,8'd211} : s = 493;
	{8'd43,8'd212} : s = 510;
	{8'd43,8'd213} : s = 1;
	{8'd43,8'd214} : s = 18;
	{8'd43,8'd215} : s = 17;
	{8'd43,8'd216} : s = 82;
	{8'd43,8'd217} : s = 12;
	{8'd43,8'd218} : s = 81;
	{8'd43,8'd219} : s = 76;
	{8'd43,8'd220} : s = 195;
	{8'd43,8'd221} : s = 10;
	{8'd43,8'd222} : s = 74;
	{8'd43,8'd223} : s = 73;
	{8'd43,8'd224} : s = 184;
	{8'd43,8'd225} : s = 70;
	{8'd43,8'd226} : s = 180;
	{8'd43,8'd227} : s = 178;
	{8'd43,8'd228} : s = 314;
	{8'd43,8'd229} : s = 9;
	{8'd43,8'd230} : s = 69;
	{8'd43,8'd231} : s = 67;
	{8'd43,8'd232} : s = 177;
	{8'd43,8'd233} : s = 56;
	{8'd43,8'd234} : s = 172;
	{8'd43,8'd235} : s = 170;
	{8'd43,8'd236} : s = 313;
	{8'd43,8'd237} : s = 52;
	{8'd43,8'd238} : s = 169;
	{8'd43,8'd239} : s = 166;
	{8'd43,8'd240} : s = 310;
	{8'd43,8'd241} : s = 165;
	{8'd43,8'd242} : s = 309;
	{8'd43,8'd243} : s = 307;
	{8'd43,8'd244} : s = 427;
	{8'd43,8'd245} : s = 6;
	{8'd43,8'd246} : s = 50;
	{8'd43,8'd247} : s = 49;
	{8'd43,8'd248} : s = 163;
	{8'd43,8'd249} : s = 44;
	{8'd43,8'd250} : s = 156;
	{8'd43,8'd251} : s = 154;
	{8'd43,8'd252} : s = 302;
	{8'd43,8'd253} : s = 42;
	{8'd43,8'd254} : s = 153;
	{8'd43,8'd255} : s = 150;
	{8'd44,8'd0} : s = 292;
	{8'd44,8'd1} : s = 424;
	{8'd44,8'd2} : s = 420;
	{8'd44,8'd3} : s = 488;
	{8'd44,8'd4} : s = 129;
	{8'd44,8'd5} : s = 290;
	{8'd44,8'd6} : s = 289;
	{8'd44,8'd7} : s = 418;
	{8'd44,8'd8} : s = 280;
	{8'd44,8'd9} : s = 417;
	{8'd44,8'd10} : s = 408;
	{8'd44,8'd11} : s = 484;
	{8'd44,8'd12} : s = 276;
	{8'd44,8'd13} : s = 404;
	{8'd44,8'd14} : s = 402;
	{8'd44,8'd15} : s = 482;
	{8'd44,8'd16} : s = 401;
	{8'd44,8'd17} : s = 481;
	{8'd44,8'd18} : s = 472;
	{8'd44,8'd19} : s = 504;
	{8'd44,8'd20} : s = 4;
	{8'd44,8'd21} : s = 96;
	{8'd44,8'd22} : s = 80;
	{8'd44,8'd23} : s = 274;
	{8'd44,8'd24} : s = 72;
	{8'd44,8'd25} : s = 273;
	{8'd44,8'd26} : s = 268;
	{8'd44,8'd27} : s = 396;
	{8'd44,8'd28} : s = 68;
	{8'd44,8'd29} : s = 266;
	{8'd44,8'd30} : s = 265;
	{8'd44,8'd31} : s = 394;
	{8'd44,8'd32} : s = 262;
	{8'd44,8'd33} : s = 393;
	{8'd44,8'd34} : s = 390;
	{8'd44,8'd35} : s = 468;
	{8'd44,8'd36} : s = 66;
	{8'd44,8'd37} : s = 261;
	{8'd44,8'd38} : s = 259;
	{8'd44,8'd39} : s = 389;
	{8'd44,8'd40} : s = 224;
	{8'd44,8'd41} : s = 387;
	{8'd44,8'd42} : s = 368;
	{8'd44,8'd43} : s = 466;
	{8'd44,8'd44} : s = 208;
	{8'd44,8'd45} : s = 360;
	{8'd44,8'd46} : s = 356;
	{8'd44,8'd47} : s = 465;
	{8'd44,8'd48} : s = 354;
	{8'd44,8'd49} : s = 460;
	{8'd44,8'd50} : s = 458;
	{8'd44,8'd51} : s = 500;
	{8'd44,8'd52} : s = 65;
	{8'd44,8'd53} : s = 200;
	{8'd44,8'd54} : s = 196;
	{8'd44,8'd55} : s = 353;
	{8'd44,8'd56} : s = 194;
	{8'd44,8'd57} : s = 344;
	{8'd44,8'd58} : s = 340;
	{8'd44,8'd59} : s = 457;
	{8'd44,8'd60} : s = 193;
	{8'd44,8'd61} : s = 338;
	{8'd44,8'd62} : s = 337;
	{8'd44,8'd63} : s = 454;
	{8'd44,8'd64} : s = 332;
	{8'd44,8'd65} : s = 453;
	{8'd44,8'd66} : s = 451;
	{8'd44,8'd67} : s = 498;
	{8'd44,8'd68} : s = 176;
	{8'd44,8'd69} : s = 330;
	{8'd44,8'd70} : s = 329;
	{8'd44,8'd71} : s = 440;
	{8'd44,8'd72} : s = 326;
	{8'd44,8'd73} : s = 436;
	{8'd44,8'd74} : s = 434;
	{8'd44,8'd75} : s = 497;
	{8'd44,8'd76} : s = 325;
	{8'd44,8'd77} : s = 433;
	{8'd44,8'd78} : s = 428;
	{8'd44,8'd79} : s = 492;
	{8'd44,8'd80} : s = 426;
	{8'd44,8'd81} : s = 490;
	{8'd44,8'd82} : s = 489;
	{8'd44,8'd83} : s = 508;
	{8'd44,8'd84} : s = 2;
	{8'd44,8'd85} : s = 48;
	{8'd44,8'd86} : s = 40;
	{8'd44,8'd87} : s = 168;
	{8'd44,8'd88} : s = 36;
	{8'd44,8'd89} : s = 164;
	{8'd44,8'd90} : s = 162;
	{8'd44,8'd91} : s = 323;
	{8'd44,8'd92} : s = 34;
	{8'd44,8'd93} : s = 161;
	{8'd44,8'd94} : s = 152;
	{8'd44,8'd95} : s = 312;
	{8'd44,8'd96} : s = 148;
	{8'd44,8'd97} : s = 308;
	{8'd44,8'd98} : s = 306;
	{8'd44,8'd99} : s = 425;
	{8'd44,8'd100} : s = 33;
	{8'd44,8'd101} : s = 146;
	{8'd44,8'd102} : s = 145;
	{8'd44,8'd103} : s = 305;
	{8'd44,8'd104} : s = 140;
	{8'd44,8'd105} : s = 300;
	{8'd44,8'd106} : s = 298;
	{8'd44,8'd107} : s = 422;
	{8'd44,8'd108} : s = 138;
	{8'd44,8'd109} : s = 297;
	{8'd44,8'd110} : s = 294;
	{8'd44,8'd111} : s = 421;
	{8'd44,8'd112} : s = 293;
	{8'd44,8'd113} : s = 419;
	{8'd44,8'd114} : s = 412;
	{8'd44,8'd115} : s = 486;
	{8'd44,8'd116} : s = 24;
	{8'd44,8'd117} : s = 137;
	{8'd44,8'd118} : s = 134;
	{8'd44,8'd119} : s = 291;
	{8'd44,8'd120} : s = 133;
	{8'd44,8'd121} : s = 284;
	{8'd44,8'd122} : s = 282;
	{8'd44,8'd123} : s = 410;
	{8'd44,8'd124} : s = 131;
	{8'd44,8'd125} : s = 281;
	{8'd44,8'd126} : s = 278;
	{8'd44,8'd127} : s = 409;
	{8'd44,8'd128} : s = 277;
	{8'd44,8'd129} : s = 406;
	{8'd44,8'd130} : s = 405;
	{8'd44,8'd131} : s = 485;
	{8'd44,8'd132} : s = 112;
	{8'd44,8'd133} : s = 275;
	{8'd44,8'd134} : s = 270;
	{8'd44,8'd135} : s = 403;
	{8'd44,8'd136} : s = 269;
	{8'd44,8'd137} : s = 398;
	{8'd44,8'd138} : s = 397;
	{8'd44,8'd139} : s = 483;
	{8'd44,8'd140} : s = 267;
	{8'd44,8'd141} : s = 395;
	{8'd44,8'd142} : s = 391;
	{8'd44,8'd143} : s = 476;
	{8'd44,8'd144} : s = 376;
	{8'd44,8'd145} : s = 474;
	{8'd44,8'd146} : s = 473;
	{8'd44,8'd147} : s = 506;
	{8'd44,8'd148} : s = 20;
	{8'd44,8'd149} : s = 104;
	{8'd44,8'd150} : s = 100;
	{8'd44,8'd151} : s = 263;
	{8'd44,8'd152} : s = 98;
	{8'd44,8'd153} : s = 240;
	{8'd44,8'd154} : s = 232;
	{8'd44,8'd155} : s = 372;
	{8'd44,8'd156} : s = 97;
	{8'd44,8'd157} : s = 228;
	{8'd44,8'd158} : s = 226;
	{8'd44,8'd159} : s = 370;
	{8'd44,8'd160} : s = 225;
	{8'd44,8'd161} : s = 369;
	{8'd44,8'd162} : s = 364;
	{8'd44,8'd163} : s = 470;
	{8'd44,8'd164} : s = 88;
	{8'd44,8'd165} : s = 216;
	{8'd44,8'd166} : s = 212;
	{8'd44,8'd167} : s = 362;
	{8'd44,8'd168} : s = 210;
	{8'd44,8'd169} : s = 361;
	{8'd44,8'd170} : s = 358;
	{8'd44,8'd171} : s = 469;
	{8'd44,8'd172} : s = 209;
	{8'd44,8'd173} : s = 357;
	{8'd44,8'd174} : s = 355;
	{8'd44,8'd175} : s = 467;
	{8'd44,8'd176} : s = 348;
	{8'd44,8'd177} : s = 462;
	{8'd44,8'd178} : s = 461;
	{8'd44,8'd179} : s = 505;
	{8'd44,8'd180} : s = 84;
	{8'd44,8'd181} : s = 204;
	{8'd44,8'd182} : s = 202;
	{8'd44,8'd183} : s = 346;
	{8'd44,8'd184} : s = 201;
	{8'd44,8'd185} : s = 345;
	{8'd44,8'd186} : s = 342;
	{8'd44,8'd187} : s = 459;
	{8'd44,8'd188} : s = 198;
	{8'd44,8'd189} : s = 341;
	{8'd44,8'd190} : s = 339;
	{8'd44,8'd191} : s = 455;
	{8'd44,8'd192} : s = 334;
	{8'd44,8'd193} : s = 444;
	{8'd44,8'd194} : s = 442;
	{8'd44,8'd195} : s = 502;
	{8'd44,8'd196} : s = 197;
	{8'd44,8'd197} : s = 333;
	{8'd44,8'd198} : s = 331;
	{8'd44,8'd199} : s = 441;
	{8'd44,8'd200} : s = 327;
	{8'd44,8'd201} : s = 438;
	{8'd44,8'd202} : s = 437;
	{8'd44,8'd203} : s = 501;
	{8'd44,8'd204} : s = 316;
	{8'd44,8'd205} : s = 435;
	{8'd44,8'd206} : s = 430;
	{8'd44,8'd207} : s = 499;
	{8'd44,8'd208} : s = 429;
	{8'd44,8'd209} : s = 494;
	{8'd44,8'd210} : s = 493;
	{8'd44,8'd211} : s = 510;
	{8'd44,8'd212} : s = 1;
	{8'd44,8'd213} : s = 18;
	{8'd44,8'd214} : s = 17;
	{8'd44,8'd215} : s = 82;
	{8'd44,8'd216} : s = 12;
	{8'd44,8'd217} : s = 81;
	{8'd44,8'd218} : s = 76;
	{8'd44,8'd219} : s = 195;
	{8'd44,8'd220} : s = 10;
	{8'd44,8'd221} : s = 74;
	{8'd44,8'd222} : s = 73;
	{8'd44,8'd223} : s = 184;
	{8'd44,8'd224} : s = 70;
	{8'd44,8'd225} : s = 180;
	{8'd44,8'd226} : s = 178;
	{8'd44,8'd227} : s = 314;
	{8'd44,8'd228} : s = 9;
	{8'd44,8'd229} : s = 69;
	{8'd44,8'd230} : s = 67;
	{8'd44,8'd231} : s = 177;
	{8'd44,8'd232} : s = 56;
	{8'd44,8'd233} : s = 172;
	{8'd44,8'd234} : s = 170;
	{8'd44,8'd235} : s = 313;
	{8'd44,8'd236} : s = 52;
	{8'd44,8'd237} : s = 169;
	{8'd44,8'd238} : s = 166;
	{8'd44,8'd239} : s = 310;
	{8'd44,8'd240} : s = 165;
	{8'd44,8'd241} : s = 309;
	{8'd44,8'd242} : s = 307;
	{8'd44,8'd243} : s = 427;
	{8'd44,8'd244} : s = 6;
	{8'd44,8'd245} : s = 50;
	{8'd44,8'd246} : s = 49;
	{8'd44,8'd247} : s = 163;
	{8'd44,8'd248} : s = 44;
	{8'd44,8'd249} : s = 156;
	{8'd44,8'd250} : s = 154;
	{8'd44,8'd251} : s = 302;
	{8'd44,8'd252} : s = 42;
	{8'd44,8'd253} : s = 153;
	{8'd44,8'd254} : s = 150;
	{8'd44,8'd255} : s = 301;
	{8'd45,8'd0} : s = 424;
	{8'd45,8'd1} : s = 420;
	{8'd45,8'd2} : s = 488;
	{8'd45,8'd3} : s = 129;
	{8'd45,8'd4} : s = 290;
	{8'd45,8'd5} : s = 289;
	{8'd45,8'd6} : s = 418;
	{8'd45,8'd7} : s = 280;
	{8'd45,8'd8} : s = 417;
	{8'd45,8'd9} : s = 408;
	{8'd45,8'd10} : s = 484;
	{8'd45,8'd11} : s = 276;
	{8'd45,8'd12} : s = 404;
	{8'd45,8'd13} : s = 402;
	{8'd45,8'd14} : s = 482;
	{8'd45,8'd15} : s = 401;
	{8'd45,8'd16} : s = 481;
	{8'd45,8'd17} : s = 472;
	{8'd45,8'd18} : s = 504;
	{8'd45,8'd19} : s = 4;
	{8'd45,8'd20} : s = 96;
	{8'd45,8'd21} : s = 80;
	{8'd45,8'd22} : s = 274;
	{8'd45,8'd23} : s = 72;
	{8'd45,8'd24} : s = 273;
	{8'd45,8'd25} : s = 268;
	{8'd45,8'd26} : s = 396;
	{8'd45,8'd27} : s = 68;
	{8'd45,8'd28} : s = 266;
	{8'd45,8'd29} : s = 265;
	{8'd45,8'd30} : s = 394;
	{8'd45,8'd31} : s = 262;
	{8'd45,8'd32} : s = 393;
	{8'd45,8'd33} : s = 390;
	{8'd45,8'd34} : s = 468;
	{8'd45,8'd35} : s = 66;
	{8'd45,8'd36} : s = 261;
	{8'd45,8'd37} : s = 259;
	{8'd45,8'd38} : s = 389;
	{8'd45,8'd39} : s = 224;
	{8'd45,8'd40} : s = 387;
	{8'd45,8'd41} : s = 368;
	{8'd45,8'd42} : s = 466;
	{8'd45,8'd43} : s = 208;
	{8'd45,8'd44} : s = 360;
	{8'd45,8'd45} : s = 356;
	{8'd45,8'd46} : s = 465;
	{8'd45,8'd47} : s = 354;
	{8'd45,8'd48} : s = 460;
	{8'd45,8'd49} : s = 458;
	{8'd45,8'd50} : s = 500;
	{8'd45,8'd51} : s = 65;
	{8'd45,8'd52} : s = 200;
	{8'd45,8'd53} : s = 196;
	{8'd45,8'd54} : s = 353;
	{8'd45,8'd55} : s = 194;
	{8'd45,8'd56} : s = 344;
	{8'd45,8'd57} : s = 340;
	{8'd45,8'd58} : s = 457;
	{8'd45,8'd59} : s = 193;
	{8'd45,8'd60} : s = 338;
	{8'd45,8'd61} : s = 337;
	{8'd45,8'd62} : s = 454;
	{8'd45,8'd63} : s = 332;
	{8'd45,8'd64} : s = 453;
	{8'd45,8'd65} : s = 451;
	{8'd45,8'd66} : s = 498;
	{8'd45,8'd67} : s = 176;
	{8'd45,8'd68} : s = 330;
	{8'd45,8'd69} : s = 329;
	{8'd45,8'd70} : s = 440;
	{8'd45,8'd71} : s = 326;
	{8'd45,8'd72} : s = 436;
	{8'd45,8'd73} : s = 434;
	{8'd45,8'd74} : s = 497;
	{8'd45,8'd75} : s = 325;
	{8'd45,8'd76} : s = 433;
	{8'd45,8'd77} : s = 428;
	{8'd45,8'd78} : s = 492;
	{8'd45,8'd79} : s = 426;
	{8'd45,8'd80} : s = 490;
	{8'd45,8'd81} : s = 489;
	{8'd45,8'd82} : s = 508;
	{8'd45,8'd83} : s = 2;
	{8'd45,8'd84} : s = 48;
	{8'd45,8'd85} : s = 40;
	{8'd45,8'd86} : s = 168;
	{8'd45,8'd87} : s = 36;
	{8'd45,8'd88} : s = 164;
	{8'd45,8'd89} : s = 162;
	{8'd45,8'd90} : s = 323;
	{8'd45,8'd91} : s = 34;
	{8'd45,8'd92} : s = 161;
	{8'd45,8'd93} : s = 152;
	{8'd45,8'd94} : s = 312;
	{8'd45,8'd95} : s = 148;
	{8'd45,8'd96} : s = 308;
	{8'd45,8'd97} : s = 306;
	{8'd45,8'd98} : s = 425;
	{8'd45,8'd99} : s = 33;
	{8'd45,8'd100} : s = 146;
	{8'd45,8'd101} : s = 145;
	{8'd45,8'd102} : s = 305;
	{8'd45,8'd103} : s = 140;
	{8'd45,8'd104} : s = 300;
	{8'd45,8'd105} : s = 298;
	{8'd45,8'd106} : s = 422;
	{8'd45,8'd107} : s = 138;
	{8'd45,8'd108} : s = 297;
	{8'd45,8'd109} : s = 294;
	{8'd45,8'd110} : s = 421;
	{8'd45,8'd111} : s = 293;
	{8'd45,8'd112} : s = 419;
	{8'd45,8'd113} : s = 412;
	{8'd45,8'd114} : s = 486;
	{8'd45,8'd115} : s = 24;
	{8'd45,8'd116} : s = 137;
	{8'd45,8'd117} : s = 134;
	{8'd45,8'd118} : s = 291;
	{8'd45,8'd119} : s = 133;
	{8'd45,8'd120} : s = 284;
	{8'd45,8'd121} : s = 282;
	{8'd45,8'd122} : s = 410;
	{8'd45,8'd123} : s = 131;
	{8'd45,8'd124} : s = 281;
	{8'd45,8'd125} : s = 278;
	{8'd45,8'd126} : s = 409;
	{8'd45,8'd127} : s = 277;
	{8'd45,8'd128} : s = 406;
	{8'd45,8'd129} : s = 405;
	{8'd45,8'd130} : s = 485;
	{8'd45,8'd131} : s = 112;
	{8'd45,8'd132} : s = 275;
	{8'd45,8'd133} : s = 270;
	{8'd45,8'd134} : s = 403;
	{8'd45,8'd135} : s = 269;
	{8'd45,8'd136} : s = 398;
	{8'd45,8'd137} : s = 397;
	{8'd45,8'd138} : s = 483;
	{8'd45,8'd139} : s = 267;
	{8'd45,8'd140} : s = 395;
	{8'd45,8'd141} : s = 391;
	{8'd45,8'd142} : s = 476;
	{8'd45,8'd143} : s = 376;
	{8'd45,8'd144} : s = 474;
	{8'd45,8'd145} : s = 473;
	{8'd45,8'd146} : s = 506;
	{8'd45,8'd147} : s = 20;
	{8'd45,8'd148} : s = 104;
	{8'd45,8'd149} : s = 100;
	{8'd45,8'd150} : s = 263;
	{8'd45,8'd151} : s = 98;
	{8'd45,8'd152} : s = 240;
	{8'd45,8'd153} : s = 232;
	{8'd45,8'd154} : s = 372;
	{8'd45,8'd155} : s = 97;
	{8'd45,8'd156} : s = 228;
	{8'd45,8'd157} : s = 226;
	{8'd45,8'd158} : s = 370;
	{8'd45,8'd159} : s = 225;
	{8'd45,8'd160} : s = 369;
	{8'd45,8'd161} : s = 364;
	{8'd45,8'd162} : s = 470;
	{8'd45,8'd163} : s = 88;
	{8'd45,8'd164} : s = 216;
	{8'd45,8'd165} : s = 212;
	{8'd45,8'd166} : s = 362;
	{8'd45,8'd167} : s = 210;
	{8'd45,8'd168} : s = 361;
	{8'd45,8'd169} : s = 358;
	{8'd45,8'd170} : s = 469;
	{8'd45,8'd171} : s = 209;
	{8'd45,8'd172} : s = 357;
	{8'd45,8'd173} : s = 355;
	{8'd45,8'd174} : s = 467;
	{8'd45,8'd175} : s = 348;
	{8'd45,8'd176} : s = 462;
	{8'd45,8'd177} : s = 461;
	{8'd45,8'd178} : s = 505;
	{8'd45,8'd179} : s = 84;
	{8'd45,8'd180} : s = 204;
	{8'd45,8'd181} : s = 202;
	{8'd45,8'd182} : s = 346;
	{8'd45,8'd183} : s = 201;
	{8'd45,8'd184} : s = 345;
	{8'd45,8'd185} : s = 342;
	{8'd45,8'd186} : s = 459;
	{8'd45,8'd187} : s = 198;
	{8'd45,8'd188} : s = 341;
	{8'd45,8'd189} : s = 339;
	{8'd45,8'd190} : s = 455;
	{8'd45,8'd191} : s = 334;
	{8'd45,8'd192} : s = 444;
	{8'd45,8'd193} : s = 442;
	{8'd45,8'd194} : s = 502;
	{8'd45,8'd195} : s = 197;
	{8'd45,8'd196} : s = 333;
	{8'd45,8'd197} : s = 331;
	{8'd45,8'd198} : s = 441;
	{8'd45,8'd199} : s = 327;
	{8'd45,8'd200} : s = 438;
	{8'd45,8'd201} : s = 437;
	{8'd45,8'd202} : s = 501;
	{8'd45,8'd203} : s = 316;
	{8'd45,8'd204} : s = 435;
	{8'd45,8'd205} : s = 430;
	{8'd45,8'd206} : s = 499;
	{8'd45,8'd207} : s = 429;
	{8'd45,8'd208} : s = 494;
	{8'd45,8'd209} : s = 493;
	{8'd45,8'd210} : s = 510;
	{8'd45,8'd211} : s = 1;
	{8'd45,8'd212} : s = 18;
	{8'd45,8'd213} : s = 17;
	{8'd45,8'd214} : s = 82;
	{8'd45,8'd215} : s = 12;
	{8'd45,8'd216} : s = 81;
	{8'd45,8'd217} : s = 76;
	{8'd45,8'd218} : s = 195;
	{8'd45,8'd219} : s = 10;
	{8'd45,8'd220} : s = 74;
	{8'd45,8'd221} : s = 73;
	{8'd45,8'd222} : s = 184;
	{8'd45,8'd223} : s = 70;
	{8'd45,8'd224} : s = 180;
	{8'd45,8'd225} : s = 178;
	{8'd45,8'd226} : s = 314;
	{8'd45,8'd227} : s = 9;
	{8'd45,8'd228} : s = 69;
	{8'd45,8'd229} : s = 67;
	{8'd45,8'd230} : s = 177;
	{8'd45,8'd231} : s = 56;
	{8'd45,8'd232} : s = 172;
	{8'd45,8'd233} : s = 170;
	{8'd45,8'd234} : s = 313;
	{8'd45,8'd235} : s = 52;
	{8'd45,8'd236} : s = 169;
	{8'd45,8'd237} : s = 166;
	{8'd45,8'd238} : s = 310;
	{8'd45,8'd239} : s = 165;
	{8'd45,8'd240} : s = 309;
	{8'd45,8'd241} : s = 307;
	{8'd45,8'd242} : s = 427;
	{8'd45,8'd243} : s = 6;
	{8'd45,8'd244} : s = 50;
	{8'd45,8'd245} : s = 49;
	{8'd45,8'd246} : s = 163;
	{8'd45,8'd247} : s = 44;
	{8'd45,8'd248} : s = 156;
	{8'd45,8'd249} : s = 154;
	{8'd45,8'd250} : s = 302;
	{8'd45,8'd251} : s = 42;
	{8'd45,8'd252} : s = 153;
	{8'd45,8'd253} : s = 150;
	{8'd45,8'd254} : s = 301;
	{8'd45,8'd255} : s = 149;
	{8'd46,8'd0} : s = 420;
	{8'd46,8'd1} : s = 488;
	{8'd46,8'd2} : s = 129;
	{8'd46,8'd3} : s = 290;
	{8'd46,8'd4} : s = 289;
	{8'd46,8'd5} : s = 418;
	{8'd46,8'd6} : s = 280;
	{8'd46,8'd7} : s = 417;
	{8'd46,8'd8} : s = 408;
	{8'd46,8'd9} : s = 484;
	{8'd46,8'd10} : s = 276;
	{8'd46,8'd11} : s = 404;
	{8'd46,8'd12} : s = 402;
	{8'd46,8'd13} : s = 482;
	{8'd46,8'd14} : s = 401;
	{8'd46,8'd15} : s = 481;
	{8'd46,8'd16} : s = 472;
	{8'd46,8'd17} : s = 504;
	{8'd46,8'd18} : s = 4;
	{8'd46,8'd19} : s = 96;
	{8'd46,8'd20} : s = 80;
	{8'd46,8'd21} : s = 274;
	{8'd46,8'd22} : s = 72;
	{8'd46,8'd23} : s = 273;
	{8'd46,8'd24} : s = 268;
	{8'd46,8'd25} : s = 396;
	{8'd46,8'd26} : s = 68;
	{8'd46,8'd27} : s = 266;
	{8'd46,8'd28} : s = 265;
	{8'd46,8'd29} : s = 394;
	{8'd46,8'd30} : s = 262;
	{8'd46,8'd31} : s = 393;
	{8'd46,8'd32} : s = 390;
	{8'd46,8'd33} : s = 468;
	{8'd46,8'd34} : s = 66;
	{8'd46,8'd35} : s = 261;
	{8'd46,8'd36} : s = 259;
	{8'd46,8'd37} : s = 389;
	{8'd46,8'd38} : s = 224;
	{8'd46,8'd39} : s = 387;
	{8'd46,8'd40} : s = 368;
	{8'd46,8'd41} : s = 466;
	{8'd46,8'd42} : s = 208;
	{8'd46,8'd43} : s = 360;
	{8'd46,8'd44} : s = 356;
	{8'd46,8'd45} : s = 465;
	{8'd46,8'd46} : s = 354;
	{8'd46,8'd47} : s = 460;
	{8'd46,8'd48} : s = 458;
	{8'd46,8'd49} : s = 500;
	{8'd46,8'd50} : s = 65;
	{8'd46,8'd51} : s = 200;
	{8'd46,8'd52} : s = 196;
	{8'd46,8'd53} : s = 353;
	{8'd46,8'd54} : s = 194;
	{8'd46,8'd55} : s = 344;
	{8'd46,8'd56} : s = 340;
	{8'd46,8'd57} : s = 457;
	{8'd46,8'd58} : s = 193;
	{8'd46,8'd59} : s = 338;
	{8'd46,8'd60} : s = 337;
	{8'd46,8'd61} : s = 454;
	{8'd46,8'd62} : s = 332;
	{8'd46,8'd63} : s = 453;
	{8'd46,8'd64} : s = 451;
	{8'd46,8'd65} : s = 498;
	{8'd46,8'd66} : s = 176;
	{8'd46,8'd67} : s = 330;
	{8'd46,8'd68} : s = 329;
	{8'd46,8'd69} : s = 440;
	{8'd46,8'd70} : s = 326;
	{8'd46,8'd71} : s = 436;
	{8'd46,8'd72} : s = 434;
	{8'd46,8'd73} : s = 497;
	{8'd46,8'd74} : s = 325;
	{8'd46,8'd75} : s = 433;
	{8'd46,8'd76} : s = 428;
	{8'd46,8'd77} : s = 492;
	{8'd46,8'd78} : s = 426;
	{8'd46,8'd79} : s = 490;
	{8'd46,8'd80} : s = 489;
	{8'd46,8'd81} : s = 508;
	{8'd46,8'd82} : s = 2;
	{8'd46,8'd83} : s = 48;
	{8'd46,8'd84} : s = 40;
	{8'd46,8'd85} : s = 168;
	{8'd46,8'd86} : s = 36;
	{8'd46,8'd87} : s = 164;
	{8'd46,8'd88} : s = 162;
	{8'd46,8'd89} : s = 323;
	{8'd46,8'd90} : s = 34;
	{8'd46,8'd91} : s = 161;
	{8'd46,8'd92} : s = 152;
	{8'd46,8'd93} : s = 312;
	{8'd46,8'd94} : s = 148;
	{8'd46,8'd95} : s = 308;
	{8'd46,8'd96} : s = 306;
	{8'd46,8'd97} : s = 425;
	{8'd46,8'd98} : s = 33;
	{8'd46,8'd99} : s = 146;
	{8'd46,8'd100} : s = 145;
	{8'd46,8'd101} : s = 305;
	{8'd46,8'd102} : s = 140;
	{8'd46,8'd103} : s = 300;
	{8'd46,8'd104} : s = 298;
	{8'd46,8'd105} : s = 422;
	{8'd46,8'd106} : s = 138;
	{8'd46,8'd107} : s = 297;
	{8'd46,8'd108} : s = 294;
	{8'd46,8'd109} : s = 421;
	{8'd46,8'd110} : s = 293;
	{8'd46,8'd111} : s = 419;
	{8'd46,8'd112} : s = 412;
	{8'd46,8'd113} : s = 486;
	{8'd46,8'd114} : s = 24;
	{8'd46,8'd115} : s = 137;
	{8'd46,8'd116} : s = 134;
	{8'd46,8'd117} : s = 291;
	{8'd46,8'd118} : s = 133;
	{8'd46,8'd119} : s = 284;
	{8'd46,8'd120} : s = 282;
	{8'd46,8'd121} : s = 410;
	{8'd46,8'd122} : s = 131;
	{8'd46,8'd123} : s = 281;
	{8'd46,8'd124} : s = 278;
	{8'd46,8'd125} : s = 409;
	{8'd46,8'd126} : s = 277;
	{8'd46,8'd127} : s = 406;
	{8'd46,8'd128} : s = 405;
	{8'd46,8'd129} : s = 485;
	{8'd46,8'd130} : s = 112;
	{8'd46,8'd131} : s = 275;
	{8'd46,8'd132} : s = 270;
	{8'd46,8'd133} : s = 403;
	{8'd46,8'd134} : s = 269;
	{8'd46,8'd135} : s = 398;
	{8'd46,8'd136} : s = 397;
	{8'd46,8'd137} : s = 483;
	{8'd46,8'd138} : s = 267;
	{8'd46,8'd139} : s = 395;
	{8'd46,8'd140} : s = 391;
	{8'd46,8'd141} : s = 476;
	{8'd46,8'd142} : s = 376;
	{8'd46,8'd143} : s = 474;
	{8'd46,8'd144} : s = 473;
	{8'd46,8'd145} : s = 506;
	{8'd46,8'd146} : s = 20;
	{8'd46,8'd147} : s = 104;
	{8'd46,8'd148} : s = 100;
	{8'd46,8'd149} : s = 263;
	{8'd46,8'd150} : s = 98;
	{8'd46,8'd151} : s = 240;
	{8'd46,8'd152} : s = 232;
	{8'd46,8'd153} : s = 372;
	{8'd46,8'd154} : s = 97;
	{8'd46,8'd155} : s = 228;
	{8'd46,8'd156} : s = 226;
	{8'd46,8'd157} : s = 370;
	{8'd46,8'd158} : s = 225;
	{8'd46,8'd159} : s = 369;
	{8'd46,8'd160} : s = 364;
	{8'd46,8'd161} : s = 470;
	{8'd46,8'd162} : s = 88;
	{8'd46,8'd163} : s = 216;
	{8'd46,8'd164} : s = 212;
	{8'd46,8'd165} : s = 362;
	{8'd46,8'd166} : s = 210;
	{8'd46,8'd167} : s = 361;
	{8'd46,8'd168} : s = 358;
	{8'd46,8'd169} : s = 469;
	{8'd46,8'd170} : s = 209;
	{8'd46,8'd171} : s = 357;
	{8'd46,8'd172} : s = 355;
	{8'd46,8'd173} : s = 467;
	{8'd46,8'd174} : s = 348;
	{8'd46,8'd175} : s = 462;
	{8'd46,8'd176} : s = 461;
	{8'd46,8'd177} : s = 505;
	{8'd46,8'd178} : s = 84;
	{8'd46,8'd179} : s = 204;
	{8'd46,8'd180} : s = 202;
	{8'd46,8'd181} : s = 346;
	{8'd46,8'd182} : s = 201;
	{8'd46,8'd183} : s = 345;
	{8'd46,8'd184} : s = 342;
	{8'd46,8'd185} : s = 459;
	{8'd46,8'd186} : s = 198;
	{8'd46,8'd187} : s = 341;
	{8'd46,8'd188} : s = 339;
	{8'd46,8'd189} : s = 455;
	{8'd46,8'd190} : s = 334;
	{8'd46,8'd191} : s = 444;
	{8'd46,8'd192} : s = 442;
	{8'd46,8'd193} : s = 502;
	{8'd46,8'd194} : s = 197;
	{8'd46,8'd195} : s = 333;
	{8'd46,8'd196} : s = 331;
	{8'd46,8'd197} : s = 441;
	{8'd46,8'd198} : s = 327;
	{8'd46,8'd199} : s = 438;
	{8'd46,8'd200} : s = 437;
	{8'd46,8'd201} : s = 501;
	{8'd46,8'd202} : s = 316;
	{8'd46,8'd203} : s = 435;
	{8'd46,8'd204} : s = 430;
	{8'd46,8'd205} : s = 499;
	{8'd46,8'd206} : s = 429;
	{8'd46,8'd207} : s = 494;
	{8'd46,8'd208} : s = 493;
	{8'd46,8'd209} : s = 510;
	{8'd46,8'd210} : s = 1;
	{8'd46,8'd211} : s = 18;
	{8'd46,8'd212} : s = 17;
	{8'd46,8'd213} : s = 82;
	{8'd46,8'd214} : s = 12;
	{8'd46,8'd215} : s = 81;
	{8'd46,8'd216} : s = 76;
	{8'd46,8'd217} : s = 195;
	{8'd46,8'd218} : s = 10;
	{8'd46,8'd219} : s = 74;
	{8'd46,8'd220} : s = 73;
	{8'd46,8'd221} : s = 184;
	{8'd46,8'd222} : s = 70;
	{8'd46,8'd223} : s = 180;
	{8'd46,8'd224} : s = 178;
	{8'd46,8'd225} : s = 314;
	{8'd46,8'd226} : s = 9;
	{8'd46,8'd227} : s = 69;
	{8'd46,8'd228} : s = 67;
	{8'd46,8'd229} : s = 177;
	{8'd46,8'd230} : s = 56;
	{8'd46,8'd231} : s = 172;
	{8'd46,8'd232} : s = 170;
	{8'd46,8'd233} : s = 313;
	{8'd46,8'd234} : s = 52;
	{8'd46,8'd235} : s = 169;
	{8'd46,8'd236} : s = 166;
	{8'd46,8'd237} : s = 310;
	{8'd46,8'd238} : s = 165;
	{8'd46,8'd239} : s = 309;
	{8'd46,8'd240} : s = 307;
	{8'd46,8'd241} : s = 427;
	{8'd46,8'd242} : s = 6;
	{8'd46,8'd243} : s = 50;
	{8'd46,8'd244} : s = 49;
	{8'd46,8'd245} : s = 163;
	{8'd46,8'd246} : s = 44;
	{8'd46,8'd247} : s = 156;
	{8'd46,8'd248} : s = 154;
	{8'd46,8'd249} : s = 302;
	{8'd46,8'd250} : s = 42;
	{8'd46,8'd251} : s = 153;
	{8'd46,8'd252} : s = 150;
	{8'd46,8'd253} : s = 301;
	{8'd46,8'd254} : s = 149;
	{8'd46,8'd255} : s = 299;
	{8'd47,8'd0} : s = 488;
	{8'd47,8'd1} : s = 129;
	{8'd47,8'd2} : s = 290;
	{8'd47,8'd3} : s = 289;
	{8'd47,8'd4} : s = 418;
	{8'd47,8'd5} : s = 280;
	{8'd47,8'd6} : s = 417;
	{8'd47,8'd7} : s = 408;
	{8'd47,8'd8} : s = 484;
	{8'd47,8'd9} : s = 276;
	{8'd47,8'd10} : s = 404;
	{8'd47,8'd11} : s = 402;
	{8'd47,8'd12} : s = 482;
	{8'd47,8'd13} : s = 401;
	{8'd47,8'd14} : s = 481;
	{8'd47,8'd15} : s = 472;
	{8'd47,8'd16} : s = 504;
	{8'd47,8'd17} : s = 4;
	{8'd47,8'd18} : s = 96;
	{8'd47,8'd19} : s = 80;
	{8'd47,8'd20} : s = 274;
	{8'd47,8'd21} : s = 72;
	{8'd47,8'd22} : s = 273;
	{8'd47,8'd23} : s = 268;
	{8'd47,8'd24} : s = 396;
	{8'd47,8'd25} : s = 68;
	{8'd47,8'd26} : s = 266;
	{8'd47,8'd27} : s = 265;
	{8'd47,8'd28} : s = 394;
	{8'd47,8'd29} : s = 262;
	{8'd47,8'd30} : s = 393;
	{8'd47,8'd31} : s = 390;
	{8'd47,8'd32} : s = 468;
	{8'd47,8'd33} : s = 66;
	{8'd47,8'd34} : s = 261;
	{8'd47,8'd35} : s = 259;
	{8'd47,8'd36} : s = 389;
	{8'd47,8'd37} : s = 224;
	{8'd47,8'd38} : s = 387;
	{8'd47,8'd39} : s = 368;
	{8'd47,8'd40} : s = 466;
	{8'd47,8'd41} : s = 208;
	{8'd47,8'd42} : s = 360;
	{8'd47,8'd43} : s = 356;
	{8'd47,8'd44} : s = 465;
	{8'd47,8'd45} : s = 354;
	{8'd47,8'd46} : s = 460;
	{8'd47,8'd47} : s = 458;
	{8'd47,8'd48} : s = 500;
	{8'd47,8'd49} : s = 65;
	{8'd47,8'd50} : s = 200;
	{8'd47,8'd51} : s = 196;
	{8'd47,8'd52} : s = 353;
	{8'd47,8'd53} : s = 194;
	{8'd47,8'd54} : s = 344;
	{8'd47,8'd55} : s = 340;
	{8'd47,8'd56} : s = 457;
	{8'd47,8'd57} : s = 193;
	{8'd47,8'd58} : s = 338;
	{8'd47,8'd59} : s = 337;
	{8'd47,8'd60} : s = 454;
	{8'd47,8'd61} : s = 332;
	{8'd47,8'd62} : s = 453;
	{8'd47,8'd63} : s = 451;
	{8'd47,8'd64} : s = 498;
	{8'd47,8'd65} : s = 176;
	{8'd47,8'd66} : s = 330;
	{8'd47,8'd67} : s = 329;
	{8'd47,8'd68} : s = 440;
	{8'd47,8'd69} : s = 326;
	{8'd47,8'd70} : s = 436;
	{8'd47,8'd71} : s = 434;
	{8'd47,8'd72} : s = 497;
	{8'd47,8'd73} : s = 325;
	{8'd47,8'd74} : s = 433;
	{8'd47,8'd75} : s = 428;
	{8'd47,8'd76} : s = 492;
	{8'd47,8'd77} : s = 426;
	{8'd47,8'd78} : s = 490;
	{8'd47,8'd79} : s = 489;
	{8'd47,8'd80} : s = 508;
	{8'd47,8'd81} : s = 2;
	{8'd47,8'd82} : s = 48;
	{8'd47,8'd83} : s = 40;
	{8'd47,8'd84} : s = 168;
	{8'd47,8'd85} : s = 36;
	{8'd47,8'd86} : s = 164;
	{8'd47,8'd87} : s = 162;
	{8'd47,8'd88} : s = 323;
	{8'd47,8'd89} : s = 34;
	{8'd47,8'd90} : s = 161;
	{8'd47,8'd91} : s = 152;
	{8'd47,8'd92} : s = 312;
	{8'd47,8'd93} : s = 148;
	{8'd47,8'd94} : s = 308;
	{8'd47,8'd95} : s = 306;
	{8'd47,8'd96} : s = 425;
	{8'd47,8'd97} : s = 33;
	{8'd47,8'd98} : s = 146;
	{8'd47,8'd99} : s = 145;
	{8'd47,8'd100} : s = 305;
	{8'd47,8'd101} : s = 140;
	{8'd47,8'd102} : s = 300;
	{8'd47,8'd103} : s = 298;
	{8'd47,8'd104} : s = 422;
	{8'd47,8'd105} : s = 138;
	{8'd47,8'd106} : s = 297;
	{8'd47,8'd107} : s = 294;
	{8'd47,8'd108} : s = 421;
	{8'd47,8'd109} : s = 293;
	{8'd47,8'd110} : s = 419;
	{8'd47,8'd111} : s = 412;
	{8'd47,8'd112} : s = 486;
	{8'd47,8'd113} : s = 24;
	{8'd47,8'd114} : s = 137;
	{8'd47,8'd115} : s = 134;
	{8'd47,8'd116} : s = 291;
	{8'd47,8'd117} : s = 133;
	{8'd47,8'd118} : s = 284;
	{8'd47,8'd119} : s = 282;
	{8'd47,8'd120} : s = 410;
	{8'd47,8'd121} : s = 131;
	{8'd47,8'd122} : s = 281;
	{8'd47,8'd123} : s = 278;
	{8'd47,8'd124} : s = 409;
	{8'd47,8'd125} : s = 277;
	{8'd47,8'd126} : s = 406;
	{8'd47,8'd127} : s = 405;
	{8'd47,8'd128} : s = 485;
	{8'd47,8'd129} : s = 112;
	{8'd47,8'd130} : s = 275;
	{8'd47,8'd131} : s = 270;
	{8'd47,8'd132} : s = 403;
	{8'd47,8'd133} : s = 269;
	{8'd47,8'd134} : s = 398;
	{8'd47,8'd135} : s = 397;
	{8'd47,8'd136} : s = 483;
	{8'd47,8'd137} : s = 267;
	{8'd47,8'd138} : s = 395;
	{8'd47,8'd139} : s = 391;
	{8'd47,8'd140} : s = 476;
	{8'd47,8'd141} : s = 376;
	{8'd47,8'd142} : s = 474;
	{8'd47,8'd143} : s = 473;
	{8'd47,8'd144} : s = 506;
	{8'd47,8'd145} : s = 20;
	{8'd47,8'd146} : s = 104;
	{8'd47,8'd147} : s = 100;
	{8'd47,8'd148} : s = 263;
	{8'd47,8'd149} : s = 98;
	{8'd47,8'd150} : s = 240;
	{8'd47,8'd151} : s = 232;
	{8'd47,8'd152} : s = 372;
	{8'd47,8'd153} : s = 97;
	{8'd47,8'd154} : s = 228;
	{8'd47,8'd155} : s = 226;
	{8'd47,8'd156} : s = 370;
	{8'd47,8'd157} : s = 225;
	{8'd47,8'd158} : s = 369;
	{8'd47,8'd159} : s = 364;
	{8'd47,8'd160} : s = 470;
	{8'd47,8'd161} : s = 88;
	{8'd47,8'd162} : s = 216;
	{8'd47,8'd163} : s = 212;
	{8'd47,8'd164} : s = 362;
	{8'd47,8'd165} : s = 210;
	{8'd47,8'd166} : s = 361;
	{8'd47,8'd167} : s = 358;
	{8'd47,8'd168} : s = 469;
	{8'd47,8'd169} : s = 209;
	{8'd47,8'd170} : s = 357;
	{8'd47,8'd171} : s = 355;
	{8'd47,8'd172} : s = 467;
	{8'd47,8'd173} : s = 348;
	{8'd47,8'd174} : s = 462;
	{8'd47,8'd175} : s = 461;
	{8'd47,8'd176} : s = 505;
	{8'd47,8'd177} : s = 84;
	{8'd47,8'd178} : s = 204;
	{8'd47,8'd179} : s = 202;
	{8'd47,8'd180} : s = 346;
	{8'd47,8'd181} : s = 201;
	{8'd47,8'd182} : s = 345;
	{8'd47,8'd183} : s = 342;
	{8'd47,8'd184} : s = 459;
	{8'd47,8'd185} : s = 198;
	{8'd47,8'd186} : s = 341;
	{8'd47,8'd187} : s = 339;
	{8'd47,8'd188} : s = 455;
	{8'd47,8'd189} : s = 334;
	{8'd47,8'd190} : s = 444;
	{8'd47,8'd191} : s = 442;
	{8'd47,8'd192} : s = 502;
	{8'd47,8'd193} : s = 197;
	{8'd47,8'd194} : s = 333;
	{8'd47,8'd195} : s = 331;
	{8'd47,8'd196} : s = 441;
	{8'd47,8'd197} : s = 327;
	{8'd47,8'd198} : s = 438;
	{8'd47,8'd199} : s = 437;
	{8'd47,8'd200} : s = 501;
	{8'd47,8'd201} : s = 316;
	{8'd47,8'd202} : s = 435;
	{8'd47,8'd203} : s = 430;
	{8'd47,8'd204} : s = 499;
	{8'd47,8'd205} : s = 429;
	{8'd47,8'd206} : s = 494;
	{8'd47,8'd207} : s = 493;
	{8'd47,8'd208} : s = 510;
	{8'd47,8'd209} : s = 1;
	{8'd47,8'd210} : s = 18;
	{8'd47,8'd211} : s = 17;
	{8'd47,8'd212} : s = 82;
	{8'd47,8'd213} : s = 12;
	{8'd47,8'd214} : s = 81;
	{8'd47,8'd215} : s = 76;
	{8'd47,8'd216} : s = 195;
	{8'd47,8'd217} : s = 10;
	{8'd47,8'd218} : s = 74;
	{8'd47,8'd219} : s = 73;
	{8'd47,8'd220} : s = 184;
	{8'd47,8'd221} : s = 70;
	{8'd47,8'd222} : s = 180;
	{8'd47,8'd223} : s = 178;
	{8'd47,8'd224} : s = 314;
	{8'd47,8'd225} : s = 9;
	{8'd47,8'd226} : s = 69;
	{8'd47,8'd227} : s = 67;
	{8'd47,8'd228} : s = 177;
	{8'd47,8'd229} : s = 56;
	{8'd47,8'd230} : s = 172;
	{8'd47,8'd231} : s = 170;
	{8'd47,8'd232} : s = 313;
	{8'd47,8'd233} : s = 52;
	{8'd47,8'd234} : s = 169;
	{8'd47,8'd235} : s = 166;
	{8'd47,8'd236} : s = 310;
	{8'd47,8'd237} : s = 165;
	{8'd47,8'd238} : s = 309;
	{8'd47,8'd239} : s = 307;
	{8'd47,8'd240} : s = 427;
	{8'd47,8'd241} : s = 6;
	{8'd47,8'd242} : s = 50;
	{8'd47,8'd243} : s = 49;
	{8'd47,8'd244} : s = 163;
	{8'd47,8'd245} : s = 44;
	{8'd47,8'd246} : s = 156;
	{8'd47,8'd247} : s = 154;
	{8'd47,8'd248} : s = 302;
	{8'd47,8'd249} : s = 42;
	{8'd47,8'd250} : s = 153;
	{8'd47,8'd251} : s = 150;
	{8'd47,8'd252} : s = 301;
	{8'd47,8'd253} : s = 149;
	{8'd47,8'd254} : s = 299;
	{8'd47,8'd255} : s = 295;
	{8'd48,8'd0} : s = 129;
	{8'd48,8'd1} : s = 290;
	{8'd48,8'd2} : s = 289;
	{8'd48,8'd3} : s = 418;
	{8'd48,8'd4} : s = 280;
	{8'd48,8'd5} : s = 417;
	{8'd48,8'd6} : s = 408;
	{8'd48,8'd7} : s = 484;
	{8'd48,8'd8} : s = 276;
	{8'd48,8'd9} : s = 404;
	{8'd48,8'd10} : s = 402;
	{8'd48,8'd11} : s = 482;
	{8'd48,8'd12} : s = 401;
	{8'd48,8'd13} : s = 481;
	{8'd48,8'd14} : s = 472;
	{8'd48,8'd15} : s = 504;
	{8'd48,8'd16} : s = 4;
	{8'd48,8'd17} : s = 96;
	{8'd48,8'd18} : s = 80;
	{8'd48,8'd19} : s = 274;
	{8'd48,8'd20} : s = 72;
	{8'd48,8'd21} : s = 273;
	{8'd48,8'd22} : s = 268;
	{8'd48,8'd23} : s = 396;
	{8'd48,8'd24} : s = 68;
	{8'd48,8'd25} : s = 266;
	{8'd48,8'd26} : s = 265;
	{8'd48,8'd27} : s = 394;
	{8'd48,8'd28} : s = 262;
	{8'd48,8'd29} : s = 393;
	{8'd48,8'd30} : s = 390;
	{8'd48,8'd31} : s = 468;
	{8'd48,8'd32} : s = 66;
	{8'd48,8'd33} : s = 261;
	{8'd48,8'd34} : s = 259;
	{8'd48,8'd35} : s = 389;
	{8'd48,8'd36} : s = 224;
	{8'd48,8'd37} : s = 387;
	{8'd48,8'd38} : s = 368;
	{8'd48,8'd39} : s = 466;
	{8'd48,8'd40} : s = 208;
	{8'd48,8'd41} : s = 360;
	{8'd48,8'd42} : s = 356;
	{8'd48,8'd43} : s = 465;
	{8'd48,8'd44} : s = 354;
	{8'd48,8'd45} : s = 460;
	{8'd48,8'd46} : s = 458;
	{8'd48,8'd47} : s = 500;
	{8'd48,8'd48} : s = 65;
	{8'd48,8'd49} : s = 200;
	{8'd48,8'd50} : s = 196;
	{8'd48,8'd51} : s = 353;
	{8'd48,8'd52} : s = 194;
	{8'd48,8'd53} : s = 344;
	{8'd48,8'd54} : s = 340;
	{8'd48,8'd55} : s = 457;
	{8'd48,8'd56} : s = 193;
	{8'd48,8'd57} : s = 338;
	{8'd48,8'd58} : s = 337;
	{8'd48,8'd59} : s = 454;
	{8'd48,8'd60} : s = 332;
	{8'd48,8'd61} : s = 453;
	{8'd48,8'd62} : s = 451;
	{8'd48,8'd63} : s = 498;
	{8'd48,8'd64} : s = 176;
	{8'd48,8'd65} : s = 330;
	{8'd48,8'd66} : s = 329;
	{8'd48,8'd67} : s = 440;
	{8'd48,8'd68} : s = 326;
	{8'd48,8'd69} : s = 436;
	{8'd48,8'd70} : s = 434;
	{8'd48,8'd71} : s = 497;
	{8'd48,8'd72} : s = 325;
	{8'd48,8'd73} : s = 433;
	{8'd48,8'd74} : s = 428;
	{8'd48,8'd75} : s = 492;
	{8'd48,8'd76} : s = 426;
	{8'd48,8'd77} : s = 490;
	{8'd48,8'd78} : s = 489;
	{8'd48,8'd79} : s = 508;
	{8'd48,8'd80} : s = 2;
	{8'd48,8'd81} : s = 48;
	{8'd48,8'd82} : s = 40;
	{8'd48,8'd83} : s = 168;
	{8'd48,8'd84} : s = 36;
	{8'd48,8'd85} : s = 164;
	{8'd48,8'd86} : s = 162;
	{8'd48,8'd87} : s = 323;
	{8'd48,8'd88} : s = 34;
	{8'd48,8'd89} : s = 161;
	{8'd48,8'd90} : s = 152;
	{8'd48,8'd91} : s = 312;
	{8'd48,8'd92} : s = 148;
	{8'd48,8'd93} : s = 308;
	{8'd48,8'd94} : s = 306;
	{8'd48,8'd95} : s = 425;
	{8'd48,8'd96} : s = 33;
	{8'd48,8'd97} : s = 146;
	{8'd48,8'd98} : s = 145;
	{8'd48,8'd99} : s = 305;
	{8'd48,8'd100} : s = 140;
	{8'd48,8'd101} : s = 300;
	{8'd48,8'd102} : s = 298;
	{8'd48,8'd103} : s = 422;
	{8'd48,8'd104} : s = 138;
	{8'd48,8'd105} : s = 297;
	{8'd48,8'd106} : s = 294;
	{8'd48,8'd107} : s = 421;
	{8'd48,8'd108} : s = 293;
	{8'd48,8'd109} : s = 419;
	{8'd48,8'd110} : s = 412;
	{8'd48,8'd111} : s = 486;
	{8'd48,8'd112} : s = 24;
	{8'd48,8'd113} : s = 137;
	{8'd48,8'd114} : s = 134;
	{8'd48,8'd115} : s = 291;
	{8'd48,8'd116} : s = 133;
	{8'd48,8'd117} : s = 284;
	{8'd48,8'd118} : s = 282;
	{8'd48,8'd119} : s = 410;
	{8'd48,8'd120} : s = 131;
	{8'd48,8'd121} : s = 281;
	{8'd48,8'd122} : s = 278;
	{8'd48,8'd123} : s = 409;
	{8'd48,8'd124} : s = 277;
	{8'd48,8'd125} : s = 406;
	{8'd48,8'd126} : s = 405;
	{8'd48,8'd127} : s = 485;
	{8'd48,8'd128} : s = 112;
	{8'd48,8'd129} : s = 275;
	{8'd48,8'd130} : s = 270;
	{8'd48,8'd131} : s = 403;
	{8'd48,8'd132} : s = 269;
	{8'd48,8'd133} : s = 398;
	{8'd48,8'd134} : s = 397;
	{8'd48,8'd135} : s = 483;
	{8'd48,8'd136} : s = 267;
	{8'd48,8'd137} : s = 395;
	{8'd48,8'd138} : s = 391;
	{8'd48,8'd139} : s = 476;
	{8'd48,8'd140} : s = 376;
	{8'd48,8'd141} : s = 474;
	{8'd48,8'd142} : s = 473;
	{8'd48,8'd143} : s = 506;
	{8'd48,8'd144} : s = 20;
	{8'd48,8'd145} : s = 104;
	{8'd48,8'd146} : s = 100;
	{8'd48,8'd147} : s = 263;
	{8'd48,8'd148} : s = 98;
	{8'd48,8'd149} : s = 240;
	{8'd48,8'd150} : s = 232;
	{8'd48,8'd151} : s = 372;
	{8'd48,8'd152} : s = 97;
	{8'd48,8'd153} : s = 228;
	{8'd48,8'd154} : s = 226;
	{8'd48,8'd155} : s = 370;
	{8'd48,8'd156} : s = 225;
	{8'd48,8'd157} : s = 369;
	{8'd48,8'd158} : s = 364;
	{8'd48,8'd159} : s = 470;
	{8'd48,8'd160} : s = 88;
	{8'd48,8'd161} : s = 216;
	{8'd48,8'd162} : s = 212;
	{8'd48,8'd163} : s = 362;
	{8'd48,8'd164} : s = 210;
	{8'd48,8'd165} : s = 361;
	{8'd48,8'd166} : s = 358;
	{8'd48,8'd167} : s = 469;
	{8'd48,8'd168} : s = 209;
	{8'd48,8'd169} : s = 357;
	{8'd48,8'd170} : s = 355;
	{8'd48,8'd171} : s = 467;
	{8'd48,8'd172} : s = 348;
	{8'd48,8'd173} : s = 462;
	{8'd48,8'd174} : s = 461;
	{8'd48,8'd175} : s = 505;
	{8'd48,8'd176} : s = 84;
	{8'd48,8'd177} : s = 204;
	{8'd48,8'd178} : s = 202;
	{8'd48,8'd179} : s = 346;
	{8'd48,8'd180} : s = 201;
	{8'd48,8'd181} : s = 345;
	{8'd48,8'd182} : s = 342;
	{8'd48,8'd183} : s = 459;
	{8'd48,8'd184} : s = 198;
	{8'd48,8'd185} : s = 341;
	{8'd48,8'd186} : s = 339;
	{8'd48,8'd187} : s = 455;
	{8'd48,8'd188} : s = 334;
	{8'd48,8'd189} : s = 444;
	{8'd48,8'd190} : s = 442;
	{8'd48,8'd191} : s = 502;
	{8'd48,8'd192} : s = 197;
	{8'd48,8'd193} : s = 333;
	{8'd48,8'd194} : s = 331;
	{8'd48,8'd195} : s = 441;
	{8'd48,8'd196} : s = 327;
	{8'd48,8'd197} : s = 438;
	{8'd48,8'd198} : s = 437;
	{8'd48,8'd199} : s = 501;
	{8'd48,8'd200} : s = 316;
	{8'd48,8'd201} : s = 435;
	{8'd48,8'd202} : s = 430;
	{8'd48,8'd203} : s = 499;
	{8'd48,8'd204} : s = 429;
	{8'd48,8'd205} : s = 494;
	{8'd48,8'd206} : s = 493;
	{8'd48,8'd207} : s = 510;
	{8'd48,8'd208} : s = 1;
	{8'd48,8'd209} : s = 18;
	{8'd48,8'd210} : s = 17;
	{8'd48,8'd211} : s = 82;
	{8'd48,8'd212} : s = 12;
	{8'd48,8'd213} : s = 81;
	{8'd48,8'd214} : s = 76;
	{8'd48,8'd215} : s = 195;
	{8'd48,8'd216} : s = 10;
	{8'd48,8'd217} : s = 74;
	{8'd48,8'd218} : s = 73;
	{8'd48,8'd219} : s = 184;
	{8'd48,8'd220} : s = 70;
	{8'd48,8'd221} : s = 180;
	{8'd48,8'd222} : s = 178;
	{8'd48,8'd223} : s = 314;
	{8'd48,8'd224} : s = 9;
	{8'd48,8'd225} : s = 69;
	{8'd48,8'd226} : s = 67;
	{8'd48,8'd227} : s = 177;
	{8'd48,8'd228} : s = 56;
	{8'd48,8'd229} : s = 172;
	{8'd48,8'd230} : s = 170;
	{8'd48,8'd231} : s = 313;
	{8'd48,8'd232} : s = 52;
	{8'd48,8'd233} : s = 169;
	{8'd48,8'd234} : s = 166;
	{8'd48,8'd235} : s = 310;
	{8'd48,8'd236} : s = 165;
	{8'd48,8'd237} : s = 309;
	{8'd48,8'd238} : s = 307;
	{8'd48,8'd239} : s = 427;
	{8'd48,8'd240} : s = 6;
	{8'd48,8'd241} : s = 50;
	{8'd48,8'd242} : s = 49;
	{8'd48,8'd243} : s = 163;
	{8'd48,8'd244} : s = 44;
	{8'd48,8'd245} : s = 156;
	{8'd48,8'd246} : s = 154;
	{8'd48,8'd247} : s = 302;
	{8'd48,8'd248} : s = 42;
	{8'd48,8'd249} : s = 153;
	{8'd48,8'd250} : s = 150;
	{8'd48,8'd251} : s = 301;
	{8'd48,8'd252} : s = 149;
	{8'd48,8'd253} : s = 299;
	{8'd48,8'd254} : s = 295;
	{8'd48,8'd255} : s = 423;
	{8'd49,8'd0} : s = 290;
	{8'd49,8'd1} : s = 289;
	{8'd49,8'd2} : s = 418;
	{8'd49,8'd3} : s = 280;
	{8'd49,8'd4} : s = 417;
	{8'd49,8'd5} : s = 408;
	{8'd49,8'd6} : s = 484;
	{8'd49,8'd7} : s = 276;
	{8'd49,8'd8} : s = 404;
	{8'd49,8'd9} : s = 402;
	{8'd49,8'd10} : s = 482;
	{8'd49,8'd11} : s = 401;
	{8'd49,8'd12} : s = 481;
	{8'd49,8'd13} : s = 472;
	{8'd49,8'd14} : s = 504;
	{8'd49,8'd15} : s = 4;
	{8'd49,8'd16} : s = 96;
	{8'd49,8'd17} : s = 80;
	{8'd49,8'd18} : s = 274;
	{8'd49,8'd19} : s = 72;
	{8'd49,8'd20} : s = 273;
	{8'd49,8'd21} : s = 268;
	{8'd49,8'd22} : s = 396;
	{8'd49,8'd23} : s = 68;
	{8'd49,8'd24} : s = 266;
	{8'd49,8'd25} : s = 265;
	{8'd49,8'd26} : s = 394;
	{8'd49,8'd27} : s = 262;
	{8'd49,8'd28} : s = 393;
	{8'd49,8'd29} : s = 390;
	{8'd49,8'd30} : s = 468;
	{8'd49,8'd31} : s = 66;
	{8'd49,8'd32} : s = 261;
	{8'd49,8'd33} : s = 259;
	{8'd49,8'd34} : s = 389;
	{8'd49,8'd35} : s = 224;
	{8'd49,8'd36} : s = 387;
	{8'd49,8'd37} : s = 368;
	{8'd49,8'd38} : s = 466;
	{8'd49,8'd39} : s = 208;
	{8'd49,8'd40} : s = 360;
	{8'd49,8'd41} : s = 356;
	{8'd49,8'd42} : s = 465;
	{8'd49,8'd43} : s = 354;
	{8'd49,8'd44} : s = 460;
	{8'd49,8'd45} : s = 458;
	{8'd49,8'd46} : s = 500;
	{8'd49,8'd47} : s = 65;
	{8'd49,8'd48} : s = 200;
	{8'd49,8'd49} : s = 196;
	{8'd49,8'd50} : s = 353;
	{8'd49,8'd51} : s = 194;
	{8'd49,8'd52} : s = 344;
	{8'd49,8'd53} : s = 340;
	{8'd49,8'd54} : s = 457;
	{8'd49,8'd55} : s = 193;
	{8'd49,8'd56} : s = 338;
	{8'd49,8'd57} : s = 337;
	{8'd49,8'd58} : s = 454;
	{8'd49,8'd59} : s = 332;
	{8'd49,8'd60} : s = 453;
	{8'd49,8'd61} : s = 451;
	{8'd49,8'd62} : s = 498;
	{8'd49,8'd63} : s = 176;
	{8'd49,8'd64} : s = 330;
	{8'd49,8'd65} : s = 329;
	{8'd49,8'd66} : s = 440;
	{8'd49,8'd67} : s = 326;
	{8'd49,8'd68} : s = 436;
	{8'd49,8'd69} : s = 434;
	{8'd49,8'd70} : s = 497;
	{8'd49,8'd71} : s = 325;
	{8'd49,8'd72} : s = 433;
	{8'd49,8'd73} : s = 428;
	{8'd49,8'd74} : s = 492;
	{8'd49,8'd75} : s = 426;
	{8'd49,8'd76} : s = 490;
	{8'd49,8'd77} : s = 489;
	{8'd49,8'd78} : s = 508;
	{8'd49,8'd79} : s = 2;
	{8'd49,8'd80} : s = 48;
	{8'd49,8'd81} : s = 40;
	{8'd49,8'd82} : s = 168;
	{8'd49,8'd83} : s = 36;
	{8'd49,8'd84} : s = 164;
	{8'd49,8'd85} : s = 162;
	{8'd49,8'd86} : s = 323;
	{8'd49,8'd87} : s = 34;
	{8'd49,8'd88} : s = 161;
	{8'd49,8'd89} : s = 152;
	{8'd49,8'd90} : s = 312;
	{8'd49,8'd91} : s = 148;
	{8'd49,8'd92} : s = 308;
	{8'd49,8'd93} : s = 306;
	{8'd49,8'd94} : s = 425;
	{8'd49,8'd95} : s = 33;
	{8'd49,8'd96} : s = 146;
	{8'd49,8'd97} : s = 145;
	{8'd49,8'd98} : s = 305;
	{8'd49,8'd99} : s = 140;
	{8'd49,8'd100} : s = 300;
	{8'd49,8'd101} : s = 298;
	{8'd49,8'd102} : s = 422;
	{8'd49,8'd103} : s = 138;
	{8'd49,8'd104} : s = 297;
	{8'd49,8'd105} : s = 294;
	{8'd49,8'd106} : s = 421;
	{8'd49,8'd107} : s = 293;
	{8'd49,8'd108} : s = 419;
	{8'd49,8'd109} : s = 412;
	{8'd49,8'd110} : s = 486;
	{8'd49,8'd111} : s = 24;
	{8'd49,8'd112} : s = 137;
	{8'd49,8'd113} : s = 134;
	{8'd49,8'd114} : s = 291;
	{8'd49,8'd115} : s = 133;
	{8'd49,8'd116} : s = 284;
	{8'd49,8'd117} : s = 282;
	{8'd49,8'd118} : s = 410;
	{8'd49,8'd119} : s = 131;
	{8'd49,8'd120} : s = 281;
	{8'd49,8'd121} : s = 278;
	{8'd49,8'd122} : s = 409;
	{8'd49,8'd123} : s = 277;
	{8'd49,8'd124} : s = 406;
	{8'd49,8'd125} : s = 405;
	{8'd49,8'd126} : s = 485;
	{8'd49,8'd127} : s = 112;
	{8'd49,8'd128} : s = 275;
	{8'd49,8'd129} : s = 270;
	{8'd49,8'd130} : s = 403;
	{8'd49,8'd131} : s = 269;
	{8'd49,8'd132} : s = 398;
	{8'd49,8'd133} : s = 397;
	{8'd49,8'd134} : s = 483;
	{8'd49,8'd135} : s = 267;
	{8'd49,8'd136} : s = 395;
	{8'd49,8'd137} : s = 391;
	{8'd49,8'd138} : s = 476;
	{8'd49,8'd139} : s = 376;
	{8'd49,8'd140} : s = 474;
	{8'd49,8'd141} : s = 473;
	{8'd49,8'd142} : s = 506;
	{8'd49,8'd143} : s = 20;
	{8'd49,8'd144} : s = 104;
	{8'd49,8'd145} : s = 100;
	{8'd49,8'd146} : s = 263;
	{8'd49,8'd147} : s = 98;
	{8'd49,8'd148} : s = 240;
	{8'd49,8'd149} : s = 232;
	{8'd49,8'd150} : s = 372;
	{8'd49,8'd151} : s = 97;
	{8'd49,8'd152} : s = 228;
	{8'd49,8'd153} : s = 226;
	{8'd49,8'd154} : s = 370;
	{8'd49,8'd155} : s = 225;
	{8'd49,8'd156} : s = 369;
	{8'd49,8'd157} : s = 364;
	{8'd49,8'd158} : s = 470;
	{8'd49,8'd159} : s = 88;
	{8'd49,8'd160} : s = 216;
	{8'd49,8'd161} : s = 212;
	{8'd49,8'd162} : s = 362;
	{8'd49,8'd163} : s = 210;
	{8'd49,8'd164} : s = 361;
	{8'd49,8'd165} : s = 358;
	{8'd49,8'd166} : s = 469;
	{8'd49,8'd167} : s = 209;
	{8'd49,8'd168} : s = 357;
	{8'd49,8'd169} : s = 355;
	{8'd49,8'd170} : s = 467;
	{8'd49,8'd171} : s = 348;
	{8'd49,8'd172} : s = 462;
	{8'd49,8'd173} : s = 461;
	{8'd49,8'd174} : s = 505;
	{8'd49,8'd175} : s = 84;
	{8'd49,8'd176} : s = 204;
	{8'd49,8'd177} : s = 202;
	{8'd49,8'd178} : s = 346;
	{8'd49,8'd179} : s = 201;
	{8'd49,8'd180} : s = 345;
	{8'd49,8'd181} : s = 342;
	{8'd49,8'd182} : s = 459;
	{8'd49,8'd183} : s = 198;
	{8'd49,8'd184} : s = 341;
	{8'd49,8'd185} : s = 339;
	{8'd49,8'd186} : s = 455;
	{8'd49,8'd187} : s = 334;
	{8'd49,8'd188} : s = 444;
	{8'd49,8'd189} : s = 442;
	{8'd49,8'd190} : s = 502;
	{8'd49,8'd191} : s = 197;
	{8'd49,8'd192} : s = 333;
	{8'd49,8'd193} : s = 331;
	{8'd49,8'd194} : s = 441;
	{8'd49,8'd195} : s = 327;
	{8'd49,8'd196} : s = 438;
	{8'd49,8'd197} : s = 437;
	{8'd49,8'd198} : s = 501;
	{8'd49,8'd199} : s = 316;
	{8'd49,8'd200} : s = 435;
	{8'd49,8'd201} : s = 430;
	{8'd49,8'd202} : s = 499;
	{8'd49,8'd203} : s = 429;
	{8'd49,8'd204} : s = 494;
	{8'd49,8'd205} : s = 493;
	{8'd49,8'd206} : s = 510;
	{8'd49,8'd207} : s = 1;
	{8'd49,8'd208} : s = 18;
	{8'd49,8'd209} : s = 17;
	{8'd49,8'd210} : s = 82;
	{8'd49,8'd211} : s = 12;
	{8'd49,8'd212} : s = 81;
	{8'd49,8'd213} : s = 76;
	{8'd49,8'd214} : s = 195;
	{8'd49,8'd215} : s = 10;
	{8'd49,8'd216} : s = 74;
	{8'd49,8'd217} : s = 73;
	{8'd49,8'd218} : s = 184;
	{8'd49,8'd219} : s = 70;
	{8'd49,8'd220} : s = 180;
	{8'd49,8'd221} : s = 178;
	{8'd49,8'd222} : s = 314;
	{8'd49,8'd223} : s = 9;
	{8'd49,8'd224} : s = 69;
	{8'd49,8'd225} : s = 67;
	{8'd49,8'd226} : s = 177;
	{8'd49,8'd227} : s = 56;
	{8'd49,8'd228} : s = 172;
	{8'd49,8'd229} : s = 170;
	{8'd49,8'd230} : s = 313;
	{8'd49,8'd231} : s = 52;
	{8'd49,8'd232} : s = 169;
	{8'd49,8'd233} : s = 166;
	{8'd49,8'd234} : s = 310;
	{8'd49,8'd235} : s = 165;
	{8'd49,8'd236} : s = 309;
	{8'd49,8'd237} : s = 307;
	{8'd49,8'd238} : s = 427;
	{8'd49,8'd239} : s = 6;
	{8'd49,8'd240} : s = 50;
	{8'd49,8'd241} : s = 49;
	{8'd49,8'd242} : s = 163;
	{8'd49,8'd243} : s = 44;
	{8'd49,8'd244} : s = 156;
	{8'd49,8'd245} : s = 154;
	{8'd49,8'd246} : s = 302;
	{8'd49,8'd247} : s = 42;
	{8'd49,8'd248} : s = 153;
	{8'd49,8'd249} : s = 150;
	{8'd49,8'd250} : s = 301;
	{8'd49,8'd251} : s = 149;
	{8'd49,8'd252} : s = 299;
	{8'd49,8'd253} : s = 295;
	{8'd49,8'd254} : s = 423;
	{8'd49,8'd255} : s = 41;
	{8'd50,8'd0} : s = 289;
	{8'd50,8'd1} : s = 418;
	{8'd50,8'd2} : s = 280;
	{8'd50,8'd3} : s = 417;
	{8'd50,8'd4} : s = 408;
	{8'd50,8'd5} : s = 484;
	{8'd50,8'd6} : s = 276;
	{8'd50,8'd7} : s = 404;
	{8'd50,8'd8} : s = 402;
	{8'd50,8'd9} : s = 482;
	{8'd50,8'd10} : s = 401;
	{8'd50,8'd11} : s = 481;
	{8'd50,8'd12} : s = 472;
	{8'd50,8'd13} : s = 504;
	{8'd50,8'd14} : s = 4;
	{8'd50,8'd15} : s = 96;
	{8'd50,8'd16} : s = 80;
	{8'd50,8'd17} : s = 274;
	{8'd50,8'd18} : s = 72;
	{8'd50,8'd19} : s = 273;
	{8'd50,8'd20} : s = 268;
	{8'd50,8'd21} : s = 396;
	{8'd50,8'd22} : s = 68;
	{8'd50,8'd23} : s = 266;
	{8'd50,8'd24} : s = 265;
	{8'd50,8'd25} : s = 394;
	{8'd50,8'd26} : s = 262;
	{8'd50,8'd27} : s = 393;
	{8'd50,8'd28} : s = 390;
	{8'd50,8'd29} : s = 468;
	{8'd50,8'd30} : s = 66;
	{8'd50,8'd31} : s = 261;
	{8'd50,8'd32} : s = 259;
	{8'd50,8'd33} : s = 389;
	{8'd50,8'd34} : s = 224;
	{8'd50,8'd35} : s = 387;
	{8'd50,8'd36} : s = 368;
	{8'd50,8'd37} : s = 466;
	{8'd50,8'd38} : s = 208;
	{8'd50,8'd39} : s = 360;
	{8'd50,8'd40} : s = 356;
	{8'd50,8'd41} : s = 465;
	{8'd50,8'd42} : s = 354;
	{8'd50,8'd43} : s = 460;
	{8'd50,8'd44} : s = 458;
	{8'd50,8'd45} : s = 500;
	{8'd50,8'd46} : s = 65;
	{8'd50,8'd47} : s = 200;
	{8'd50,8'd48} : s = 196;
	{8'd50,8'd49} : s = 353;
	{8'd50,8'd50} : s = 194;
	{8'd50,8'd51} : s = 344;
	{8'd50,8'd52} : s = 340;
	{8'd50,8'd53} : s = 457;
	{8'd50,8'd54} : s = 193;
	{8'd50,8'd55} : s = 338;
	{8'd50,8'd56} : s = 337;
	{8'd50,8'd57} : s = 454;
	{8'd50,8'd58} : s = 332;
	{8'd50,8'd59} : s = 453;
	{8'd50,8'd60} : s = 451;
	{8'd50,8'd61} : s = 498;
	{8'd50,8'd62} : s = 176;
	{8'd50,8'd63} : s = 330;
	{8'd50,8'd64} : s = 329;
	{8'd50,8'd65} : s = 440;
	{8'd50,8'd66} : s = 326;
	{8'd50,8'd67} : s = 436;
	{8'd50,8'd68} : s = 434;
	{8'd50,8'd69} : s = 497;
	{8'd50,8'd70} : s = 325;
	{8'd50,8'd71} : s = 433;
	{8'd50,8'd72} : s = 428;
	{8'd50,8'd73} : s = 492;
	{8'd50,8'd74} : s = 426;
	{8'd50,8'd75} : s = 490;
	{8'd50,8'd76} : s = 489;
	{8'd50,8'd77} : s = 508;
	{8'd50,8'd78} : s = 2;
	{8'd50,8'd79} : s = 48;
	{8'd50,8'd80} : s = 40;
	{8'd50,8'd81} : s = 168;
	{8'd50,8'd82} : s = 36;
	{8'd50,8'd83} : s = 164;
	{8'd50,8'd84} : s = 162;
	{8'd50,8'd85} : s = 323;
	{8'd50,8'd86} : s = 34;
	{8'd50,8'd87} : s = 161;
	{8'd50,8'd88} : s = 152;
	{8'd50,8'd89} : s = 312;
	{8'd50,8'd90} : s = 148;
	{8'd50,8'd91} : s = 308;
	{8'd50,8'd92} : s = 306;
	{8'd50,8'd93} : s = 425;
	{8'd50,8'd94} : s = 33;
	{8'd50,8'd95} : s = 146;
	{8'd50,8'd96} : s = 145;
	{8'd50,8'd97} : s = 305;
	{8'd50,8'd98} : s = 140;
	{8'd50,8'd99} : s = 300;
	{8'd50,8'd100} : s = 298;
	{8'd50,8'd101} : s = 422;
	{8'd50,8'd102} : s = 138;
	{8'd50,8'd103} : s = 297;
	{8'd50,8'd104} : s = 294;
	{8'd50,8'd105} : s = 421;
	{8'd50,8'd106} : s = 293;
	{8'd50,8'd107} : s = 419;
	{8'd50,8'd108} : s = 412;
	{8'd50,8'd109} : s = 486;
	{8'd50,8'd110} : s = 24;
	{8'd50,8'd111} : s = 137;
	{8'd50,8'd112} : s = 134;
	{8'd50,8'd113} : s = 291;
	{8'd50,8'd114} : s = 133;
	{8'd50,8'd115} : s = 284;
	{8'd50,8'd116} : s = 282;
	{8'd50,8'd117} : s = 410;
	{8'd50,8'd118} : s = 131;
	{8'd50,8'd119} : s = 281;
	{8'd50,8'd120} : s = 278;
	{8'd50,8'd121} : s = 409;
	{8'd50,8'd122} : s = 277;
	{8'd50,8'd123} : s = 406;
	{8'd50,8'd124} : s = 405;
	{8'd50,8'd125} : s = 485;
	{8'd50,8'd126} : s = 112;
	{8'd50,8'd127} : s = 275;
	{8'd50,8'd128} : s = 270;
	{8'd50,8'd129} : s = 403;
	{8'd50,8'd130} : s = 269;
	{8'd50,8'd131} : s = 398;
	{8'd50,8'd132} : s = 397;
	{8'd50,8'd133} : s = 483;
	{8'd50,8'd134} : s = 267;
	{8'd50,8'd135} : s = 395;
	{8'd50,8'd136} : s = 391;
	{8'd50,8'd137} : s = 476;
	{8'd50,8'd138} : s = 376;
	{8'd50,8'd139} : s = 474;
	{8'd50,8'd140} : s = 473;
	{8'd50,8'd141} : s = 506;
	{8'd50,8'd142} : s = 20;
	{8'd50,8'd143} : s = 104;
	{8'd50,8'd144} : s = 100;
	{8'd50,8'd145} : s = 263;
	{8'd50,8'd146} : s = 98;
	{8'd50,8'd147} : s = 240;
	{8'd50,8'd148} : s = 232;
	{8'd50,8'd149} : s = 372;
	{8'd50,8'd150} : s = 97;
	{8'd50,8'd151} : s = 228;
	{8'd50,8'd152} : s = 226;
	{8'd50,8'd153} : s = 370;
	{8'd50,8'd154} : s = 225;
	{8'd50,8'd155} : s = 369;
	{8'd50,8'd156} : s = 364;
	{8'd50,8'd157} : s = 470;
	{8'd50,8'd158} : s = 88;
	{8'd50,8'd159} : s = 216;
	{8'd50,8'd160} : s = 212;
	{8'd50,8'd161} : s = 362;
	{8'd50,8'd162} : s = 210;
	{8'd50,8'd163} : s = 361;
	{8'd50,8'd164} : s = 358;
	{8'd50,8'd165} : s = 469;
	{8'd50,8'd166} : s = 209;
	{8'd50,8'd167} : s = 357;
	{8'd50,8'd168} : s = 355;
	{8'd50,8'd169} : s = 467;
	{8'd50,8'd170} : s = 348;
	{8'd50,8'd171} : s = 462;
	{8'd50,8'd172} : s = 461;
	{8'd50,8'd173} : s = 505;
	{8'd50,8'd174} : s = 84;
	{8'd50,8'd175} : s = 204;
	{8'd50,8'd176} : s = 202;
	{8'd50,8'd177} : s = 346;
	{8'd50,8'd178} : s = 201;
	{8'd50,8'd179} : s = 345;
	{8'd50,8'd180} : s = 342;
	{8'd50,8'd181} : s = 459;
	{8'd50,8'd182} : s = 198;
	{8'd50,8'd183} : s = 341;
	{8'd50,8'd184} : s = 339;
	{8'd50,8'd185} : s = 455;
	{8'd50,8'd186} : s = 334;
	{8'd50,8'd187} : s = 444;
	{8'd50,8'd188} : s = 442;
	{8'd50,8'd189} : s = 502;
	{8'd50,8'd190} : s = 197;
	{8'd50,8'd191} : s = 333;
	{8'd50,8'd192} : s = 331;
	{8'd50,8'd193} : s = 441;
	{8'd50,8'd194} : s = 327;
	{8'd50,8'd195} : s = 438;
	{8'd50,8'd196} : s = 437;
	{8'd50,8'd197} : s = 501;
	{8'd50,8'd198} : s = 316;
	{8'd50,8'd199} : s = 435;
	{8'd50,8'd200} : s = 430;
	{8'd50,8'd201} : s = 499;
	{8'd50,8'd202} : s = 429;
	{8'd50,8'd203} : s = 494;
	{8'd50,8'd204} : s = 493;
	{8'd50,8'd205} : s = 510;
	{8'd50,8'd206} : s = 1;
	{8'd50,8'd207} : s = 18;
	{8'd50,8'd208} : s = 17;
	{8'd50,8'd209} : s = 82;
	{8'd50,8'd210} : s = 12;
	{8'd50,8'd211} : s = 81;
	{8'd50,8'd212} : s = 76;
	{8'd50,8'd213} : s = 195;
	{8'd50,8'd214} : s = 10;
	{8'd50,8'd215} : s = 74;
	{8'd50,8'd216} : s = 73;
	{8'd50,8'd217} : s = 184;
	{8'd50,8'd218} : s = 70;
	{8'd50,8'd219} : s = 180;
	{8'd50,8'd220} : s = 178;
	{8'd50,8'd221} : s = 314;
	{8'd50,8'd222} : s = 9;
	{8'd50,8'd223} : s = 69;
	{8'd50,8'd224} : s = 67;
	{8'd50,8'd225} : s = 177;
	{8'd50,8'd226} : s = 56;
	{8'd50,8'd227} : s = 172;
	{8'd50,8'd228} : s = 170;
	{8'd50,8'd229} : s = 313;
	{8'd50,8'd230} : s = 52;
	{8'd50,8'd231} : s = 169;
	{8'd50,8'd232} : s = 166;
	{8'd50,8'd233} : s = 310;
	{8'd50,8'd234} : s = 165;
	{8'd50,8'd235} : s = 309;
	{8'd50,8'd236} : s = 307;
	{8'd50,8'd237} : s = 427;
	{8'd50,8'd238} : s = 6;
	{8'd50,8'd239} : s = 50;
	{8'd50,8'd240} : s = 49;
	{8'd50,8'd241} : s = 163;
	{8'd50,8'd242} : s = 44;
	{8'd50,8'd243} : s = 156;
	{8'd50,8'd244} : s = 154;
	{8'd50,8'd245} : s = 302;
	{8'd50,8'd246} : s = 42;
	{8'd50,8'd247} : s = 153;
	{8'd50,8'd248} : s = 150;
	{8'd50,8'd249} : s = 301;
	{8'd50,8'd250} : s = 149;
	{8'd50,8'd251} : s = 299;
	{8'd50,8'd252} : s = 295;
	{8'd50,8'd253} : s = 423;
	{8'd50,8'd254} : s = 41;
	{8'd50,8'd255} : s = 147;
	{8'd51,8'd0} : s = 418;
	{8'd51,8'd1} : s = 280;
	{8'd51,8'd2} : s = 417;
	{8'd51,8'd3} : s = 408;
	{8'd51,8'd4} : s = 484;
	{8'd51,8'd5} : s = 276;
	{8'd51,8'd6} : s = 404;
	{8'd51,8'd7} : s = 402;
	{8'd51,8'd8} : s = 482;
	{8'd51,8'd9} : s = 401;
	{8'd51,8'd10} : s = 481;
	{8'd51,8'd11} : s = 472;
	{8'd51,8'd12} : s = 504;
	{8'd51,8'd13} : s = 4;
	{8'd51,8'd14} : s = 96;
	{8'd51,8'd15} : s = 80;
	{8'd51,8'd16} : s = 274;
	{8'd51,8'd17} : s = 72;
	{8'd51,8'd18} : s = 273;
	{8'd51,8'd19} : s = 268;
	{8'd51,8'd20} : s = 396;
	{8'd51,8'd21} : s = 68;
	{8'd51,8'd22} : s = 266;
	{8'd51,8'd23} : s = 265;
	{8'd51,8'd24} : s = 394;
	{8'd51,8'd25} : s = 262;
	{8'd51,8'd26} : s = 393;
	{8'd51,8'd27} : s = 390;
	{8'd51,8'd28} : s = 468;
	{8'd51,8'd29} : s = 66;
	{8'd51,8'd30} : s = 261;
	{8'd51,8'd31} : s = 259;
	{8'd51,8'd32} : s = 389;
	{8'd51,8'd33} : s = 224;
	{8'd51,8'd34} : s = 387;
	{8'd51,8'd35} : s = 368;
	{8'd51,8'd36} : s = 466;
	{8'd51,8'd37} : s = 208;
	{8'd51,8'd38} : s = 360;
	{8'd51,8'd39} : s = 356;
	{8'd51,8'd40} : s = 465;
	{8'd51,8'd41} : s = 354;
	{8'd51,8'd42} : s = 460;
	{8'd51,8'd43} : s = 458;
	{8'd51,8'd44} : s = 500;
	{8'd51,8'd45} : s = 65;
	{8'd51,8'd46} : s = 200;
	{8'd51,8'd47} : s = 196;
	{8'd51,8'd48} : s = 353;
	{8'd51,8'd49} : s = 194;
	{8'd51,8'd50} : s = 344;
	{8'd51,8'd51} : s = 340;
	{8'd51,8'd52} : s = 457;
	{8'd51,8'd53} : s = 193;
	{8'd51,8'd54} : s = 338;
	{8'd51,8'd55} : s = 337;
	{8'd51,8'd56} : s = 454;
	{8'd51,8'd57} : s = 332;
	{8'd51,8'd58} : s = 453;
	{8'd51,8'd59} : s = 451;
	{8'd51,8'd60} : s = 498;
	{8'd51,8'd61} : s = 176;
	{8'd51,8'd62} : s = 330;
	{8'd51,8'd63} : s = 329;
	{8'd51,8'd64} : s = 440;
	{8'd51,8'd65} : s = 326;
	{8'd51,8'd66} : s = 436;
	{8'd51,8'd67} : s = 434;
	{8'd51,8'd68} : s = 497;
	{8'd51,8'd69} : s = 325;
	{8'd51,8'd70} : s = 433;
	{8'd51,8'd71} : s = 428;
	{8'd51,8'd72} : s = 492;
	{8'd51,8'd73} : s = 426;
	{8'd51,8'd74} : s = 490;
	{8'd51,8'd75} : s = 489;
	{8'd51,8'd76} : s = 508;
	{8'd51,8'd77} : s = 2;
	{8'd51,8'd78} : s = 48;
	{8'd51,8'd79} : s = 40;
	{8'd51,8'd80} : s = 168;
	{8'd51,8'd81} : s = 36;
	{8'd51,8'd82} : s = 164;
	{8'd51,8'd83} : s = 162;
	{8'd51,8'd84} : s = 323;
	{8'd51,8'd85} : s = 34;
	{8'd51,8'd86} : s = 161;
	{8'd51,8'd87} : s = 152;
	{8'd51,8'd88} : s = 312;
	{8'd51,8'd89} : s = 148;
	{8'd51,8'd90} : s = 308;
	{8'd51,8'd91} : s = 306;
	{8'd51,8'd92} : s = 425;
	{8'd51,8'd93} : s = 33;
	{8'd51,8'd94} : s = 146;
	{8'd51,8'd95} : s = 145;
	{8'd51,8'd96} : s = 305;
	{8'd51,8'd97} : s = 140;
	{8'd51,8'd98} : s = 300;
	{8'd51,8'd99} : s = 298;
	{8'd51,8'd100} : s = 422;
	{8'd51,8'd101} : s = 138;
	{8'd51,8'd102} : s = 297;
	{8'd51,8'd103} : s = 294;
	{8'd51,8'd104} : s = 421;
	{8'd51,8'd105} : s = 293;
	{8'd51,8'd106} : s = 419;
	{8'd51,8'd107} : s = 412;
	{8'd51,8'd108} : s = 486;
	{8'd51,8'd109} : s = 24;
	{8'd51,8'd110} : s = 137;
	{8'd51,8'd111} : s = 134;
	{8'd51,8'd112} : s = 291;
	{8'd51,8'd113} : s = 133;
	{8'd51,8'd114} : s = 284;
	{8'd51,8'd115} : s = 282;
	{8'd51,8'd116} : s = 410;
	{8'd51,8'd117} : s = 131;
	{8'd51,8'd118} : s = 281;
	{8'd51,8'd119} : s = 278;
	{8'd51,8'd120} : s = 409;
	{8'd51,8'd121} : s = 277;
	{8'd51,8'd122} : s = 406;
	{8'd51,8'd123} : s = 405;
	{8'd51,8'd124} : s = 485;
	{8'd51,8'd125} : s = 112;
	{8'd51,8'd126} : s = 275;
	{8'd51,8'd127} : s = 270;
	{8'd51,8'd128} : s = 403;
	{8'd51,8'd129} : s = 269;
	{8'd51,8'd130} : s = 398;
	{8'd51,8'd131} : s = 397;
	{8'd51,8'd132} : s = 483;
	{8'd51,8'd133} : s = 267;
	{8'd51,8'd134} : s = 395;
	{8'd51,8'd135} : s = 391;
	{8'd51,8'd136} : s = 476;
	{8'd51,8'd137} : s = 376;
	{8'd51,8'd138} : s = 474;
	{8'd51,8'd139} : s = 473;
	{8'd51,8'd140} : s = 506;
	{8'd51,8'd141} : s = 20;
	{8'd51,8'd142} : s = 104;
	{8'd51,8'd143} : s = 100;
	{8'd51,8'd144} : s = 263;
	{8'd51,8'd145} : s = 98;
	{8'd51,8'd146} : s = 240;
	{8'd51,8'd147} : s = 232;
	{8'd51,8'd148} : s = 372;
	{8'd51,8'd149} : s = 97;
	{8'd51,8'd150} : s = 228;
	{8'd51,8'd151} : s = 226;
	{8'd51,8'd152} : s = 370;
	{8'd51,8'd153} : s = 225;
	{8'd51,8'd154} : s = 369;
	{8'd51,8'd155} : s = 364;
	{8'd51,8'd156} : s = 470;
	{8'd51,8'd157} : s = 88;
	{8'd51,8'd158} : s = 216;
	{8'd51,8'd159} : s = 212;
	{8'd51,8'd160} : s = 362;
	{8'd51,8'd161} : s = 210;
	{8'd51,8'd162} : s = 361;
	{8'd51,8'd163} : s = 358;
	{8'd51,8'd164} : s = 469;
	{8'd51,8'd165} : s = 209;
	{8'd51,8'd166} : s = 357;
	{8'd51,8'd167} : s = 355;
	{8'd51,8'd168} : s = 467;
	{8'd51,8'd169} : s = 348;
	{8'd51,8'd170} : s = 462;
	{8'd51,8'd171} : s = 461;
	{8'd51,8'd172} : s = 505;
	{8'd51,8'd173} : s = 84;
	{8'd51,8'd174} : s = 204;
	{8'd51,8'd175} : s = 202;
	{8'd51,8'd176} : s = 346;
	{8'd51,8'd177} : s = 201;
	{8'd51,8'd178} : s = 345;
	{8'd51,8'd179} : s = 342;
	{8'd51,8'd180} : s = 459;
	{8'd51,8'd181} : s = 198;
	{8'd51,8'd182} : s = 341;
	{8'd51,8'd183} : s = 339;
	{8'd51,8'd184} : s = 455;
	{8'd51,8'd185} : s = 334;
	{8'd51,8'd186} : s = 444;
	{8'd51,8'd187} : s = 442;
	{8'd51,8'd188} : s = 502;
	{8'd51,8'd189} : s = 197;
	{8'd51,8'd190} : s = 333;
	{8'd51,8'd191} : s = 331;
	{8'd51,8'd192} : s = 441;
	{8'd51,8'd193} : s = 327;
	{8'd51,8'd194} : s = 438;
	{8'd51,8'd195} : s = 437;
	{8'd51,8'd196} : s = 501;
	{8'd51,8'd197} : s = 316;
	{8'd51,8'd198} : s = 435;
	{8'd51,8'd199} : s = 430;
	{8'd51,8'd200} : s = 499;
	{8'd51,8'd201} : s = 429;
	{8'd51,8'd202} : s = 494;
	{8'd51,8'd203} : s = 493;
	{8'd51,8'd204} : s = 510;
	{8'd51,8'd205} : s = 1;
	{8'd51,8'd206} : s = 18;
	{8'd51,8'd207} : s = 17;
	{8'd51,8'd208} : s = 82;
	{8'd51,8'd209} : s = 12;
	{8'd51,8'd210} : s = 81;
	{8'd51,8'd211} : s = 76;
	{8'd51,8'd212} : s = 195;
	{8'd51,8'd213} : s = 10;
	{8'd51,8'd214} : s = 74;
	{8'd51,8'd215} : s = 73;
	{8'd51,8'd216} : s = 184;
	{8'd51,8'd217} : s = 70;
	{8'd51,8'd218} : s = 180;
	{8'd51,8'd219} : s = 178;
	{8'd51,8'd220} : s = 314;
	{8'd51,8'd221} : s = 9;
	{8'd51,8'd222} : s = 69;
	{8'd51,8'd223} : s = 67;
	{8'd51,8'd224} : s = 177;
	{8'd51,8'd225} : s = 56;
	{8'd51,8'd226} : s = 172;
	{8'd51,8'd227} : s = 170;
	{8'd51,8'd228} : s = 313;
	{8'd51,8'd229} : s = 52;
	{8'd51,8'd230} : s = 169;
	{8'd51,8'd231} : s = 166;
	{8'd51,8'd232} : s = 310;
	{8'd51,8'd233} : s = 165;
	{8'd51,8'd234} : s = 309;
	{8'd51,8'd235} : s = 307;
	{8'd51,8'd236} : s = 427;
	{8'd51,8'd237} : s = 6;
	{8'd51,8'd238} : s = 50;
	{8'd51,8'd239} : s = 49;
	{8'd51,8'd240} : s = 163;
	{8'd51,8'd241} : s = 44;
	{8'd51,8'd242} : s = 156;
	{8'd51,8'd243} : s = 154;
	{8'd51,8'd244} : s = 302;
	{8'd51,8'd245} : s = 42;
	{8'd51,8'd246} : s = 153;
	{8'd51,8'd247} : s = 150;
	{8'd51,8'd248} : s = 301;
	{8'd51,8'd249} : s = 149;
	{8'd51,8'd250} : s = 299;
	{8'd51,8'd251} : s = 295;
	{8'd51,8'd252} : s = 423;
	{8'd51,8'd253} : s = 41;
	{8'd51,8'd254} : s = 147;
	{8'd51,8'd255} : s = 142;
	{8'd52,8'd0} : s = 280;
	{8'd52,8'd1} : s = 417;
	{8'd52,8'd2} : s = 408;
	{8'd52,8'd3} : s = 484;
	{8'd52,8'd4} : s = 276;
	{8'd52,8'd5} : s = 404;
	{8'd52,8'd6} : s = 402;
	{8'd52,8'd7} : s = 482;
	{8'd52,8'd8} : s = 401;
	{8'd52,8'd9} : s = 481;
	{8'd52,8'd10} : s = 472;
	{8'd52,8'd11} : s = 504;
	{8'd52,8'd12} : s = 4;
	{8'd52,8'd13} : s = 96;
	{8'd52,8'd14} : s = 80;
	{8'd52,8'd15} : s = 274;
	{8'd52,8'd16} : s = 72;
	{8'd52,8'd17} : s = 273;
	{8'd52,8'd18} : s = 268;
	{8'd52,8'd19} : s = 396;
	{8'd52,8'd20} : s = 68;
	{8'd52,8'd21} : s = 266;
	{8'd52,8'd22} : s = 265;
	{8'd52,8'd23} : s = 394;
	{8'd52,8'd24} : s = 262;
	{8'd52,8'd25} : s = 393;
	{8'd52,8'd26} : s = 390;
	{8'd52,8'd27} : s = 468;
	{8'd52,8'd28} : s = 66;
	{8'd52,8'd29} : s = 261;
	{8'd52,8'd30} : s = 259;
	{8'd52,8'd31} : s = 389;
	{8'd52,8'd32} : s = 224;
	{8'd52,8'd33} : s = 387;
	{8'd52,8'd34} : s = 368;
	{8'd52,8'd35} : s = 466;
	{8'd52,8'd36} : s = 208;
	{8'd52,8'd37} : s = 360;
	{8'd52,8'd38} : s = 356;
	{8'd52,8'd39} : s = 465;
	{8'd52,8'd40} : s = 354;
	{8'd52,8'd41} : s = 460;
	{8'd52,8'd42} : s = 458;
	{8'd52,8'd43} : s = 500;
	{8'd52,8'd44} : s = 65;
	{8'd52,8'd45} : s = 200;
	{8'd52,8'd46} : s = 196;
	{8'd52,8'd47} : s = 353;
	{8'd52,8'd48} : s = 194;
	{8'd52,8'd49} : s = 344;
	{8'd52,8'd50} : s = 340;
	{8'd52,8'd51} : s = 457;
	{8'd52,8'd52} : s = 193;
	{8'd52,8'd53} : s = 338;
	{8'd52,8'd54} : s = 337;
	{8'd52,8'd55} : s = 454;
	{8'd52,8'd56} : s = 332;
	{8'd52,8'd57} : s = 453;
	{8'd52,8'd58} : s = 451;
	{8'd52,8'd59} : s = 498;
	{8'd52,8'd60} : s = 176;
	{8'd52,8'd61} : s = 330;
	{8'd52,8'd62} : s = 329;
	{8'd52,8'd63} : s = 440;
	{8'd52,8'd64} : s = 326;
	{8'd52,8'd65} : s = 436;
	{8'd52,8'd66} : s = 434;
	{8'd52,8'd67} : s = 497;
	{8'd52,8'd68} : s = 325;
	{8'd52,8'd69} : s = 433;
	{8'd52,8'd70} : s = 428;
	{8'd52,8'd71} : s = 492;
	{8'd52,8'd72} : s = 426;
	{8'd52,8'd73} : s = 490;
	{8'd52,8'd74} : s = 489;
	{8'd52,8'd75} : s = 508;
	{8'd52,8'd76} : s = 2;
	{8'd52,8'd77} : s = 48;
	{8'd52,8'd78} : s = 40;
	{8'd52,8'd79} : s = 168;
	{8'd52,8'd80} : s = 36;
	{8'd52,8'd81} : s = 164;
	{8'd52,8'd82} : s = 162;
	{8'd52,8'd83} : s = 323;
	{8'd52,8'd84} : s = 34;
	{8'd52,8'd85} : s = 161;
	{8'd52,8'd86} : s = 152;
	{8'd52,8'd87} : s = 312;
	{8'd52,8'd88} : s = 148;
	{8'd52,8'd89} : s = 308;
	{8'd52,8'd90} : s = 306;
	{8'd52,8'd91} : s = 425;
	{8'd52,8'd92} : s = 33;
	{8'd52,8'd93} : s = 146;
	{8'd52,8'd94} : s = 145;
	{8'd52,8'd95} : s = 305;
	{8'd52,8'd96} : s = 140;
	{8'd52,8'd97} : s = 300;
	{8'd52,8'd98} : s = 298;
	{8'd52,8'd99} : s = 422;
	{8'd52,8'd100} : s = 138;
	{8'd52,8'd101} : s = 297;
	{8'd52,8'd102} : s = 294;
	{8'd52,8'd103} : s = 421;
	{8'd52,8'd104} : s = 293;
	{8'd52,8'd105} : s = 419;
	{8'd52,8'd106} : s = 412;
	{8'd52,8'd107} : s = 486;
	{8'd52,8'd108} : s = 24;
	{8'd52,8'd109} : s = 137;
	{8'd52,8'd110} : s = 134;
	{8'd52,8'd111} : s = 291;
	{8'd52,8'd112} : s = 133;
	{8'd52,8'd113} : s = 284;
	{8'd52,8'd114} : s = 282;
	{8'd52,8'd115} : s = 410;
	{8'd52,8'd116} : s = 131;
	{8'd52,8'd117} : s = 281;
	{8'd52,8'd118} : s = 278;
	{8'd52,8'd119} : s = 409;
	{8'd52,8'd120} : s = 277;
	{8'd52,8'd121} : s = 406;
	{8'd52,8'd122} : s = 405;
	{8'd52,8'd123} : s = 485;
	{8'd52,8'd124} : s = 112;
	{8'd52,8'd125} : s = 275;
	{8'd52,8'd126} : s = 270;
	{8'd52,8'd127} : s = 403;
	{8'd52,8'd128} : s = 269;
	{8'd52,8'd129} : s = 398;
	{8'd52,8'd130} : s = 397;
	{8'd52,8'd131} : s = 483;
	{8'd52,8'd132} : s = 267;
	{8'd52,8'd133} : s = 395;
	{8'd52,8'd134} : s = 391;
	{8'd52,8'd135} : s = 476;
	{8'd52,8'd136} : s = 376;
	{8'd52,8'd137} : s = 474;
	{8'd52,8'd138} : s = 473;
	{8'd52,8'd139} : s = 506;
	{8'd52,8'd140} : s = 20;
	{8'd52,8'd141} : s = 104;
	{8'd52,8'd142} : s = 100;
	{8'd52,8'd143} : s = 263;
	{8'd52,8'd144} : s = 98;
	{8'd52,8'd145} : s = 240;
	{8'd52,8'd146} : s = 232;
	{8'd52,8'd147} : s = 372;
	{8'd52,8'd148} : s = 97;
	{8'd52,8'd149} : s = 228;
	{8'd52,8'd150} : s = 226;
	{8'd52,8'd151} : s = 370;
	{8'd52,8'd152} : s = 225;
	{8'd52,8'd153} : s = 369;
	{8'd52,8'd154} : s = 364;
	{8'd52,8'd155} : s = 470;
	{8'd52,8'd156} : s = 88;
	{8'd52,8'd157} : s = 216;
	{8'd52,8'd158} : s = 212;
	{8'd52,8'd159} : s = 362;
	{8'd52,8'd160} : s = 210;
	{8'd52,8'd161} : s = 361;
	{8'd52,8'd162} : s = 358;
	{8'd52,8'd163} : s = 469;
	{8'd52,8'd164} : s = 209;
	{8'd52,8'd165} : s = 357;
	{8'd52,8'd166} : s = 355;
	{8'd52,8'd167} : s = 467;
	{8'd52,8'd168} : s = 348;
	{8'd52,8'd169} : s = 462;
	{8'd52,8'd170} : s = 461;
	{8'd52,8'd171} : s = 505;
	{8'd52,8'd172} : s = 84;
	{8'd52,8'd173} : s = 204;
	{8'd52,8'd174} : s = 202;
	{8'd52,8'd175} : s = 346;
	{8'd52,8'd176} : s = 201;
	{8'd52,8'd177} : s = 345;
	{8'd52,8'd178} : s = 342;
	{8'd52,8'd179} : s = 459;
	{8'd52,8'd180} : s = 198;
	{8'd52,8'd181} : s = 341;
	{8'd52,8'd182} : s = 339;
	{8'd52,8'd183} : s = 455;
	{8'd52,8'd184} : s = 334;
	{8'd52,8'd185} : s = 444;
	{8'd52,8'd186} : s = 442;
	{8'd52,8'd187} : s = 502;
	{8'd52,8'd188} : s = 197;
	{8'd52,8'd189} : s = 333;
	{8'd52,8'd190} : s = 331;
	{8'd52,8'd191} : s = 441;
	{8'd52,8'd192} : s = 327;
	{8'd52,8'd193} : s = 438;
	{8'd52,8'd194} : s = 437;
	{8'd52,8'd195} : s = 501;
	{8'd52,8'd196} : s = 316;
	{8'd52,8'd197} : s = 435;
	{8'd52,8'd198} : s = 430;
	{8'd52,8'd199} : s = 499;
	{8'd52,8'd200} : s = 429;
	{8'd52,8'd201} : s = 494;
	{8'd52,8'd202} : s = 493;
	{8'd52,8'd203} : s = 510;
	{8'd52,8'd204} : s = 1;
	{8'd52,8'd205} : s = 18;
	{8'd52,8'd206} : s = 17;
	{8'd52,8'd207} : s = 82;
	{8'd52,8'd208} : s = 12;
	{8'd52,8'd209} : s = 81;
	{8'd52,8'd210} : s = 76;
	{8'd52,8'd211} : s = 195;
	{8'd52,8'd212} : s = 10;
	{8'd52,8'd213} : s = 74;
	{8'd52,8'd214} : s = 73;
	{8'd52,8'd215} : s = 184;
	{8'd52,8'd216} : s = 70;
	{8'd52,8'd217} : s = 180;
	{8'd52,8'd218} : s = 178;
	{8'd52,8'd219} : s = 314;
	{8'd52,8'd220} : s = 9;
	{8'd52,8'd221} : s = 69;
	{8'd52,8'd222} : s = 67;
	{8'd52,8'd223} : s = 177;
	{8'd52,8'd224} : s = 56;
	{8'd52,8'd225} : s = 172;
	{8'd52,8'd226} : s = 170;
	{8'd52,8'd227} : s = 313;
	{8'd52,8'd228} : s = 52;
	{8'd52,8'd229} : s = 169;
	{8'd52,8'd230} : s = 166;
	{8'd52,8'd231} : s = 310;
	{8'd52,8'd232} : s = 165;
	{8'd52,8'd233} : s = 309;
	{8'd52,8'd234} : s = 307;
	{8'd52,8'd235} : s = 427;
	{8'd52,8'd236} : s = 6;
	{8'd52,8'd237} : s = 50;
	{8'd52,8'd238} : s = 49;
	{8'd52,8'd239} : s = 163;
	{8'd52,8'd240} : s = 44;
	{8'd52,8'd241} : s = 156;
	{8'd52,8'd242} : s = 154;
	{8'd52,8'd243} : s = 302;
	{8'd52,8'd244} : s = 42;
	{8'd52,8'd245} : s = 153;
	{8'd52,8'd246} : s = 150;
	{8'd52,8'd247} : s = 301;
	{8'd52,8'd248} : s = 149;
	{8'd52,8'd249} : s = 299;
	{8'd52,8'd250} : s = 295;
	{8'd52,8'd251} : s = 423;
	{8'd52,8'd252} : s = 41;
	{8'd52,8'd253} : s = 147;
	{8'd52,8'd254} : s = 142;
	{8'd52,8'd255} : s = 286;
	{8'd53,8'd0} : s = 417;
	{8'd53,8'd1} : s = 408;
	{8'd53,8'd2} : s = 484;
	{8'd53,8'd3} : s = 276;
	{8'd53,8'd4} : s = 404;
	{8'd53,8'd5} : s = 402;
	{8'd53,8'd6} : s = 482;
	{8'd53,8'd7} : s = 401;
	{8'd53,8'd8} : s = 481;
	{8'd53,8'd9} : s = 472;
	{8'd53,8'd10} : s = 504;
	{8'd53,8'd11} : s = 4;
	{8'd53,8'd12} : s = 96;
	{8'd53,8'd13} : s = 80;
	{8'd53,8'd14} : s = 274;
	{8'd53,8'd15} : s = 72;
	{8'd53,8'd16} : s = 273;
	{8'd53,8'd17} : s = 268;
	{8'd53,8'd18} : s = 396;
	{8'd53,8'd19} : s = 68;
	{8'd53,8'd20} : s = 266;
	{8'd53,8'd21} : s = 265;
	{8'd53,8'd22} : s = 394;
	{8'd53,8'd23} : s = 262;
	{8'd53,8'd24} : s = 393;
	{8'd53,8'd25} : s = 390;
	{8'd53,8'd26} : s = 468;
	{8'd53,8'd27} : s = 66;
	{8'd53,8'd28} : s = 261;
	{8'd53,8'd29} : s = 259;
	{8'd53,8'd30} : s = 389;
	{8'd53,8'd31} : s = 224;
	{8'd53,8'd32} : s = 387;
	{8'd53,8'd33} : s = 368;
	{8'd53,8'd34} : s = 466;
	{8'd53,8'd35} : s = 208;
	{8'd53,8'd36} : s = 360;
	{8'd53,8'd37} : s = 356;
	{8'd53,8'd38} : s = 465;
	{8'd53,8'd39} : s = 354;
	{8'd53,8'd40} : s = 460;
	{8'd53,8'd41} : s = 458;
	{8'd53,8'd42} : s = 500;
	{8'd53,8'd43} : s = 65;
	{8'd53,8'd44} : s = 200;
	{8'd53,8'd45} : s = 196;
	{8'd53,8'd46} : s = 353;
	{8'd53,8'd47} : s = 194;
	{8'd53,8'd48} : s = 344;
	{8'd53,8'd49} : s = 340;
	{8'd53,8'd50} : s = 457;
	{8'd53,8'd51} : s = 193;
	{8'd53,8'd52} : s = 338;
	{8'd53,8'd53} : s = 337;
	{8'd53,8'd54} : s = 454;
	{8'd53,8'd55} : s = 332;
	{8'd53,8'd56} : s = 453;
	{8'd53,8'd57} : s = 451;
	{8'd53,8'd58} : s = 498;
	{8'd53,8'd59} : s = 176;
	{8'd53,8'd60} : s = 330;
	{8'd53,8'd61} : s = 329;
	{8'd53,8'd62} : s = 440;
	{8'd53,8'd63} : s = 326;
	{8'd53,8'd64} : s = 436;
	{8'd53,8'd65} : s = 434;
	{8'd53,8'd66} : s = 497;
	{8'd53,8'd67} : s = 325;
	{8'd53,8'd68} : s = 433;
	{8'd53,8'd69} : s = 428;
	{8'd53,8'd70} : s = 492;
	{8'd53,8'd71} : s = 426;
	{8'd53,8'd72} : s = 490;
	{8'd53,8'd73} : s = 489;
	{8'd53,8'd74} : s = 508;
	{8'd53,8'd75} : s = 2;
	{8'd53,8'd76} : s = 48;
	{8'd53,8'd77} : s = 40;
	{8'd53,8'd78} : s = 168;
	{8'd53,8'd79} : s = 36;
	{8'd53,8'd80} : s = 164;
	{8'd53,8'd81} : s = 162;
	{8'd53,8'd82} : s = 323;
	{8'd53,8'd83} : s = 34;
	{8'd53,8'd84} : s = 161;
	{8'd53,8'd85} : s = 152;
	{8'd53,8'd86} : s = 312;
	{8'd53,8'd87} : s = 148;
	{8'd53,8'd88} : s = 308;
	{8'd53,8'd89} : s = 306;
	{8'd53,8'd90} : s = 425;
	{8'd53,8'd91} : s = 33;
	{8'd53,8'd92} : s = 146;
	{8'd53,8'd93} : s = 145;
	{8'd53,8'd94} : s = 305;
	{8'd53,8'd95} : s = 140;
	{8'd53,8'd96} : s = 300;
	{8'd53,8'd97} : s = 298;
	{8'd53,8'd98} : s = 422;
	{8'd53,8'd99} : s = 138;
	{8'd53,8'd100} : s = 297;
	{8'd53,8'd101} : s = 294;
	{8'd53,8'd102} : s = 421;
	{8'd53,8'd103} : s = 293;
	{8'd53,8'd104} : s = 419;
	{8'd53,8'd105} : s = 412;
	{8'd53,8'd106} : s = 486;
	{8'd53,8'd107} : s = 24;
	{8'd53,8'd108} : s = 137;
	{8'd53,8'd109} : s = 134;
	{8'd53,8'd110} : s = 291;
	{8'd53,8'd111} : s = 133;
	{8'd53,8'd112} : s = 284;
	{8'd53,8'd113} : s = 282;
	{8'd53,8'd114} : s = 410;
	{8'd53,8'd115} : s = 131;
	{8'd53,8'd116} : s = 281;
	{8'd53,8'd117} : s = 278;
	{8'd53,8'd118} : s = 409;
	{8'd53,8'd119} : s = 277;
	{8'd53,8'd120} : s = 406;
	{8'd53,8'd121} : s = 405;
	{8'd53,8'd122} : s = 485;
	{8'd53,8'd123} : s = 112;
	{8'd53,8'd124} : s = 275;
	{8'd53,8'd125} : s = 270;
	{8'd53,8'd126} : s = 403;
	{8'd53,8'd127} : s = 269;
	{8'd53,8'd128} : s = 398;
	{8'd53,8'd129} : s = 397;
	{8'd53,8'd130} : s = 483;
	{8'd53,8'd131} : s = 267;
	{8'd53,8'd132} : s = 395;
	{8'd53,8'd133} : s = 391;
	{8'd53,8'd134} : s = 476;
	{8'd53,8'd135} : s = 376;
	{8'd53,8'd136} : s = 474;
	{8'd53,8'd137} : s = 473;
	{8'd53,8'd138} : s = 506;
	{8'd53,8'd139} : s = 20;
	{8'd53,8'd140} : s = 104;
	{8'd53,8'd141} : s = 100;
	{8'd53,8'd142} : s = 263;
	{8'd53,8'd143} : s = 98;
	{8'd53,8'd144} : s = 240;
	{8'd53,8'd145} : s = 232;
	{8'd53,8'd146} : s = 372;
	{8'd53,8'd147} : s = 97;
	{8'd53,8'd148} : s = 228;
	{8'd53,8'd149} : s = 226;
	{8'd53,8'd150} : s = 370;
	{8'd53,8'd151} : s = 225;
	{8'd53,8'd152} : s = 369;
	{8'd53,8'd153} : s = 364;
	{8'd53,8'd154} : s = 470;
	{8'd53,8'd155} : s = 88;
	{8'd53,8'd156} : s = 216;
	{8'd53,8'd157} : s = 212;
	{8'd53,8'd158} : s = 362;
	{8'd53,8'd159} : s = 210;
	{8'd53,8'd160} : s = 361;
	{8'd53,8'd161} : s = 358;
	{8'd53,8'd162} : s = 469;
	{8'd53,8'd163} : s = 209;
	{8'd53,8'd164} : s = 357;
	{8'd53,8'd165} : s = 355;
	{8'd53,8'd166} : s = 467;
	{8'd53,8'd167} : s = 348;
	{8'd53,8'd168} : s = 462;
	{8'd53,8'd169} : s = 461;
	{8'd53,8'd170} : s = 505;
	{8'd53,8'd171} : s = 84;
	{8'd53,8'd172} : s = 204;
	{8'd53,8'd173} : s = 202;
	{8'd53,8'd174} : s = 346;
	{8'd53,8'd175} : s = 201;
	{8'd53,8'd176} : s = 345;
	{8'd53,8'd177} : s = 342;
	{8'd53,8'd178} : s = 459;
	{8'd53,8'd179} : s = 198;
	{8'd53,8'd180} : s = 341;
	{8'd53,8'd181} : s = 339;
	{8'd53,8'd182} : s = 455;
	{8'd53,8'd183} : s = 334;
	{8'd53,8'd184} : s = 444;
	{8'd53,8'd185} : s = 442;
	{8'd53,8'd186} : s = 502;
	{8'd53,8'd187} : s = 197;
	{8'd53,8'd188} : s = 333;
	{8'd53,8'd189} : s = 331;
	{8'd53,8'd190} : s = 441;
	{8'd53,8'd191} : s = 327;
	{8'd53,8'd192} : s = 438;
	{8'd53,8'd193} : s = 437;
	{8'd53,8'd194} : s = 501;
	{8'd53,8'd195} : s = 316;
	{8'd53,8'd196} : s = 435;
	{8'd53,8'd197} : s = 430;
	{8'd53,8'd198} : s = 499;
	{8'd53,8'd199} : s = 429;
	{8'd53,8'd200} : s = 494;
	{8'd53,8'd201} : s = 493;
	{8'd53,8'd202} : s = 510;
	{8'd53,8'd203} : s = 1;
	{8'd53,8'd204} : s = 18;
	{8'd53,8'd205} : s = 17;
	{8'd53,8'd206} : s = 82;
	{8'd53,8'd207} : s = 12;
	{8'd53,8'd208} : s = 81;
	{8'd53,8'd209} : s = 76;
	{8'd53,8'd210} : s = 195;
	{8'd53,8'd211} : s = 10;
	{8'd53,8'd212} : s = 74;
	{8'd53,8'd213} : s = 73;
	{8'd53,8'd214} : s = 184;
	{8'd53,8'd215} : s = 70;
	{8'd53,8'd216} : s = 180;
	{8'd53,8'd217} : s = 178;
	{8'd53,8'd218} : s = 314;
	{8'd53,8'd219} : s = 9;
	{8'd53,8'd220} : s = 69;
	{8'd53,8'd221} : s = 67;
	{8'd53,8'd222} : s = 177;
	{8'd53,8'd223} : s = 56;
	{8'd53,8'd224} : s = 172;
	{8'd53,8'd225} : s = 170;
	{8'd53,8'd226} : s = 313;
	{8'd53,8'd227} : s = 52;
	{8'd53,8'd228} : s = 169;
	{8'd53,8'd229} : s = 166;
	{8'd53,8'd230} : s = 310;
	{8'd53,8'd231} : s = 165;
	{8'd53,8'd232} : s = 309;
	{8'd53,8'd233} : s = 307;
	{8'd53,8'd234} : s = 427;
	{8'd53,8'd235} : s = 6;
	{8'd53,8'd236} : s = 50;
	{8'd53,8'd237} : s = 49;
	{8'd53,8'd238} : s = 163;
	{8'd53,8'd239} : s = 44;
	{8'd53,8'd240} : s = 156;
	{8'd53,8'd241} : s = 154;
	{8'd53,8'd242} : s = 302;
	{8'd53,8'd243} : s = 42;
	{8'd53,8'd244} : s = 153;
	{8'd53,8'd245} : s = 150;
	{8'd53,8'd246} : s = 301;
	{8'd53,8'd247} : s = 149;
	{8'd53,8'd248} : s = 299;
	{8'd53,8'd249} : s = 295;
	{8'd53,8'd250} : s = 423;
	{8'd53,8'd251} : s = 41;
	{8'd53,8'd252} : s = 147;
	{8'd53,8'd253} : s = 142;
	{8'd53,8'd254} : s = 286;
	{8'd53,8'd255} : s = 141;
	{8'd54,8'd0} : s = 408;
	{8'd54,8'd1} : s = 484;
	{8'd54,8'd2} : s = 276;
	{8'd54,8'd3} : s = 404;
	{8'd54,8'd4} : s = 402;
	{8'd54,8'd5} : s = 482;
	{8'd54,8'd6} : s = 401;
	{8'd54,8'd7} : s = 481;
	{8'd54,8'd8} : s = 472;
	{8'd54,8'd9} : s = 504;
	{8'd54,8'd10} : s = 4;
	{8'd54,8'd11} : s = 96;
	{8'd54,8'd12} : s = 80;
	{8'd54,8'd13} : s = 274;
	{8'd54,8'd14} : s = 72;
	{8'd54,8'd15} : s = 273;
	{8'd54,8'd16} : s = 268;
	{8'd54,8'd17} : s = 396;
	{8'd54,8'd18} : s = 68;
	{8'd54,8'd19} : s = 266;
	{8'd54,8'd20} : s = 265;
	{8'd54,8'd21} : s = 394;
	{8'd54,8'd22} : s = 262;
	{8'd54,8'd23} : s = 393;
	{8'd54,8'd24} : s = 390;
	{8'd54,8'd25} : s = 468;
	{8'd54,8'd26} : s = 66;
	{8'd54,8'd27} : s = 261;
	{8'd54,8'd28} : s = 259;
	{8'd54,8'd29} : s = 389;
	{8'd54,8'd30} : s = 224;
	{8'd54,8'd31} : s = 387;
	{8'd54,8'd32} : s = 368;
	{8'd54,8'd33} : s = 466;
	{8'd54,8'd34} : s = 208;
	{8'd54,8'd35} : s = 360;
	{8'd54,8'd36} : s = 356;
	{8'd54,8'd37} : s = 465;
	{8'd54,8'd38} : s = 354;
	{8'd54,8'd39} : s = 460;
	{8'd54,8'd40} : s = 458;
	{8'd54,8'd41} : s = 500;
	{8'd54,8'd42} : s = 65;
	{8'd54,8'd43} : s = 200;
	{8'd54,8'd44} : s = 196;
	{8'd54,8'd45} : s = 353;
	{8'd54,8'd46} : s = 194;
	{8'd54,8'd47} : s = 344;
	{8'd54,8'd48} : s = 340;
	{8'd54,8'd49} : s = 457;
	{8'd54,8'd50} : s = 193;
	{8'd54,8'd51} : s = 338;
	{8'd54,8'd52} : s = 337;
	{8'd54,8'd53} : s = 454;
	{8'd54,8'd54} : s = 332;
	{8'd54,8'd55} : s = 453;
	{8'd54,8'd56} : s = 451;
	{8'd54,8'd57} : s = 498;
	{8'd54,8'd58} : s = 176;
	{8'd54,8'd59} : s = 330;
	{8'd54,8'd60} : s = 329;
	{8'd54,8'd61} : s = 440;
	{8'd54,8'd62} : s = 326;
	{8'd54,8'd63} : s = 436;
	{8'd54,8'd64} : s = 434;
	{8'd54,8'd65} : s = 497;
	{8'd54,8'd66} : s = 325;
	{8'd54,8'd67} : s = 433;
	{8'd54,8'd68} : s = 428;
	{8'd54,8'd69} : s = 492;
	{8'd54,8'd70} : s = 426;
	{8'd54,8'd71} : s = 490;
	{8'd54,8'd72} : s = 489;
	{8'd54,8'd73} : s = 508;
	{8'd54,8'd74} : s = 2;
	{8'd54,8'd75} : s = 48;
	{8'd54,8'd76} : s = 40;
	{8'd54,8'd77} : s = 168;
	{8'd54,8'd78} : s = 36;
	{8'd54,8'd79} : s = 164;
	{8'd54,8'd80} : s = 162;
	{8'd54,8'd81} : s = 323;
	{8'd54,8'd82} : s = 34;
	{8'd54,8'd83} : s = 161;
	{8'd54,8'd84} : s = 152;
	{8'd54,8'd85} : s = 312;
	{8'd54,8'd86} : s = 148;
	{8'd54,8'd87} : s = 308;
	{8'd54,8'd88} : s = 306;
	{8'd54,8'd89} : s = 425;
	{8'd54,8'd90} : s = 33;
	{8'd54,8'd91} : s = 146;
	{8'd54,8'd92} : s = 145;
	{8'd54,8'd93} : s = 305;
	{8'd54,8'd94} : s = 140;
	{8'd54,8'd95} : s = 300;
	{8'd54,8'd96} : s = 298;
	{8'd54,8'd97} : s = 422;
	{8'd54,8'd98} : s = 138;
	{8'd54,8'd99} : s = 297;
	{8'd54,8'd100} : s = 294;
	{8'd54,8'd101} : s = 421;
	{8'd54,8'd102} : s = 293;
	{8'd54,8'd103} : s = 419;
	{8'd54,8'd104} : s = 412;
	{8'd54,8'd105} : s = 486;
	{8'd54,8'd106} : s = 24;
	{8'd54,8'd107} : s = 137;
	{8'd54,8'd108} : s = 134;
	{8'd54,8'd109} : s = 291;
	{8'd54,8'd110} : s = 133;
	{8'd54,8'd111} : s = 284;
	{8'd54,8'd112} : s = 282;
	{8'd54,8'd113} : s = 410;
	{8'd54,8'd114} : s = 131;
	{8'd54,8'd115} : s = 281;
	{8'd54,8'd116} : s = 278;
	{8'd54,8'd117} : s = 409;
	{8'd54,8'd118} : s = 277;
	{8'd54,8'd119} : s = 406;
	{8'd54,8'd120} : s = 405;
	{8'd54,8'd121} : s = 485;
	{8'd54,8'd122} : s = 112;
	{8'd54,8'd123} : s = 275;
	{8'd54,8'd124} : s = 270;
	{8'd54,8'd125} : s = 403;
	{8'd54,8'd126} : s = 269;
	{8'd54,8'd127} : s = 398;
	{8'd54,8'd128} : s = 397;
	{8'd54,8'd129} : s = 483;
	{8'd54,8'd130} : s = 267;
	{8'd54,8'd131} : s = 395;
	{8'd54,8'd132} : s = 391;
	{8'd54,8'd133} : s = 476;
	{8'd54,8'd134} : s = 376;
	{8'd54,8'd135} : s = 474;
	{8'd54,8'd136} : s = 473;
	{8'd54,8'd137} : s = 506;
	{8'd54,8'd138} : s = 20;
	{8'd54,8'd139} : s = 104;
	{8'd54,8'd140} : s = 100;
	{8'd54,8'd141} : s = 263;
	{8'd54,8'd142} : s = 98;
	{8'd54,8'd143} : s = 240;
	{8'd54,8'd144} : s = 232;
	{8'd54,8'd145} : s = 372;
	{8'd54,8'd146} : s = 97;
	{8'd54,8'd147} : s = 228;
	{8'd54,8'd148} : s = 226;
	{8'd54,8'd149} : s = 370;
	{8'd54,8'd150} : s = 225;
	{8'd54,8'd151} : s = 369;
	{8'd54,8'd152} : s = 364;
	{8'd54,8'd153} : s = 470;
	{8'd54,8'd154} : s = 88;
	{8'd54,8'd155} : s = 216;
	{8'd54,8'd156} : s = 212;
	{8'd54,8'd157} : s = 362;
	{8'd54,8'd158} : s = 210;
	{8'd54,8'd159} : s = 361;
	{8'd54,8'd160} : s = 358;
	{8'd54,8'd161} : s = 469;
	{8'd54,8'd162} : s = 209;
	{8'd54,8'd163} : s = 357;
	{8'd54,8'd164} : s = 355;
	{8'd54,8'd165} : s = 467;
	{8'd54,8'd166} : s = 348;
	{8'd54,8'd167} : s = 462;
	{8'd54,8'd168} : s = 461;
	{8'd54,8'd169} : s = 505;
	{8'd54,8'd170} : s = 84;
	{8'd54,8'd171} : s = 204;
	{8'd54,8'd172} : s = 202;
	{8'd54,8'd173} : s = 346;
	{8'd54,8'd174} : s = 201;
	{8'd54,8'd175} : s = 345;
	{8'd54,8'd176} : s = 342;
	{8'd54,8'd177} : s = 459;
	{8'd54,8'd178} : s = 198;
	{8'd54,8'd179} : s = 341;
	{8'd54,8'd180} : s = 339;
	{8'd54,8'd181} : s = 455;
	{8'd54,8'd182} : s = 334;
	{8'd54,8'd183} : s = 444;
	{8'd54,8'd184} : s = 442;
	{8'd54,8'd185} : s = 502;
	{8'd54,8'd186} : s = 197;
	{8'd54,8'd187} : s = 333;
	{8'd54,8'd188} : s = 331;
	{8'd54,8'd189} : s = 441;
	{8'd54,8'd190} : s = 327;
	{8'd54,8'd191} : s = 438;
	{8'd54,8'd192} : s = 437;
	{8'd54,8'd193} : s = 501;
	{8'd54,8'd194} : s = 316;
	{8'd54,8'd195} : s = 435;
	{8'd54,8'd196} : s = 430;
	{8'd54,8'd197} : s = 499;
	{8'd54,8'd198} : s = 429;
	{8'd54,8'd199} : s = 494;
	{8'd54,8'd200} : s = 493;
	{8'd54,8'd201} : s = 510;
	{8'd54,8'd202} : s = 1;
	{8'd54,8'd203} : s = 18;
	{8'd54,8'd204} : s = 17;
	{8'd54,8'd205} : s = 82;
	{8'd54,8'd206} : s = 12;
	{8'd54,8'd207} : s = 81;
	{8'd54,8'd208} : s = 76;
	{8'd54,8'd209} : s = 195;
	{8'd54,8'd210} : s = 10;
	{8'd54,8'd211} : s = 74;
	{8'd54,8'd212} : s = 73;
	{8'd54,8'd213} : s = 184;
	{8'd54,8'd214} : s = 70;
	{8'd54,8'd215} : s = 180;
	{8'd54,8'd216} : s = 178;
	{8'd54,8'd217} : s = 314;
	{8'd54,8'd218} : s = 9;
	{8'd54,8'd219} : s = 69;
	{8'd54,8'd220} : s = 67;
	{8'd54,8'd221} : s = 177;
	{8'd54,8'd222} : s = 56;
	{8'd54,8'd223} : s = 172;
	{8'd54,8'd224} : s = 170;
	{8'd54,8'd225} : s = 313;
	{8'd54,8'd226} : s = 52;
	{8'd54,8'd227} : s = 169;
	{8'd54,8'd228} : s = 166;
	{8'd54,8'd229} : s = 310;
	{8'd54,8'd230} : s = 165;
	{8'd54,8'd231} : s = 309;
	{8'd54,8'd232} : s = 307;
	{8'd54,8'd233} : s = 427;
	{8'd54,8'd234} : s = 6;
	{8'd54,8'd235} : s = 50;
	{8'd54,8'd236} : s = 49;
	{8'd54,8'd237} : s = 163;
	{8'd54,8'd238} : s = 44;
	{8'd54,8'd239} : s = 156;
	{8'd54,8'd240} : s = 154;
	{8'd54,8'd241} : s = 302;
	{8'd54,8'd242} : s = 42;
	{8'd54,8'd243} : s = 153;
	{8'd54,8'd244} : s = 150;
	{8'd54,8'd245} : s = 301;
	{8'd54,8'd246} : s = 149;
	{8'd54,8'd247} : s = 299;
	{8'd54,8'd248} : s = 295;
	{8'd54,8'd249} : s = 423;
	{8'd54,8'd250} : s = 41;
	{8'd54,8'd251} : s = 147;
	{8'd54,8'd252} : s = 142;
	{8'd54,8'd253} : s = 286;
	{8'd54,8'd254} : s = 141;
	{8'd54,8'd255} : s = 285;
	{8'd55,8'd0} : s = 484;
	{8'd55,8'd1} : s = 276;
	{8'd55,8'd2} : s = 404;
	{8'd55,8'd3} : s = 402;
	{8'd55,8'd4} : s = 482;
	{8'd55,8'd5} : s = 401;
	{8'd55,8'd6} : s = 481;
	{8'd55,8'd7} : s = 472;
	{8'd55,8'd8} : s = 504;
	{8'd55,8'd9} : s = 4;
	{8'd55,8'd10} : s = 96;
	{8'd55,8'd11} : s = 80;
	{8'd55,8'd12} : s = 274;
	{8'd55,8'd13} : s = 72;
	{8'd55,8'd14} : s = 273;
	{8'd55,8'd15} : s = 268;
	{8'd55,8'd16} : s = 396;
	{8'd55,8'd17} : s = 68;
	{8'd55,8'd18} : s = 266;
	{8'd55,8'd19} : s = 265;
	{8'd55,8'd20} : s = 394;
	{8'd55,8'd21} : s = 262;
	{8'd55,8'd22} : s = 393;
	{8'd55,8'd23} : s = 390;
	{8'd55,8'd24} : s = 468;
	{8'd55,8'd25} : s = 66;
	{8'd55,8'd26} : s = 261;
	{8'd55,8'd27} : s = 259;
	{8'd55,8'd28} : s = 389;
	{8'd55,8'd29} : s = 224;
	{8'd55,8'd30} : s = 387;
	{8'd55,8'd31} : s = 368;
	{8'd55,8'd32} : s = 466;
	{8'd55,8'd33} : s = 208;
	{8'd55,8'd34} : s = 360;
	{8'd55,8'd35} : s = 356;
	{8'd55,8'd36} : s = 465;
	{8'd55,8'd37} : s = 354;
	{8'd55,8'd38} : s = 460;
	{8'd55,8'd39} : s = 458;
	{8'd55,8'd40} : s = 500;
	{8'd55,8'd41} : s = 65;
	{8'd55,8'd42} : s = 200;
	{8'd55,8'd43} : s = 196;
	{8'd55,8'd44} : s = 353;
	{8'd55,8'd45} : s = 194;
	{8'd55,8'd46} : s = 344;
	{8'd55,8'd47} : s = 340;
	{8'd55,8'd48} : s = 457;
	{8'd55,8'd49} : s = 193;
	{8'd55,8'd50} : s = 338;
	{8'd55,8'd51} : s = 337;
	{8'd55,8'd52} : s = 454;
	{8'd55,8'd53} : s = 332;
	{8'd55,8'd54} : s = 453;
	{8'd55,8'd55} : s = 451;
	{8'd55,8'd56} : s = 498;
	{8'd55,8'd57} : s = 176;
	{8'd55,8'd58} : s = 330;
	{8'd55,8'd59} : s = 329;
	{8'd55,8'd60} : s = 440;
	{8'd55,8'd61} : s = 326;
	{8'd55,8'd62} : s = 436;
	{8'd55,8'd63} : s = 434;
	{8'd55,8'd64} : s = 497;
	{8'd55,8'd65} : s = 325;
	{8'd55,8'd66} : s = 433;
	{8'd55,8'd67} : s = 428;
	{8'd55,8'd68} : s = 492;
	{8'd55,8'd69} : s = 426;
	{8'd55,8'd70} : s = 490;
	{8'd55,8'd71} : s = 489;
	{8'd55,8'd72} : s = 508;
	{8'd55,8'd73} : s = 2;
	{8'd55,8'd74} : s = 48;
	{8'd55,8'd75} : s = 40;
	{8'd55,8'd76} : s = 168;
	{8'd55,8'd77} : s = 36;
	{8'd55,8'd78} : s = 164;
	{8'd55,8'd79} : s = 162;
	{8'd55,8'd80} : s = 323;
	{8'd55,8'd81} : s = 34;
	{8'd55,8'd82} : s = 161;
	{8'd55,8'd83} : s = 152;
	{8'd55,8'd84} : s = 312;
	{8'd55,8'd85} : s = 148;
	{8'd55,8'd86} : s = 308;
	{8'd55,8'd87} : s = 306;
	{8'd55,8'd88} : s = 425;
	{8'd55,8'd89} : s = 33;
	{8'd55,8'd90} : s = 146;
	{8'd55,8'd91} : s = 145;
	{8'd55,8'd92} : s = 305;
	{8'd55,8'd93} : s = 140;
	{8'd55,8'd94} : s = 300;
	{8'd55,8'd95} : s = 298;
	{8'd55,8'd96} : s = 422;
	{8'd55,8'd97} : s = 138;
	{8'd55,8'd98} : s = 297;
	{8'd55,8'd99} : s = 294;
	{8'd55,8'd100} : s = 421;
	{8'd55,8'd101} : s = 293;
	{8'd55,8'd102} : s = 419;
	{8'd55,8'd103} : s = 412;
	{8'd55,8'd104} : s = 486;
	{8'd55,8'd105} : s = 24;
	{8'd55,8'd106} : s = 137;
	{8'd55,8'd107} : s = 134;
	{8'd55,8'd108} : s = 291;
	{8'd55,8'd109} : s = 133;
	{8'd55,8'd110} : s = 284;
	{8'd55,8'd111} : s = 282;
	{8'd55,8'd112} : s = 410;
	{8'd55,8'd113} : s = 131;
	{8'd55,8'd114} : s = 281;
	{8'd55,8'd115} : s = 278;
	{8'd55,8'd116} : s = 409;
	{8'd55,8'd117} : s = 277;
	{8'd55,8'd118} : s = 406;
	{8'd55,8'd119} : s = 405;
	{8'd55,8'd120} : s = 485;
	{8'd55,8'd121} : s = 112;
	{8'd55,8'd122} : s = 275;
	{8'd55,8'd123} : s = 270;
	{8'd55,8'd124} : s = 403;
	{8'd55,8'd125} : s = 269;
	{8'd55,8'd126} : s = 398;
	{8'd55,8'd127} : s = 397;
	{8'd55,8'd128} : s = 483;
	{8'd55,8'd129} : s = 267;
	{8'd55,8'd130} : s = 395;
	{8'd55,8'd131} : s = 391;
	{8'd55,8'd132} : s = 476;
	{8'd55,8'd133} : s = 376;
	{8'd55,8'd134} : s = 474;
	{8'd55,8'd135} : s = 473;
	{8'd55,8'd136} : s = 506;
	{8'd55,8'd137} : s = 20;
	{8'd55,8'd138} : s = 104;
	{8'd55,8'd139} : s = 100;
	{8'd55,8'd140} : s = 263;
	{8'd55,8'd141} : s = 98;
	{8'd55,8'd142} : s = 240;
	{8'd55,8'd143} : s = 232;
	{8'd55,8'd144} : s = 372;
	{8'd55,8'd145} : s = 97;
	{8'd55,8'd146} : s = 228;
	{8'd55,8'd147} : s = 226;
	{8'd55,8'd148} : s = 370;
	{8'd55,8'd149} : s = 225;
	{8'd55,8'd150} : s = 369;
	{8'd55,8'd151} : s = 364;
	{8'd55,8'd152} : s = 470;
	{8'd55,8'd153} : s = 88;
	{8'd55,8'd154} : s = 216;
	{8'd55,8'd155} : s = 212;
	{8'd55,8'd156} : s = 362;
	{8'd55,8'd157} : s = 210;
	{8'd55,8'd158} : s = 361;
	{8'd55,8'd159} : s = 358;
	{8'd55,8'd160} : s = 469;
	{8'd55,8'd161} : s = 209;
	{8'd55,8'd162} : s = 357;
	{8'd55,8'd163} : s = 355;
	{8'd55,8'd164} : s = 467;
	{8'd55,8'd165} : s = 348;
	{8'd55,8'd166} : s = 462;
	{8'd55,8'd167} : s = 461;
	{8'd55,8'd168} : s = 505;
	{8'd55,8'd169} : s = 84;
	{8'd55,8'd170} : s = 204;
	{8'd55,8'd171} : s = 202;
	{8'd55,8'd172} : s = 346;
	{8'd55,8'd173} : s = 201;
	{8'd55,8'd174} : s = 345;
	{8'd55,8'd175} : s = 342;
	{8'd55,8'd176} : s = 459;
	{8'd55,8'd177} : s = 198;
	{8'd55,8'd178} : s = 341;
	{8'd55,8'd179} : s = 339;
	{8'd55,8'd180} : s = 455;
	{8'd55,8'd181} : s = 334;
	{8'd55,8'd182} : s = 444;
	{8'd55,8'd183} : s = 442;
	{8'd55,8'd184} : s = 502;
	{8'd55,8'd185} : s = 197;
	{8'd55,8'd186} : s = 333;
	{8'd55,8'd187} : s = 331;
	{8'd55,8'd188} : s = 441;
	{8'd55,8'd189} : s = 327;
	{8'd55,8'd190} : s = 438;
	{8'd55,8'd191} : s = 437;
	{8'd55,8'd192} : s = 501;
	{8'd55,8'd193} : s = 316;
	{8'd55,8'd194} : s = 435;
	{8'd55,8'd195} : s = 430;
	{8'd55,8'd196} : s = 499;
	{8'd55,8'd197} : s = 429;
	{8'd55,8'd198} : s = 494;
	{8'd55,8'd199} : s = 493;
	{8'd55,8'd200} : s = 510;
	{8'd55,8'd201} : s = 1;
	{8'd55,8'd202} : s = 18;
	{8'd55,8'd203} : s = 17;
	{8'd55,8'd204} : s = 82;
	{8'd55,8'd205} : s = 12;
	{8'd55,8'd206} : s = 81;
	{8'd55,8'd207} : s = 76;
	{8'd55,8'd208} : s = 195;
	{8'd55,8'd209} : s = 10;
	{8'd55,8'd210} : s = 74;
	{8'd55,8'd211} : s = 73;
	{8'd55,8'd212} : s = 184;
	{8'd55,8'd213} : s = 70;
	{8'd55,8'd214} : s = 180;
	{8'd55,8'd215} : s = 178;
	{8'd55,8'd216} : s = 314;
	{8'd55,8'd217} : s = 9;
	{8'd55,8'd218} : s = 69;
	{8'd55,8'd219} : s = 67;
	{8'd55,8'd220} : s = 177;
	{8'd55,8'd221} : s = 56;
	{8'd55,8'd222} : s = 172;
	{8'd55,8'd223} : s = 170;
	{8'd55,8'd224} : s = 313;
	{8'd55,8'd225} : s = 52;
	{8'd55,8'd226} : s = 169;
	{8'd55,8'd227} : s = 166;
	{8'd55,8'd228} : s = 310;
	{8'd55,8'd229} : s = 165;
	{8'd55,8'd230} : s = 309;
	{8'd55,8'd231} : s = 307;
	{8'd55,8'd232} : s = 427;
	{8'd55,8'd233} : s = 6;
	{8'd55,8'd234} : s = 50;
	{8'd55,8'd235} : s = 49;
	{8'd55,8'd236} : s = 163;
	{8'd55,8'd237} : s = 44;
	{8'd55,8'd238} : s = 156;
	{8'd55,8'd239} : s = 154;
	{8'd55,8'd240} : s = 302;
	{8'd55,8'd241} : s = 42;
	{8'd55,8'd242} : s = 153;
	{8'd55,8'd243} : s = 150;
	{8'd55,8'd244} : s = 301;
	{8'd55,8'd245} : s = 149;
	{8'd55,8'd246} : s = 299;
	{8'd55,8'd247} : s = 295;
	{8'd55,8'd248} : s = 423;
	{8'd55,8'd249} : s = 41;
	{8'd55,8'd250} : s = 147;
	{8'd55,8'd251} : s = 142;
	{8'd55,8'd252} : s = 286;
	{8'd55,8'd253} : s = 141;
	{8'd55,8'd254} : s = 285;
	{8'd55,8'd255} : s = 283;
	{8'd56,8'd0} : s = 276;
	{8'd56,8'd1} : s = 404;
	{8'd56,8'd2} : s = 402;
	{8'd56,8'd3} : s = 482;
	{8'd56,8'd4} : s = 401;
	{8'd56,8'd5} : s = 481;
	{8'd56,8'd6} : s = 472;
	{8'd56,8'd7} : s = 504;
	{8'd56,8'd8} : s = 4;
	{8'd56,8'd9} : s = 96;
	{8'd56,8'd10} : s = 80;
	{8'd56,8'd11} : s = 274;
	{8'd56,8'd12} : s = 72;
	{8'd56,8'd13} : s = 273;
	{8'd56,8'd14} : s = 268;
	{8'd56,8'd15} : s = 396;
	{8'd56,8'd16} : s = 68;
	{8'd56,8'd17} : s = 266;
	{8'd56,8'd18} : s = 265;
	{8'd56,8'd19} : s = 394;
	{8'd56,8'd20} : s = 262;
	{8'd56,8'd21} : s = 393;
	{8'd56,8'd22} : s = 390;
	{8'd56,8'd23} : s = 468;
	{8'd56,8'd24} : s = 66;
	{8'd56,8'd25} : s = 261;
	{8'd56,8'd26} : s = 259;
	{8'd56,8'd27} : s = 389;
	{8'd56,8'd28} : s = 224;
	{8'd56,8'd29} : s = 387;
	{8'd56,8'd30} : s = 368;
	{8'd56,8'd31} : s = 466;
	{8'd56,8'd32} : s = 208;
	{8'd56,8'd33} : s = 360;
	{8'd56,8'd34} : s = 356;
	{8'd56,8'd35} : s = 465;
	{8'd56,8'd36} : s = 354;
	{8'd56,8'd37} : s = 460;
	{8'd56,8'd38} : s = 458;
	{8'd56,8'd39} : s = 500;
	{8'd56,8'd40} : s = 65;
	{8'd56,8'd41} : s = 200;
	{8'd56,8'd42} : s = 196;
	{8'd56,8'd43} : s = 353;
	{8'd56,8'd44} : s = 194;
	{8'd56,8'd45} : s = 344;
	{8'd56,8'd46} : s = 340;
	{8'd56,8'd47} : s = 457;
	{8'd56,8'd48} : s = 193;
	{8'd56,8'd49} : s = 338;
	{8'd56,8'd50} : s = 337;
	{8'd56,8'd51} : s = 454;
	{8'd56,8'd52} : s = 332;
	{8'd56,8'd53} : s = 453;
	{8'd56,8'd54} : s = 451;
	{8'd56,8'd55} : s = 498;
	{8'd56,8'd56} : s = 176;
	{8'd56,8'd57} : s = 330;
	{8'd56,8'd58} : s = 329;
	{8'd56,8'd59} : s = 440;
	{8'd56,8'd60} : s = 326;
	{8'd56,8'd61} : s = 436;
	{8'd56,8'd62} : s = 434;
	{8'd56,8'd63} : s = 497;
	{8'd56,8'd64} : s = 325;
	{8'd56,8'd65} : s = 433;
	{8'd56,8'd66} : s = 428;
	{8'd56,8'd67} : s = 492;
	{8'd56,8'd68} : s = 426;
	{8'd56,8'd69} : s = 490;
	{8'd56,8'd70} : s = 489;
	{8'd56,8'd71} : s = 508;
	{8'd56,8'd72} : s = 2;
	{8'd56,8'd73} : s = 48;
	{8'd56,8'd74} : s = 40;
	{8'd56,8'd75} : s = 168;
	{8'd56,8'd76} : s = 36;
	{8'd56,8'd77} : s = 164;
	{8'd56,8'd78} : s = 162;
	{8'd56,8'd79} : s = 323;
	{8'd56,8'd80} : s = 34;
	{8'd56,8'd81} : s = 161;
	{8'd56,8'd82} : s = 152;
	{8'd56,8'd83} : s = 312;
	{8'd56,8'd84} : s = 148;
	{8'd56,8'd85} : s = 308;
	{8'd56,8'd86} : s = 306;
	{8'd56,8'd87} : s = 425;
	{8'd56,8'd88} : s = 33;
	{8'd56,8'd89} : s = 146;
	{8'd56,8'd90} : s = 145;
	{8'd56,8'd91} : s = 305;
	{8'd56,8'd92} : s = 140;
	{8'd56,8'd93} : s = 300;
	{8'd56,8'd94} : s = 298;
	{8'd56,8'd95} : s = 422;
	{8'd56,8'd96} : s = 138;
	{8'd56,8'd97} : s = 297;
	{8'd56,8'd98} : s = 294;
	{8'd56,8'd99} : s = 421;
	{8'd56,8'd100} : s = 293;
	{8'd56,8'd101} : s = 419;
	{8'd56,8'd102} : s = 412;
	{8'd56,8'd103} : s = 486;
	{8'd56,8'd104} : s = 24;
	{8'd56,8'd105} : s = 137;
	{8'd56,8'd106} : s = 134;
	{8'd56,8'd107} : s = 291;
	{8'd56,8'd108} : s = 133;
	{8'd56,8'd109} : s = 284;
	{8'd56,8'd110} : s = 282;
	{8'd56,8'd111} : s = 410;
	{8'd56,8'd112} : s = 131;
	{8'd56,8'd113} : s = 281;
	{8'd56,8'd114} : s = 278;
	{8'd56,8'd115} : s = 409;
	{8'd56,8'd116} : s = 277;
	{8'd56,8'd117} : s = 406;
	{8'd56,8'd118} : s = 405;
	{8'd56,8'd119} : s = 485;
	{8'd56,8'd120} : s = 112;
	{8'd56,8'd121} : s = 275;
	{8'd56,8'd122} : s = 270;
	{8'd56,8'd123} : s = 403;
	{8'd56,8'd124} : s = 269;
	{8'd56,8'd125} : s = 398;
	{8'd56,8'd126} : s = 397;
	{8'd56,8'd127} : s = 483;
	{8'd56,8'd128} : s = 267;
	{8'd56,8'd129} : s = 395;
	{8'd56,8'd130} : s = 391;
	{8'd56,8'd131} : s = 476;
	{8'd56,8'd132} : s = 376;
	{8'd56,8'd133} : s = 474;
	{8'd56,8'd134} : s = 473;
	{8'd56,8'd135} : s = 506;
	{8'd56,8'd136} : s = 20;
	{8'd56,8'd137} : s = 104;
	{8'd56,8'd138} : s = 100;
	{8'd56,8'd139} : s = 263;
	{8'd56,8'd140} : s = 98;
	{8'd56,8'd141} : s = 240;
	{8'd56,8'd142} : s = 232;
	{8'd56,8'd143} : s = 372;
	{8'd56,8'd144} : s = 97;
	{8'd56,8'd145} : s = 228;
	{8'd56,8'd146} : s = 226;
	{8'd56,8'd147} : s = 370;
	{8'd56,8'd148} : s = 225;
	{8'd56,8'd149} : s = 369;
	{8'd56,8'd150} : s = 364;
	{8'd56,8'd151} : s = 470;
	{8'd56,8'd152} : s = 88;
	{8'd56,8'd153} : s = 216;
	{8'd56,8'd154} : s = 212;
	{8'd56,8'd155} : s = 362;
	{8'd56,8'd156} : s = 210;
	{8'd56,8'd157} : s = 361;
	{8'd56,8'd158} : s = 358;
	{8'd56,8'd159} : s = 469;
	{8'd56,8'd160} : s = 209;
	{8'd56,8'd161} : s = 357;
	{8'd56,8'd162} : s = 355;
	{8'd56,8'd163} : s = 467;
	{8'd56,8'd164} : s = 348;
	{8'd56,8'd165} : s = 462;
	{8'd56,8'd166} : s = 461;
	{8'd56,8'd167} : s = 505;
	{8'd56,8'd168} : s = 84;
	{8'd56,8'd169} : s = 204;
	{8'd56,8'd170} : s = 202;
	{8'd56,8'd171} : s = 346;
	{8'd56,8'd172} : s = 201;
	{8'd56,8'd173} : s = 345;
	{8'd56,8'd174} : s = 342;
	{8'd56,8'd175} : s = 459;
	{8'd56,8'd176} : s = 198;
	{8'd56,8'd177} : s = 341;
	{8'd56,8'd178} : s = 339;
	{8'd56,8'd179} : s = 455;
	{8'd56,8'd180} : s = 334;
	{8'd56,8'd181} : s = 444;
	{8'd56,8'd182} : s = 442;
	{8'd56,8'd183} : s = 502;
	{8'd56,8'd184} : s = 197;
	{8'd56,8'd185} : s = 333;
	{8'd56,8'd186} : s = 331;
	{8'd56,8'd187} : s = 441;
	{8'd56,8'd188} : s = 327;
	{8'd56,8'd189} : s = 438;
	{8'd56,8'd190} : s = 437;
	{8'd56,8'd191} : s = 501;
	{8'd56,8'd192} : s = 316;
	{8'd56,8'd193} : s = 435;
	{8'd56,8'd194} : s = 430;
	{8'd56,8'd195} : s = 499;
	{8'd56,8'd196} : s = 429;
	{8'd56,8'd197} : s = 494;
	{8'd56,8'd198} : s = 493;
	{8'd56,8'd199} : s = 510;
	{8'd56,8'd200} : s = 1;
	{8'd56,8'd201} : s = 18;
	{8'd56,8'd202} : s = 17;
	{8'd56,8'd203} : s = 82;
	{8'd56,8'd204} : s = 12;
	{8'd56,8'd205} : s = 81;
	{8'd56,8'd206} : s = 76;
	{8'd56,8'd207} : s = 195;
	{8'd56,8'd208} : s = 10;
	{8'd56,8'd209} : s = 74;
	{8'd56,8'd210} : s = 73;
	{8'd56,8'd211} : s = 184;
	{8'd56,8'd212} : s = 70;
	{8'd56,8'd213} : s = 180;
	{8'd56,8'd214} : s = 178;
	{8'd56,8'd215} : s = 314;
	{8'd56,8'd216} : s = 9;
	{8'd56,8'd217} : s = 69;
	{8'd56,8'd218} : s = 67;
	{8'd56,8'd219} : s = 177;
	{8'd56,8'd220} : s = 56;
	{8'd56,8'd221} : s = 172;
	{8'd56,8'd222} : s = 170;
	{8'd56,8'd223} : s = 313;
	{8'd56,8'd224} : s = 52;
	{8'd56,8'd225} : s = 169;
	{8'd56,8'd226} : s = 166;
	{8'd56,8'd227} : s = 310;
	{8'd56,8'd228} : s = 165;
	{8'd56,8'd229} : s = 309;
	{8'd56,8'd230} : s = 307;
	{8'd56,8'd231} : s = 427;
	{8'd56,8'd232} : s = 6;
	{8'd56,8'd233} : s = 50;
	{8'd56,8'd234} : s = 49;
	{8'd56,8'd235} : s = 163;
	{8'd56,8'd236} : s = 44;
	{8'd56,8'd237} : s = 156;
	{8'd56,8'd238} : s = 154;
	{8'd56,8'd239} : s = 302;
	{8'd56,8'd240} : s = 42;
	{8'd56,8'd241} : s = 153;
	{8'd56,8'd242} : s = 150;
	{8'd56,8'd243} : s = 301;
	{8'd56,8'd244} : s = 149;
	{8'd56,8'd245} : s = 299;
	{8'd56,8'd246} : s = 295;
	{8'd56,8'd247} : s = 423;
	{8'd56,8'd248} : s = 41;
	{8'd56,8'd249} : s = 147;
	{8'd56,8'd250} : s = 142;
	{8'd56,8'd251} : s = 286;
	{8'd56,8'd252} : s = 141;
	{8'd56,8'd253} : s = 285;
	{8'd56,8'd254} : s = 283;
	{8'd56,8'd255} : s = 414;
	{8'd57,8'd0} : s = 404;
	{8'd57,8'd1} : s = 402;
	{8'd57,8'd2} : s = 482;
	{8'd57,8'd3} : s = 401;
	{8'd57,8'd4} : s = 481;
	{8'd57,8'd5} : s = 472;
	{8'd57,8'd6} : s = 504;
	{8'd57,8'd7} : s = 4;
	{8'd57,8'd8} : s = 96;
	{8'd57,8'd9} : s = 80;
	{8'd57,8'd10} : s = 274;
	{8'd57,8'd11} : s = 72;
	{8'd57,8'd12} : s = 273;
	{8'd57,8'd13} : s = 268;
	{8'd57,8'd14} : s = 396;
	{8'd57,8'd15} : s = 68;
	{8'd57,8'd16} : s = 266;
	{8'd57,8'd17} : s = 265;
	{8'd57,8'd18} : s = 394;
	{8'd57,8'd19} : s = 262;
	{8'd57,8'd20} : s = 393;
	{8'd57,8'd21} : s = 390;
	{8'd57,8'd22} : s = 468;
	{8'd57,8'd23} : s = 66;
	{8'd57,8'd24} : s = 261;
	{8'd57,8'd25} : s = 259;
	{8'd57,8'd26} : s = 389;
	{8'd57,8'd27} : s = 224;
	{8'd57,8'd28} : s = 387;
	{8'd57,8'd29} : s = 368;
	{8'd57,8'd30} : s = 466;
	{8'd57,8'd31} : s = 208;
	{8'd57,8'd32} : s = 360;
	{8'd57,8'd33} : s = 356;
	{8'd57,8'd34} : s = 465;
	{8'd57,8'd35} : s = 354;
	{8'd57,8'd36} : s = 460;
	{8'd57,8'd37} : s = 458;
	{8'd57,8'd38} : s = 500;
	{8'd57,8'd39} : s = 65;
	{8'd57,8'd40} : s = 200;
	{8'd57,8'd41} : s = 196;
	{8'd57,8'd42} : s = 353;
	{8'd57,8'd43} : s = 194;
	{8'd57,8'd44} : s = 344;
	{8'd57,8'd45} : s = 340;
	{8'd57,8'd46} : s = 457;
	{8'd57,8'd47} : s = 193;
	{8'd57,8'd48} : s = 338;
	{8'd57,8'd49} : s = 337;
	{8'd57,8'd50} : s = 454;
	{8'd57,8'd51} : s = 332;
	{8'd57,8'd52} : s = 453;
	{8'd57,8'd53} : s = 451;
	{8'd57,8'd54} : s = 498;
	{8'd57,8'd55} : s = 176;
	{8'd57,8'd56} : s = 330;
	{8'd57,8'd57} : s = 329;
	{8'd57,8'd58} : s = 440;
	{8'd57,8'd59} : s = 326;
	{8'd57,8'd60} : s = 436;
	{8'd57,8'd61} : s = 434;
	{8'd57,8'd62} : s = 497;
	{8'd57,8'd63} : s = 325;
	{8'd57,8'd64} : s = 433;
	{8'd57,8'd65} : s = 428;
	{8'd57,8'd66} : s = 492;
	{8'd57,8'd67} : s = 426;
	{8'd57,8'd68} : s = 490;
	{8'd57,8'd69} : s = 489;
	{8'd57,8'd70} : s = 508;
	{8'd57,8'd71} : s = 2;
	{8'd57,8'd72} : s = 48;
	{8'd57,8'd73} : s = 40;
	{8'd57,8'd74} : s = 168;
	{8'd57,8'd75} : s = 36;
	{8'd57,8'd76} : s = 164;
	{8'd57,8'd77} : s = 162;
	{8'd57,8'd78} : s = 323;
	{8'd57,8'd79} : s = 34;
	{8'd57,8'd80} : s = 161;
	{8'd57,8'd81} : s = 152;
	{8'd57,8'd82} : s = 312;
	{8'd57,8'd83} : s = 148;
	{8'd57,8'd84} : s = 308;
	{8'd57,8'd85} : s = 306;
	{8'd57,8'd86} : s = 425;
	{8'd57,8'd87} : s = 33;
	{8'd57,8'd88} : s = 146;
	{8'd57,8'd89} : s = 145;
	{8'd57,8'd90} : s = 305;
	{8'd57,8'd91} : s = 140;
	{8'd57,8'd92} : s = 300;
	{8'd57,8'd93} : s = 298;
	{8'd57,8'd94} : s = 422;
	{8'd57,8'd95} : s = 138;
	{8'd57,8'd96} : s = 297;
	{8'd57,8'd97} : s = 294;
	{8'd57,8'd98} : s = 421;
	{8'd57,8'd99} : s = 293;
	{8'd57,8'd100} : s = 419;
	{8'd57,8'd101} : s = 412;
	{8'd57,8'd102} : s = 486;
	{8'd57,8'd103} : s = 24;
	{8'd57,8'd104} : s = 137;
	{8'd57,8'd105} : s = 134;
	{8'd57,8'd106} : s = 291;
	{8'd57,8'd107} : s = 133;
	{8'd57,8'd108} : s = 284;
	{8'd57,8'd109} : s = 282;
	{8'd57,8'd110} : s = 410;
	{8'd57,8'd111} : s = 131;
	{8'd57,8'd112} : s = 281;
	{8'd57,8'd113} : s = 278;
	{8'd57,8'd114} : s = 409;
	{8'd57,8'd115} : s = 277;
	{8'd57,8'd116} : s = 406;
	{8'd57,8'd117} : s = 405;
	{8'd57,8'd118} : s = 485;
	{8'd57,8'd119} : s = 112;
	{8'd57,8'd120} : s = 275;
	{8'd57,8'd121} : s = 270;
	{8'd57,8'd122} : s = 403;
	{8'd57,8'd123} : s = 269;
	{8'd57,8'd124} : s = 398;
	{8'd57,8'd125} : s = 397;
	{8'd57,8'd126} : s = 483;
	{8'd57,8'd127} : s = 267;
	{8'd57,8'd128} : s = 395;
	{8'd57,8'd129} : s = 391;
	{8'd57,8'd130} : s = 476;
	{8'd57,8'd131} : s = 376;
	{8'd57,8'd132} : s = 474;
	{8'd57,8'd133} : s = 473;
	{8'd57,8'd134} : s = 506;
	{8'd57,8'd135} : s = 20;
	{8'd57,8'd136} : s = 104;
	{8'd57,8'd137} : s = 100;
	{8'd57,8'd138} : s = 263;
	{8'd57,8'd139} : s = 98;
	{8'd57,8'd140} : s = 240;
	{8'd57,8'd141} : s = 232;
	{8'd57,8'd142} : s = 372;
	{8'd57,8'd143} : s = 97;
	{8'd57,8'd144} : s = 228;
	{8'd57,8'd145} : s = 226;
	{8'd57,8'd146} : s = 370;
	{8'd57,8'd147} : s = 225;
	{8'd57,8'd148} : s = 369;
	{8'd57,8'd149} : s = 364;
	{8'd57,8'd150} : s = 470;
	{8'd57,8'd151} : s = 88;
	{8'd57,8'd152} : s = 216;
	{8'd57,8'd153} : s = 212;
	{8'd57,8'd154} : s = 362;
	{8'd57,8'd155} : s = 210;
	{8'd57,8'd156} : s = 361;
	{8'd57,8'd157} : s = 358;
	{8'd57,8'd158} : s = 469;
	{8'd57,8'd159} : s = 209;
	{8'd57,8'd160} : s = 357;
	{8'd57,8'd161} : s = 355;
	{8'd57,8'd162} : s = 467;
	{8'd57,8'd163} : s = 348;
	{8'd57,8'd164} : s = 462;
	{8'd57,8'd165} : s = 461;
	{8'd57,8'd166} : s = 505;
	{8'd57,8'd167} : s = 84;
	{8'd57,8'd168} : s = 204;
	{8'd57,8'd169} : s = 202;
	{8'd57,8'd170} : s = 346;
	{8'd57,8'd171} : s = 201;
	{8'd57,8'd172} : s = 345;
	{8'd57,8'd173} : s = 342;
	{8'd57,8'd174} : s = 459;
	{8'd57,8'd175} : s = 198;
	{8'd57,8'd176} : s = 341;
	{8'd57,8'd177} : s = 339;
	{8'd57,8'd178} : s = 455;
	{8'd57,8'd179} : s = 334;
	{8'd57,8'd180} : s = 444;
	{8'd57,8'd181} : s = 442;
	{8'd57,8'd182} : s = 502;
	{8'd57,8'd183} : s = 197;
	{8'd57,8'd184} : s = 333;
	{8'd57,8'd185} : s = 331;
	{8'd57,8'd186} : s = 441;
	{8'd57,8'd187} : s = 327;
	{8'd57,8'd188} : s = 438;
	{8'd57,8'd189} : s = 437;
	{8'd57,8'd190} : s = 501;
	{8'd57,8'd191} : s = 316;
	{8'd57,8'd192} : s = 435;
	{8'd57,8'd193} : s = 430;
	{8'd57,8'd194} : s = 499;
	{8'd57,8'd195} : s = 429;
	{8'd57,8'd196} : s = 494;
	{8'd57,8'd197} : s = 493;
	{8'd57,8'd198} : s = 510;
	{8'd57,8'd199} : s = 1;
	{8'd57,8'd200} : s = 18;
	{8'd57,8'd201} : s = 17;
	{8'd57,8'd202} : s = 82;
	{8'd57,8'd203} : s = 12;
	{8'd57,8'd204} : s = 81;
	{8'd57,8'd205} : s = 76;
	{8'd57,8'd206} : s = 195;
	{8'd57,8'd207} : s = 10;
	{8'd57,8'd208} : s = 74;
	{8'd57,8'd209} : s = 73;
	{8'd57,8'd210} : s = 184;
	{8'd57,8'd211} : s = 70;
	{8'd57,8'd212} : s = 180;
	{8'd57,8'd213} : s = 178;
	{8'd57,8'd214} : s = 314;
	{8'd57,8'd215} : s = 9;
	{8'd57,8'd216} : s = 69;
	{8'd57,8'd217} : s = 67;
	{8'd57,8'd218} : s = 177;
	{8'd57,8'd219} : s = 56;
	{8'd57,8'd220} : s = 172;
	{8'd57,8'd221} : s = 170;
	{8'd57,8'd222} : s = 313;
	{8'd57,8'd223} : s = 52;
	{8'd57,8'd224} : s = 169;
	{8'd57,8'd225} : s = 166;
	{8'd57,8'd226} : s = 310;
	{8'd57,8'd227} : s = 165;
	{8'd57,8'd228} : s = 309;
	{8'd57,8'd229} : s = 307;
	{8'd57,8'd230} : s = 427;
	{8'd57,8'd231} : s = 6;
	{8'd57,8'd232} : s = 50;
	{8'd57,8'd233} : s = 49;
	{8'd57,8'd234} : s = 163;
	{8'd57,8'd235} : s = 44;
	{8'd57,8'd236} : s = 156;
	{8'd57,8'd237} : s = 154;
	{8'd57,8'd238} : s = 302;
	{8'd57,8'd239} : s = 42;
	{8'd57,8'd240} : s = 153;
	{8'd57,8'd241} : s = 150;
	{8'd57,8'd242} : s = 301;
	{8'd57,8'd243} : s = 149;
	{8'd57,8'd244} : s = 299;
	{8'd57,8'd245} : s = 295;
	{8'd57,8'd246} : s = 423;
	{8'd57,8'd247} : s = 41;
	{8'd57,8'd248} : s = 147;
	{8'd57,8'd249} : s = 142;
	{8'd57,8'd250} : s = 286;
	{8'd57,8'd251} : s = 141;
	{8'd57,8'd252} : s = 285;
	{8'd57,8'd253} : s = 283;
	{8'd57,8'd254} : s = 414;
	{8'd57,8'd255} : s = 139;
	{8'd58,8'd0} : s = 402;
	{8'd58,8'd1} : s = 482;
	{8'd58,8'd2} : s = 401;
	{8'd58,8'd3} : s = 481;
	{8'd58,8'd4} : s = 472;
	{8'd58,8'd5} : s = 504;
	{8'd58,8'd6} : s = 4;
	{8'd58,8'd7} : s = 96;
	{8'd58,8'd8} : s = 80;
	{8'd58,8'd9} : s = 274;
	{8'd58,8'd10} : s = 72;
	{8'd58,8'd11} : s = 273;
	{8'd58,8'd12} : s = 268;
	{8'd58,8'd13} : s = 396;
	{8'd58,8'd14} : s = 68;
	{8'd58,8'd15} : s = 266;
	{8'd58,8'd16} : s = 265;
	{8'd58,8'd17} : s = 394;
	{8'd58,8'd18} : s = 262;
	{8'd58,8'd19} : s = 393;
	{8'd58,8'd20} : s = 390;
	{8'd58,8'd21} : s = 468;
	{8'd58,8'd22} : s = 66;
	{8'd58,8'd23} : s = 261;
	{8'd58,8'd24} : s = 259;
	{8'd58,8'd25} : s = 389;
	{8'd58,8'd26} : s = 224;
	{8'd58,8'd27} : s = 387;
	{8'd58,8'd28} : s = 368;
	{8'd58,8'd29} : s = 466;
	{8'd58,8'd30} : s = 208;
	{8'd58,8'd31} : s = 360;
	{8'd58,8'd32} : s = 356;
	{8'd58,8'd33} : s = 465;
	{8'd58,8'd34} : s = 354;
	{8'd58,8'd35} : s = 460;
	{8'd58,8'd36} : s = 458;
	{8'd58,8'd37} : s = 500;
	{8'd58,8'd38} : s = 65;
	{8'd58,8'd39} : s = 200;
	{8'd58,8'd40} : s = 196;
	{8'd58,8'd41} : s = 353;
	{8'd58,8'd42} : s = 194;
	{8'd58,8'd43} : s = 344;
	{8'd58,8'd44} : s = 340;
	{8'd58,8'd45} : s = 457;
	{8'd58,8'd46} : s = 193;
	{8'd58,8'd47} : s = 338;
	{8'd58,8'd48} : s = 337;
	{8'd58,8'd49} : s = 454;
	{8'd58,8'd50} : s = 332;
	{8'd58,8'd51} : s = 453;
	{8'd58,8'd52} : s = 451;
	{8'd58,8'd53} : s = 498;
	{8'd58,8'd54} : s = 176;
	{8'd58,8'd55} : s = 330;
	{8'd58,8'd56} : s = 329;
	{8'd58,8'd57} : s = 440;
	{8'd58,8'd58} : s = 326;
	{8'd58,8'd59} : s = 436;
	{8'd58,8'd60} : s = 434;
	{8'd58,8'd61} : s = 497;
	{8'd58,8'd62} : s = 325;
	{8'd58,8'd63} : s = 433;
	{8'd58,8'd64} : s = 428;
	{8'd58,8'd65} : s = 492;
	{8'd58,8'd66} : s = 426;
	{8'd58,8'd67} : s = 490;
	{8'd58,8'd68} : s = 489;
	{8'd58,8'd69} : s = 508;
	{8'd58,8'd70} : s = 2;
	{8'd58,8'd71} : s = 48;
	{8'd58,8'd72} : s = 40;
	{8'd58,8'd73} : s = 168;
	{8'd58,8'd74} : s = 36;
	{8'd58,8'd75} : s = 164;
	{8'd58,8'd76} : s = 162;
	{8'd58,8'd77} : s = 323;
	{8'd58,8'd78} : s = 34;
	{8'd58,8'd79} : s = 161;
	{8'd58,8'd80} : s = 152;
	{8'd58,8'd81} : s = 312;
	{8'd58,8'd82} : s = 148;
	{8'd58,8'd83} : s = 308;
	{8'd58,8'd84} : s = 306;
	{8'd58,8'd85} : s = 425;
	{8'd58,8'd86} : s = 33;
	{8'd58,8'd87} : s = 146;
	{8'd58,8'd88} : s = 145;
	{8'd58,8'd89} : s = 305;
	{8'd58,8'd90} : s = 140;
	{8'd58,8'd91} : s = 300;
	{8'd58,8'd92} : s = 298;
	{8'd58,8'd93} : s = 422;
	{8'd58,8'd94} : s = 138;
	{8'd58,8'd95} : s = 297;
	{8'd58,8'd96} : s = 294;
	{8'd58,8'd97} : s = 421;
	{8'd58,8'd98} : s = 293;
	{8'd58,8'd99} : s = 419;
	{8'd58,8'd100} : s = 412;
	{8'd58,8'd101} : s = 486;
	{8'd58,8'd102} : s = 24;
	{8'd58,8'd103} : s = 137;
	{8'd58,8'd104} : s = 134;
	{8'd58,8'd105} : s = 291;
	{8'd58,8'd106} : s = 133;
	{8'd58,8'd107} : s = 284;
	{8'd58,8'd108} : s = 282;
	{8'd58,8'd109} : s = 410;
	{8'd58,8'd110} : s = 131;
	{8'd58,8'd111} : s = 281;
	{8'd58,8'd112} : s = 278;
	{8'd58,8'd113} : s = 409;
	{8'd58,8'd114} : s = 277;
	{8'd58,8'd115} : s = 406;
	{8'd58,8'd116} : s = 405;
	{8'd58,8'd117} : s = 485;
	{8'd58,8'd118} : s = 112;
	{8'd58,8'd119} : s = 275;
	{8'd58,8'd120} : s = 270;
	{8'd58,8'd121} : s = 403;
	{8'd58,8'd122} : s = 269;
	{8'd58,8'd123} : s = 398;
	{8'd58,8'd124} : s = 397;
	{8'd58,8'd125} : s = 483;
	{8'd58,8'd126} : s = 267;
	{8'd58,8'd127} : s = 395;
	{8'd58,8'd128} : s = 391;
	{8'd58,8'd129} : s = 476;
	{8'd58,8'd130} : s = 376;
	{8'd58,8'd131} : s = 474;
	{8'd58,8'd132} : s = 473;
	{8'd58,8'd133} : s = 506;
	{8'd58,8'd134} : s = 20;
	{8'd58,8'd135} : s = 104;
	{8'd58,8'd136} : s = 100;
	{8'd58,8'd137} : s = 263;
	{8'd58,8'd138} : s = 98;
	{8'd58,8'd139} : s = 240;
	{8'd58,8'd140} : s = 232;
	{8'd58,8'd141} : s = 372;
	{8'd58,8'd142} : s = 97;
	{8'd58,8'd143} : s = 228;
	{8'd58,8'd144} : s = 226;
	{8'd58,8'd145} : s = 370;
	{8'd58,8'd146} : s = 225;
	{8'd58,8'd147} : s = 369;
	{8'd58,8'd148} : s = 364;
	{8'd58,8'd149} : s = 470;
	{8'd58,8'd150} : s = 88;
	{8'd58,8'd151} : s = 216;
	{8'd58,8'd152} : s = 212;
	{8'd58,8'd153} : s = 362;
	{8'd58,8'd154} : s = 210;
	{8'd58,8'd155} : s = 361;
	{8'd58,8'd156} : s = 358;
	{8'd58,8'd157} : s = 469;
	{8'd58,8'd158} : s = 209;
	{8'd58,8'd159} : s = 357;
	{8'd58,8'd160} : s = 355;
	{8'd58,8'd161} : s = 467;
	{8'd58,8'd162} : s = 348;
	{8'd58,8'd163} : s = 462;
	{8'd58,8'd164} : s = 461;
	{8'd58,8'd165} : s = 505;
	{8'd58,8'd166} : s = 84;
	{8'd58,8'd167} : s = 204;
	{8'd58,8'd168} : s = 202;
	{8'd58,8'd169} : s = 346;
	{8'd58,8'd170} : s = 201;
	{8'd58,8'd171} : s = 345;
	{8'd58,8'd172} : s = 342;
	{8'd58,8'd173} : s = 459;
	{8'd58,8'd174} : s = 198;
	{8'd58,8'd175} : s = 341;
	{8'd58,8'd176} : s = 339;
	{8'd58,8'd177} : s = 455;
	{8'd58,8'd178} : s = 334;
	{8'd58,8'd179} : s = 444;
	{8'd58,8'd180} : s = 442;
	{8'd58,8'd181} : s = 502;
	{8'd58,8'd182} : s = 197;
	{8'd58,8'd183} : s = 333;
	{8'd58,8'd184} : s = 331;
	{8'd58,8'd185} : s = 441;
	{8'd58,8'd186} : s = 327;
	{8'd58,8'd187} : s = 438;
	{8'd58,8'd188} : s = 437;
	{8'd58,8'd189} : s = 501;
	{8'd58,8'd190} : s = 316;
	{8'd58,8'd191} : s = 435;
	{8'd58,8'd192} : s = 430;
	{8'd58,8'd193} : s = 499;
	{8'd58,8'd194} : s = 429;
	{8'd58,8'd195} : s = 494;
	{8'd58,8'd196} : s = 493;
	{8'd58,8'd197} : s = 510;
	{8'd58,8'd198} : s = 1;
	{8'd58,8'd199} : s = 18;
	{8'd58,8'd200} : s = 17;
	{8'd58,8'd201} : s = 82;
	{8'd58,8'd202} : s = 12;
	{8'd58,8'd203} : s = 81;
	{8'd58,8'd204} : s = 76;
	{8'd58,8'd205} : s = 195;
	{8'd58,8'd206} : s = 10;
	{8'd58,8'd207} : s = 74;
	{8'd58,8'd208} : s = 73;
	{8'd58,8'd209} : s = 184;
	{8'd58,8'd210} : s = 70;
	{8'd58,8'd211} : s = 180;
	{8'd58,8'd212} : s = 178;
	{8'd58,8'd213} : s = 314;
	{8'd58,8'd214} : s = 9;
	{8'd58,8'd215} : s = 69;
	{8'd58,8'd216} : s = 67;
	{8'd58,8'd217} : s = 177;
	{8'd58,8'd218} : s = 56;
	{8'd58,8'd219} : s = 172;
	{8'd58,8'd220} : s = 170;
	{8'd58,8'd221} : s = 313;
	{8'd58,8'd222} : s = 52;
	{8'd58,8'd223} : s = 169;
	{8'd58,8'd224} : s = 166;
	{8'd58,8'd225} : s = 310;
	{8'd58,8'd226} : s = 165;
	{8'd58,8'd227} : s = 309;
	{8'd58,8'd228} : s = 307;
	{8'd58,8'd229} : s = 427;
	{8'd58,8'd230} : s = 6;
	{8'd58,8'd231} : s = 50;
	{8'd58,8'd232} : s = 49;
	{8'd58,8'd233} : s = 163;
	{8'd58,8'd234} : s = 44;
	{8'd58,8'd235} : s = 156;
	{8'd58,8'd236} : s = 154;
	{8'd58,8'd237} : s = 302;
	{8'd58,8'd238} : s = 42;
	{8'd58,8'd239} : s = 153;
	{8'd58,8'd240} : s = 150;
	{8'd58,8'd241} : s = 301;
	{8'd58,8'd242} : s = 149;
	{8'd58,8'd243} : s = 299;
	{8'd58,8'd244} : s = 295;
	{8'd58,8'd245} : s = 423;
	{8'd58,8'd246} : s = 41;
	{8'd58,8'd247} : s = 147;
	{8'd58,8'd248} : s = 142;
	{8'd58,8'd249} : s = 286;
	{8'd58,8'd250} : s = 141;
	{8'd58,8'd251} : s = 285;
	{8'd58,8'd252} : s = 283;
	{8'd58,8'd253} : s = 414;
	{8'd58,8'd254} : s = 139;
	{8'd58,8'd255} : s = 279;
	{8'd59,8'd0} : s = 482;
	{8'd59,8'd1} : s = 401;
	{8'd59,8'd2} : s = 481;
	{8'd59,8'd3} : s = 472;
	{8'd59,8'd4} : s = 504;
	{8'd59,8'd5} : s = 4;
	{8'd59,8'd6} : s = 96;
	{8'd59,8'd7} : s = 80;
	{8'd59,8'd8} : s = 274;
	{8'd59,8'd9} : s = 72;
	{8'd59,8'd10} : s = 273;
	{8'd59,8'd11} : s = 268;
	{8'd59,8'd12} : s = 396;
	{8'd59,8'd13} : s = 68;
	{8'd59,8'd14} : s = 266;
	{8'd59,8'd15} : s = 265;
	{8'd59,8'd16} : s = 394;
	{8'd59,8'd17} : s = 262;
	{8'd59,8'd18} : s = 393;
	{8'd59,8'd19} : s = 390;
	{8'd59,8'd20} : s = 468;
	{8'd59,8'd21} : s = 66;
	{8'd59,8'd22} : s = 261;
	{8'd59,8'd23} : s = 259;
	{8'd59,8'd24} : s = 389;
	{8'd59,8'd25} : s = 224;
	{8'd59,8'd26} : s = 387;
	{8'd59,8'd27} : s = 368;
	{8'd59,8'd28} : s = 466;
	{8'd59,8'd29} : s = 208;
	{8'd59,8'd30} : s = 360;
	{8'd59,8'd31} : s = 356;
	{8'd59,8'd32} : s = 465;
	{8'd59,8'd33} : s = 354;
	{8'd59,8'd34} : s = 460;
	{8'd59,8'd35} : s = 458;
	{8'd59,8'd36} : s = 500;
	{8'd59,8'd37} : s = 65;
	{8'd59,8'd38} : s = 200;
	{8'd59,8'd39} : s = 196;
	{8'd59,8'd40} : s = 353;
	{8'd59,8'd41} : s = 194;
	{8'd59,8'd42} : s = 344;
	{8'd59,8'd43} : s = 340;
	{8'd59,8'd44} : s = 457;
	{8'd59,8'd45} : s = 193;
	{8'd59,8'd46} : s = 338;
	{8'd59,8'd47} : s = 337;
	{8'd59,8'd48} : s = 454;
	{8'd59,8'd49} : s = 332;
	{8'd59,8'd50} : s = 453;
	{8'd59,8'd51} : s = 451;
	{8'd59,8'd52} : s = 498;
	{8'd59,8'd53} : s = 176;
	{8'd59,8'd54} : s = 330;
	{8'd59,8'd55} : s = 329;
	{8'd59,8'd56} : s = 440;
	{8'd59,8'd57} : s = 326;
	{8'd59,8'd58} : s = 436;
	{8'd59,8'd59} : s = 434;
	{8'd59,8'd60} : s = 497;
	{8'd59,8'd61} : s = 325;
	{8'd59,8'd62} : s = 433;
	{8'd59,8'd63} : s = 428;
	{8'd59,8'd64} : s = 492;
	{8'd59,8'd65} : s = 426;
	{8'd59,8'd66} : s = 490;
	{8'd59,8'd67} : s = 489;
	{8'd59,8'd68} : s = 508;
	{8'd59,8'd69} : s = 2;
	{8'd59,8'd70} : s = 48;
	{8'd59,8'd71} : s = 40;
	{8'd59,8'd72} : s = 168;
	{8'd59,8'd73} : s = 36;
	{8'd59,8'd74} : s = 164;
	{8'd59,8'd75} : s = 162;
	{8'd59,8'd76} : s = 323;
	{8'd59,8'd77} : s = 34;
	{8'd59,8'd78} : s = 161;
	{8'd59,8'd79} : s = 152;
	{8'd59,8'd80} : s = 312;
	{8'd59,8'd81} : s = 148;
	{8'd59,8'd82} : s = 308;
	{8'd59,8'd83} : s = 306;
	{8'd59,8'd84} : s = 425;
	{8'd59,8'd85} : s = 33;
	{8'd59,8'd86} : s = 146;
	{8'd59,8'd87} : s = 145;
	{8'd59,8'd88} : s = 305;
	{8'd59,8'd89} : s = 140;
	{8'd59,8'd90} : s = 300;
	{8'd59,8'd91} : s = 298;
	{8'd59,8'd92} : s = 422;
	{8'd59,8'd93} : s = 138;
	{8'd59,8'd94} : s = 297;
	{8'd59,8'd95} : s = 294;
	{8'd59,8'd96} : s = 421;
	{8'd59,8'd97} : s = 293;
	{8'd59,8'd98} : s = 419;
	{8'd59,8'd99} : s = 412;
	{8'd59,8'd100} : s = 486;
	{8'd59,8'd101} : s = 24;
	{8'd59,8'd102} : s = 137;
	{8'd59,8'd103} : s = 134;
	{8'd59,8'd104} : s = 291;
	{8'd59,8'd105} : s = 133;
	{8'd59,8'd106} : s = 284;
	{8'd59,8'd107} : s = 282;
	{8'd59,8'd108} : s = 410;
	{8'd59,8'd109} : s = 131;
	{8'd59,8'd110} : s = 281;
	{8'd59,8'd111} : s = 278;
	{8'd59,8'd112} : s = 409;
	{8'd59,8'd113} : s = 277;
	{8'd59,8'd114} : s = 406;
	{8'd59,8'd115} : s = 405;
	{8'd59,8'd116} : s = 485;
	{8'd59,8'd117} : s = 112;
	{8'd59,8'd118} : s = 275;
	{8'd59,8'd119} : s = 270;
	{8'd59,8'd120} : s = 403;
	{8'd59,8'd121} : s = 269;
	{8'd59,8'd122} : s = 398;
	{8'd59,8'd123} : s = 397;
	{8'd59,8'd124} : s = 483;
	{8'd59,8'd125} : s = 267;
	{8'd59,8'd126} : s = 395;
	{8'd59,8'd127} : s = 391;
	{8'd59,8'd128} : s = 476;
	{8'd59,8'd129} : s = 376;
	{8'd59,8'd130} : s = 474;
	{8'd59,8'd131} : s = 473;
	{8'd59,8'd132} : s = 506;
	{8'd59,8'd133} : s = 20;
	{8'd59,8'd134} : s = 104;
	{8'd59,8'd135} : s = 100;
	{8'd59,8'd136} : s = 263;
	{8'd59,8'd137} : s = 98;
	{8'd59,8'd138} : s = 240;
	{8'd59,8'd139} : s = 232;
	{8'd59,8'd140} : s = 372;
	{8'd59,8'd141} : s = 97;
	{8'd59,8'd142} : s = 228;
	{8'd59,8'd143} : s = 226;
	{8'd59,8'd144} : s = 370;
	{8'd59,8'd145} : s = 225;
	{8'd59,8'd146} : s = 369;
	{8'd59,8'd147} : s = 364;
	{8'd59,8'd148} : s = 470;
	{8'd59,8'd149} : s = 88;
	{8'd59,8'd150} : s = 216;
	{8'd59,8'd151} : s = 212;
	{8'd59,8'd152} : s = 362;
	{8'd59,8'd153} : s = 210;
	{8'd59,8'd154} : s = 361;
	{8'd59,8'd155} : s = 358;
	{8'd59,8'd156} : s = 469;
	{8'd59,8'd157} : s = 209;
	{8'd59,8'd158} : s = 357;
	{8'd59,8'd159} : s = 355;
	{8'd59,8'd160} : s = 467;
	{8'd59,8'd161} : s = 348;
	{8'd59,8'd162} : s = 462;
	{8'd59,8'd163} : s = 461;
	{8'd59,8'd164} : s = 505;
	{8'd59,8'd165} : s = 84;
	{8'd59,8'd166} : s = 204;
	{8'd59,8'd167} : s = 202;
	{8'd59,8'd168} : s = 346;
	{8'd59,8'd169} : s = 201;
	{8'd59,8'd170} : s = 345;
	{8'd59,8'd171} : s = 342;
	{8'd59,8'd172} : s = 459;
	{8'd59,8'd173} : s = 198;
	{8'd59,8'd174} : s = 341;
	{8'd59,8'd175} : s = 339;
	{8'd59,8'd176} : s = 455;
	{8'd59,8'd177} : s = 334;
	{8'd59,8'd178} : s = 444;
	{8'd59,8'd179} : s = 442;
	{8'd59,8'd180} : s = 502;
	{8'd59,8'd181} : s = 197;
	{8'd59,8'd182} : s = 333;
	{8'd59,8'd183} : s = 331;
	{8'd59,8'd184} : s = 441;
	{8'd59,8'd185} : s = 327;
	{8'd59,8'd186} : s = 438;
	{8'd59,8'd187} : s = 437;
	{8'd59,8'd188} : s = 501;
	{8'd59,8'd189} : s = 316;
	{8'd59,8'd190} : s = 435;
	{8'd59,8'd191} : s = 430;
	{8'd59,8'd192} : s = 499;
	{8'd59,8'd193} : s = 429;
	{8'd59,8'd194} : s = 494;
	{8'd59,8'd195} : s = 493;
	{8'd59,8'd196} : s = 510;
	{8'd59,8'd197} : s = 1;
	{8'd59,8'd198} : s = 18;
	{8'd59,8'd199} : s = 17;
	{8'd59,8'd200} : s = 82;
	{8'd59,8'd201} : s = 12;
	{8'd59,8'd202} : s = 81;
	{8'd59,8'd203} : s = 76;
	{8'd59,8'd204} : s = 195;
	{8'd59,8'd205} : s = 10;
	{8'd59,8'd206} : s = 74;
	{8'd59,8'd207} : s = 73;
	{8'd59,8'd208} : s = 184;
	{8'd59,8'd209} : s = 70;
	{8'd59,8'd210} : s = 180;
	{8'd59,8'd211} : s = 178;
	{8'd59,8'd212} : s = 314;
	{8'd59,8'd213} : s = 9;
	{8'd59,8'd214} : s = 69;
	{8'd59,8'd215} : s = 67;
	{8'd59,8'd216} : s = 177;
	{8'd59,8'd217} : s = 56;
	{8'd59,8'd218} : s = 172;
	{8'd59,8'd219} : s = 170;
	{8'd59,8'd220} : s = 313;
	{8'd59,8'd221} : s = 52;
	{8'd59,8'd222} : s = 169;
	{8'd59,8'd223} : s = 166;
	{8'd59,8'd224} : s = 310;
	{8'd59,8'd225} : s = 165;
	{8'd59,8'd226} : s = 309;
	{8'd59,8'd227} : s = 307;
	{8'd59,8'd228} : s = 427;
	{8'd59,8'd229} : s = 6;
	{8'd59,8'd230} : s = 50;
	{8'd59,8'd231} : s = 49;
	{8'd59,8'd232} : s = 163;
	{8'd59,8'd233} : s = 44;
	{8'd59,8'd234} : s = 156;
	{8'd59,8'd235} : s = 154;
	{8'd59,8'd236} : s = 302;
	{8'd59,8'd237} : s = 42;
	{8'd59,8'd238} : s = 153;
	{8'd59,8'd239} : s = 150;
	{8'd59,8'd240} : s = 301;
	{8'd59,8'd241} : s = 149;
	{8'd59,8'd242} : s = 299;
	{8'd59,8'd243} : s = 295;
	{8'd59,8'd244} : s = 423;
	{8'd59,8'd245} : s = 41;
	{8'd59,8'd246} : s = 147;
	{8'd59,8'd247} : s = 142;
	{8'd59,8'd248} : s = 286;
	{8'd59,8'd249} : s = 141;
	{8'd59,8'd250} : s = 285;
	{8'd59,8'd251} : s = 283;
	{8'd59,8'd252} : s = 414;
	{8'd59,8'd253} : s = 139;
	{8'd59,8'd254} : s = 279;
	{8'd59,8'd255} : s = 271;
	{8'd60,8'd0} : s = 401;
	{8'd60,8'd1} : s = 481;
	{8'd60,8'd2} : s = 472;
	{8'd60,8'd3} : s = 504;
	{8'd60,8'd4} : s = 4;
	{8'd60,8'd5} : s = 96;
	{8'd60,8'd6} : s = 80;
	{8'd60,8'd7} : s = 274;
	{8'd60,8'd8} : s = 72;
	{8'd60,8'd9} : s = 273;
	{8'd60,8'd10} : s = 268;
	{8'd60,8'd11} : s = 396;
	{8'd60,8'd12} : s = 68;
	{8'd60,8'd13} : s = 266;
	{8'd60,8'd14} : s = 265;
	{8'd60,8'd15} : s = 394;
	{8'd60,8'd16} : s = 262;
	{8'd60,8'd17} : s = 393;
	{8'd60,8'd18} : s = 390;
	{8'd60,8'd19} : s = 468;
	{8'd60,8'd20} : s = 66;
	{8'd60,8'd21} : s = 261;
	{8'd60,8'd22} : s = 259;
	{8'd60,8'd23} : s = 389;
	{8'd60,8'd24} : s = 224;
	{8'd60,8'd25} : s = 387;
	{8'd60,8'd26} : s = 368;
	{8'd60,8'd27} : s = 466;
	{8'd60,8'd28} : s = 208;
	{8'd60,8'd29} : s = 360;
	{8'd60,8'd30} : s = 356;
	{8'd60,8'd31} : s = 465;
	{8'd60,8'd32} : s = 354;
	{8'd60,8'd33} : s = 460;
	{8'd60,8'd34} : s = 458;
	{8'd60,8'd35} : s = 500;
	{8'd60,8'd36} : s = 65;
	{8'd60,8'd37} : s = 200;
	{8'd60,8'd38} : s = 196;
	{8'd60,8'd39} : s = 353;
	{8'd60,8'd40} : s = 194;
	{8'd60,8'd41} : s = 344;
	{8'd60,8'd42} : s = 340;
	{8'd60,8'd43} : s = 457;
	{8'd60,8'd44} : s = 193;
	{8'd60,8'd45} : s = 338;
	{8'd60,8'd46} : s = 337;
	{8'd60,8'd47} : s = 454;
	{8'd60,8'd48} : s = 332;
	{8'd60,8'd49} : s = 453;
	{8'd60,8'd50} : s = 451;
	{8'd60,8'd51} : s = 498;
	{8'd60,8'd52} : s = 176;
	{8'd60,8'd53} : s = 330;
	{8'd60,8'd54} : s = 329;
	{8'd60,8'd55} : s = 440;
	{8'd60,8'd56} : s = 326;
	{8'd60,8'd57} : s = 436;
	{8'd60,8'd58} : s = 434;
	{8'd60,8'd59} : s = 497;
	{8'd60,8'd60} : s = 325;
	{8'd60,8'd61} : s = 433;
	{8'd60,8'd62} : s = 428;
	{8'd60,8'd63} : s = 492;
	{8'd60,8'd64} : s = 426;
	{8'd60,8'd65} : s = 490;
	{8'd60,8'd66} : s = 489;
	{8'd60,8'd67} : s = 508;
	{8'd60,8'd68} : s = 2;
	{8'd60,8'd69} : s = 48;
	{8'd60,8'd70} : s = 40;
	{8'd60,8'd71} : s = 168;
	{8'd60,8'd72} : s = 36;
	{8'd60,8'd73} : s = 164;
	{8'd60,8'd74} : s = 162;
	{8'd60,8'd75} : s = 323;
	{8'd60,8'd76} : s = 34;
	{8'd60,8'd77} : s = 161;
	{8'd60,8'd78} : s = 152;
	{8'd60,8'd79} : s = 312;
	{8'd60,8'd80} : s = 148;
	{8'd60,8'd81} : s = 308;
	{8'd60,8'd82} : s = 306;
	{8'd60,8'd83} : s = 425;
	{8'd60,8'd84} : s = 33;
	{8'd60,8'd85} : s = 146;
	{8'd60,8'd86} : s = 145;
	{8'd60,8'd87} : s = 305;
	{8'd60,8'd88} : s = 140;
	{8'd60,8'd89} : s = 300;
	{8'd60,8'd90} : s = 298;
	{8'd60,8'd91} : s = 422;
	{8'd60,8'd92} : s = 138;
	{8'd60,8'd93} : s = 297;
	{8'd60,8'd94} : s = 294;
	{8'd60,8'd95} : s = 421;
	{8'd60,8'd96} : s = 293;
	{8'd60,8'd97} : s = 419;
	{8'd60,8'd98} : s = 412;
	{8'd60,8'd99} : s = 486;
	{8'd60,8'd100} : s = 24;
	{8'd60,8'd101} : s = 137;
	{8'd60,8'd102} : s = 134;
	{8'd60,8'd103} : s = 291;
	{8'd60,8'd104} : s = 133;
	{8'd60,8'd105} : s = 284;
	{8'd60,8'd106} : s = 282;
	{8'd60,8'd107} : s = 410;
	{8'd60,8'd108} : s = 131;
	{8'd60,8'd109} : s = 281;
	{8'd60,8'd110} : s = 278;
	{8'd60,8'd111} : s = 409;
	{8'd60,8'd112} : s = 277;
	{8'd60,8'd113} : s = 406;
	{8'd60,8'd114} : s = 405;
	{8'd60,8'd115} : s = 485;
	{8'd60,8'd116} : s = 112;
	{8'd60,8'd117} : s = 275;
	{8'd60,8'd118} : s = 270;
	{8'd60,8'd119} : s = 403;
	{8'd60,8'd120} : s = 269;
	{8'd60,8'd121} : s = 398;
	{8'd60,8'd122} : s = 397;
	{8'd60,8'd123} : s = 483;
	{8'd60,8'd124} : s = 267;
	{8'd60,8'd125} : s = 395;
	{8'd60,8'd126} : s = 391;
	{8'd60,8'd127} : s = 476;
	{8'd60,8'd128} : s = 376;
	{8'd60,8'd129} : s = 474;
	{8'd60,8'd130} : s = 473;
	{8'd60,8'd131} : s = 506;
	{8'd60,8'd132} : s = 20;
	{8'd60,8'd133} : s = 104;
	{8'd60,8'd134} : s = 100;
	{8'd60,8'd135} : s = 263;
	{8'd60,8'd136} : s = 98;
	{8'd60,8'd137} : s = 240;
	{8'd60,8'd138} : s = 232;
	{8'd60,8'd139} : s = 372;
	{8'd60,8'd140} : s = 97;
	{8'd60,8'd141} : s = 228;
	{8'd60,8'd142} : s = 226;
	{8'd60,8'd143} : s = 370;
	{8'd60,8'd144} : s = 225;
	{8'd60,8'd145} : s = 369;
	{8'd60,8'd146} : s = 364;
	{8'd60,8'd147} : s = 470;
	{8'd60,8'd148} : s = 88;
	{8'd60,8'd149} : s = 216;
	{8'd60,8'd150} : s = 212;
	{8'd60,8'd151} : s = 362;
	{8'd60,8'd152} : s = 210;
	{8'd60,8'd153} : s = 361;
	{8'd60,8'd154} : s = 358;
	{8'd60,8'd155} : s = 469;
	{8'd60,8'd156} : s = 209;
	{8'd60,8'd157} : s = 357;
	{8'd60,8'd158} : s = 355;
	{8'd60,8'd159} : s = 467;
	{8'd60,8'd160} : s = 348;
	{8'd60,8'd161} : s = 462;
	{8'd60,8'd162} : s = 461;
	{8'd60,8'd163} : s = 505;
	{8'd60,8'd164} : s = 84;
	{8'd60,8'd165} : s = 204;
	{8'd60,8'd166} : s = 202;
	{8'd60,8'd167} : s = 346;
	{8'd60,8'd168} : s = 201;
	{8'd60,8'd169} : s = 345;
	{8'd60,8'd170} : s = 342;
	{8'd60,8'd171} : s = 459;
	{8'd60,8'd172} : s = 198;
	{8'd60,8'd173} : s = 341;
	{8'd60,8'd174} : s = 339;
	{8'd60,8'd175} : s = 455;
	{8'd60,8'd176} : s = 334;
	{8'd60,8'd177} : s = 444;
	{8'd60,8'd178} : s = 442;
	{8'd60,8'd179} : s = 502;
	{8'd60,8'd180} : s = 197;
	{8'd60,8'd181} : s = 333;
	{8'd60,8'd182} : s = 331;
	{8'd60,8'd183} : s = 441;
	{8'd60,8'd184} : s = 327;
	{8'd60,8'd185} : s = 438;
	{8'd60,8'd186} : s = 437;
	{8'd60,8'd187} : s = 501;
	{8'd60,8'd188} : s = 316;
	{8'd60,8'd189} : s = 435;
	{8'd60,8'd190} : s = 430;
	{8'd60,8'd191} : s = 499;
	{8'd60,8'd192} : s = 429;
	{8'd60,8'd193} : s = 494;
	{8'd60,8'd194} : s = 493;
	{8'd60,8'd195} : s = 510;
	{8'd60,8'd196} : s = 1;
	{8'd60,8'd197} : s = 18;
	{8'd60,8'd198} : s = 17;
	{8'd60,8'd199} : s = 82;
	{8'd60,8'd200} : s = 12;
	{8'd60,8'd201} : s = 81;
	{8'd60,8'd202} : s = 76;
	{8'd60,8'd203} : s = 195;
	{8'd60,8'd204} : s = 10;
	{8'd60,8'd205} : s = 74;
	{8'd60,8'd206} : s = 73;
	{8'd60,8'd207} : s = 184;
	{8'd60,8'd208} : s = 70;
	{8'd60,8'd209} : s = 180;
	{8'd60,8'd210} : s = 178;
	{8'd60,8'd211} : s = 314;
	{8'd60,8'd212} : s = 9;
	{8'd60,8'd213} : s = 69;
	{8'd60,8'd214} : s = 67;
	{8'd60,8'd215} : s = 177;
	{8'd60,8'd216} : s = 56;
	{8'd60,8'd217} : s = 172;
	{8'd60,8'd218} : s = 170;
	{8'd60,8'd219} : s = 313;
	{8'd60,8'd220} : s = 52;
	{8'd60,8'd221} : s = 169;
	{8'd60,8'd222} : s = 166;
	{8'd60,8'd223} : s = 310;
	{8'd60,8'd224} : s = 165;
	{8'd60,8'd225} : s = 309;
	{8'd60,8'd226} : s = 307;
	{8'd60,8'd227} : s = 427;
	{8'd60,8'd228} : s = 6;
	{8'd60,8'd229} : s = 50;
	{8'd60,8'd230} : s = 49;
	{8'd60,8'd231} : s = 163;
	{8'd60,8'd232} : s = 44;
	{8'd60,8'd233} : s = 156;
	{8'd60,8'd234} : s = 154;
	{8'd60,8'd235} : s = 302;
	{8'd60,8'd236} : s = 42;
	{8'd60,8'd237} : s = 153;
	{8'd60,8'd238} : s = 150;
	{8'd60,8'd239} : s = 301;
	{8'd60,8'd240} : s = 149;
	{8'd60,8'd241} : s = 299;
	{8'd60,8'd242} : s = 295;
	{8'd60,8'd243} : s = 423;
	{8'd60,8'd244} : s = 41;
	{8'd60,8'd245} : s = 147;
	{8'd60,8'd246} : s = 142;
	{8'd60,8'd247} : s = 286;
	{8'd60,8'd248} : s = 141;
	{8'd60,8'd249} : s = 285;
	{8'd60,8'd250} : s = 283;
	{8'd60,8'd251} : s = 414;
	{8'd60,8'd252} : s = 139;
	{8'd60,8'd253} : s = 279;
	{8'd60,8'd254} : s = 271;
	{8'd60,8'd255} : s = 413;
	{8'd61,8'd0} : s = 481;
	{8'd61,8'd1} : s = 472;
	{8'd61,8'd2} : s = 504;
	{8'd61,8'd3} : s = 4;
	{8'd61,8'd4} : s = 96;
	{8'd61,8'd5} : s = 80;
	{8'd61,8'd6} : s = 274;
	{8'd61,8'd7} : s = 72;
	{8'd61,8'd8} : s = 273;
	{8'd61,8'd9} : s = 268;
	{8'd61,8'd10} : s = 396;
	{8'd61,8'd11} : s = 68;
	{8'd61,8'd12} : s = 266;
	{8'd61,8'd13} : s = 265;
	{8'd61,8'd14} : s = 394;
	{8'd61,8'd15} : s = 262;
	{8'd61,8'd16} : s = 393;
	{8'd61,8'd17} : s = 390;
	{8'd61,8'd18} : s = 468;
	{8'd61,8'd19} : s = 66;
	{8'd61,8'd20} : s = 261;
	{8'd61,8'd21} : s = 259;
	{8'd61,8'd22} : s = 389;
	{8'd61,8'd23} : s = 224;
	{8'd61,8'd24} : s = 387;
	{8'd61,8'd25} : s = 368;
	{8'd61,8'd26} : s = 466;
	{8'd61,8'd27} : s = 208;
	{8'd61,8'd28} : s = 360;
	{8'd61,8'd29} : s = 356;
	{8'd61,8'd30} : s = 465;
	{8'd61,8'd31} : s = 354;
	{8'd61,8'd32} : s = 460;
	{8'd61,8'd33} : s = 458;
	{8'd61,8'd34} : s = 500;
	{8'd61,8'd35} : s = 65;
	{8'd61,8'd36} : s = 200;
	{8'd61,8'd37} : s = 196;
	{8'd61,8'd38} : s = 353;
	{8'd61,8'd39} : s = 194;
	{8'd61,8'd40} : s = 344;
	{8'd61,8'd41} : s = 340;
	{8'd61,8'd42} : s = 457;
	{8'd61,8'd43} : s = 193;
	{8'd61,8'd44} : s = 338;
	{8'd61,8'd45} : s = 337;
	{8'd61,8'd46} : s = 454;
	{8'd61,8'd47} : s = 332;
	{8'd61,8'd48} : s = 453;
	{8'd61,8'd49} : s = 451;
	{8'd61,8'd50} : s = 498;
	{8'd61,8'd51} : s = 176;
	{8'd61,8'd52} : s = 330;
	{8'd61,8'd53} : s = 329;
	{8'd61,8'd54} : s = 440;
	{8'd61,8'd55} : s = 326;
	{8'd61,8'd56} : s = 436;
	{8'd61,8'd57} : s = 434;
	{8'd61,8'd58} : s = 497;
	{8'd61,8'd59} : s = 325;
	{8'd61,8'd60} : s = 433;
	{8'd61,8'd61} : s = 428;
	{8'd61,8'd62} : s = 492;
	{8'd61,8'd63} : s = 426;
	{8'd61,8'd64} : s = 490;
	{8'd61,8'd65} : s = 489;
	{8'd61,8'd66} : s = 508;
	{8'd61,8'd67} : s = 2;
	{8'd61,8'd68} : s = 48;
	{8'd61,8'd69} : s = 40;
	{8'd61,8'd70} : s = 168;
	{8'd61,8'd71} : s = 36;
	{8'd61,8'd72} : s = 164;
	{8'd61,8'd73} : s = 162;
	{8'd61,8'd74} : s = 323;
	{8'd61,8'd75} : s = 34;
	{8'd61,8'd76} : s = 161;
	{8'd61,8'd77} : s = 152;
	{8'd61,8'd78} : s = 312;
	{8'd61,8'd79} : s = 148;
	{8'd61,8'd80} : s = 308;
	{8'd61,8'd81} : s = 306;
	{8'd61,8'd82} : s = 425;
	{8'd61,8'd83} : s = 33;
	{8'd61,8'd84} : s = 146;
	{8'd61,8'd85} : s = 145;
	{8'd61,8'd86} : s = 305;
	{8'd61,8'd87} : s = 140;
	{8'd61,8'd88} : s = 300;
	{8'd61,8'd89} : s = 298;
	{8'd61,8'd90} : s = 422;
	{8'd61,8'd91} : s = 138;
	{8'd61,8'd92} : s = 297;
	{8'd61,8'd93} : s = 294;
	{8'd61,8'd94} : s = 421;
	{8'd61,8'd95} : s = 293;
	{8'd61,8'd96} : s = 419;
	{8'd61,8'd97} : s = 412;
	{8'd61,8'd98} : s = 486;
	{8'd61,8'd99} : s = 24;
	{8'd61,8'd100} : s = 137;
	{8'd61,8'd101} : s = 134;
	{8'd61,8'd102} : s = 291;
	{8'd61,8'd103} : s = 133;
	{8'd61,8'd104} : s = 284;
	{8'd61,8'd105} : s = 282;
	{8'd61,8'd106} : s = 410;
	{8'd61,8'd107} : s = 131;
	{8'd61,8'd108} : s = 281;
	{8'd61,8'd109} : s = 278;
	{8'd61,8'd110} : s = 409;
	{8'd61,8'd111} : s = 277;
	{8'd61,8'd112} : s = 406;
	{8'd61,8'd113} : s = 405;
	{8'd61,8'd114} : s = 485;
	{8'd61,8'd115} : s = 112;
	{8'd61,8'd116} : s = 275;
	{8'd61,8'd117} : s = 270;
	{8'd61,8'd118} : s = 403;
	{8'd61,8'd119} : s = 269;
	{8'd61,8'd120} : s = 398;
	{8'd61,8'd121} : s = 397;
	{8'd61,8'd122} : s = 483;
	{8'd61,8'd123} : s = 267;
	{8'd61,8'd124} : s = 395;
	{8'd61,8'd125} : s = 391;
	{8'd61,8'd126} : s = 476;
	{8'd61,8'd127} : s = 376;
	{8'd61,8'd128} : s = 474;
	{8'd61,8'd129} : s = 473;
	{8'd61,8'd130} : s = 506;
	{8'd61,8'd131} : s = 20;
	{8'd61,8'd132} : s = 104;
	{8'd61,8'd133} : s = 100;
	{8'd61,8'd134} : s = 263;
	{8'd61,8'd135} : s = 98;
	{8'd61,8'd136} : s = 240;
	{8'd61,8'd137} : s = 232;
	{8'd61,8'd138} : s = 372;
	{8'd61,8'd139} : s = 97;
	{8'd61,8'd140} : s = 228;
	{8'd61,8'd141} : s = 226;
	{8'd61,8'd142} : s = 370;
	{8'd61,8'd143} : s = 225;
	{8'd61,8'd144} : s = 369;
	{8'd61,8'd145} : s = 364;
	{8'd61,8'd146} : s = 470;
	{8'd61,8'd147} : s = 88;
	{8'd61,8'd148} : s = 216;
	{8'd61,8'd149} : s = 212;
	{8'd61,8'd150} : s = 362;
	{8'd61,8'd151} : s = 210;
	{8'd61,8'd152} : s = 361;
	{8'd61,8'd153} : s = 358;
	{8'd61,8'd154} : s = 469;
	{8'd61,8'd155} : s = 209;
	{8'd61,8'd156} : s = 357;
	{8'd61,8'd157} : s = 355;
	{8'd61,8'd158} : s = 467;
	{8'd61,8'd159} : s = 348;
	{8'd61,8'd160} : s = 462;
	{8'd61,8'd161} : s = 461;
	{8'd61,8'd162} : s = 505;
	{8'd61,8'd163} : s = 84;
	{8'd61,8'd164} : s = 204;
	{8'd61,8'd165} : s = 202;
	{8'd61,8'd166} : s = 346;
	{8'd61,8'd167} : s = 201;
	{8'd61,8'd168} : s = 345;
	{8'd61,8'd169} : s = 342;
	{8'd61,8'd170} : s = 459;
	{8'd61,8'd171} : s = 198;
	{8'd61,8'd172} : s = 341;
	{8'd61,8'd173} : s = 339;
	{8'd61,8'd174} : s = 455;
	{8'd61,8'd175} : s = 334;
	{8'd61,8'd176} : s = 444;
	{8'd61,8'd177} : s = 442;
	{8'd61,8'd178} : s = 502;
	{8'd61,8'd179} : s = 197;
	{8'd61,8'd180} : s = 333;
	{8'd61,8'd181} : s = 331;
	{8'd61,8'd182} : s = 441;
	{8'd61,8'd183} : s = 327;
	{8'd61,8'd184} : s = 438;
	{8'd61,8'd185} : s = 437;
	{8'd61,8'd186} : s = 501;
	{8'd61,8'd187} : s = 316;
	{8'd61,8'd188} : s = 435;
	{8'd61,8'd189} : s = 430;
	{8'd61,8'd190} : s = 499;
	{8'd61,8'd191} : s = 429;
	{8'd61,8'd192} : s = 494;
	{8'd61,8'd193} : s = 493;
	{8'd61,8'd194} : s = 510;
	{8'd61,8'd195} : s = 1;
	{8'd61,8'd196} : s = 18;
	{8'd61,8'd197} : s = 17;
	{8'd61,8'd198} : s = 82;
	{8'd61,8'd199} : s = 12;
	{8'd61,8'd200} : s = 81;
	{8'd61,8'd201} : s = 76;
	{8'd61,8'd202} : s = 195;
	{8'd61,8'd203} : s = 10;
	{8'd61,8'd204} : s = 74;
	{8'd61,8'd205} : s = 73;
	{8'd61,8'd206} : s = 184;
	{8'd61,8'd207} : s = 70;
	{8'd61,8'd208} : s = 180;
	{8'd61,8'd209} : s = 178;
	{8'd61,8'd210} : s = 314;
	{8'd61,8'd211} : s = 9;
	{8'd61,8'd212} : s = 69;
	{8'd61,8'd213} : s = 67;
	{8'd61,8'd214} : s = 177;
	{8'd61,8'd215} : s = 56;
	{8'd61,8'd216} : s = 172;
	{8'd61,8'd217} : s = 170;
	{8'd61,8'd218} : s = 313;
	{8'd61,8'd219} : s = 52;
	{8'd61,8'd220} : s = 169;
	{8'd61,8'd221} : s = 166;
	{8'd61,8'd222} : s = 310;
	{8'd61,8'd223} : s = 165;
	{8'd61,8'd224} : s = 309;
	{8'd61,8'd225} : s = 307;
	{8'd61,8'd226} : s = 427;
	{8'd61,8'd227} : s = 6;
	{8'd61,8'd228} : s = 50;
	{8'd61,8'd229} : s = 49;
	{8'd61,8'd230} : s = 163;
	{8'd61,8'd231} : s = 44;
	{8'd61,8'd232} : s = 156;
	{8'd61,8'd233} : s = 154;
	{8'd61,8'd234} : s = 302;
	{8'd61,8'd235} : s = 42;
	{8'd61,8'd236} : s = 153;
	{8'd61,8'd237} : s = 150;
	{8'd61,8'd238} : s = 301;
	{8'd61,8'd239} : s = 149;
	{8'd61,8'd240} : s = 299;
	{8'd61,8'd241} : s = 295;
	{8'd61,8'd242} : s = 423;
	{8'd61,8'd243} : s = 41;
	{8'd61,8'd244} : s = 147;
	{8'd61,8'd245} : s = 142;
	{8'd61,8'd246} : s = 286;
	{8'd61,8'd247} : s = 141;
	{8'd61,8'd248} : s = 285;
	{8'd61,8'd249} : s = 283;
	{8'd61,8'd250} : s = 414;
	{8'd61,8'd251} : s = 139;
	{8'd61,8'd252} : s = 279;
	{8'd61,8'd253} : s = 271;
	{8'd61,8'd254} : s = 413;
	{8'd61,8'd255} : s = 248;
	{8'd62,8'd0} : s = 472;
	{8'd62,8'd1} : s = 504;
	{8'd62,8'd2} : s = 4;
	{8'd62,8'd3} : s = 96;
	{8'd62,8'd4} : s = 80;
	{8'd62,8'd5} : s = 274;
	{8'd62,8'd6} : s = 72;
	{8'd62,8'd7} : s = 273;
	{8'd62,8'd8} : s = 268;
	{8'd62,8'd9} : s = 396;
	{8'd62,8'd10} : s = 68;
	{8'd62,8'd11} : s = 266;
	{8'd62,8'd12} : s = 265;
	{8'd62,8'd13} : s = 394;
	{8'd62,8'd14} : s = 262;
	{8'd62,8'd15} : s = 393;
	{8'd62,8'd16} : s = 390;
	{8'd62,8'd17} : s = 468;
	{8'd62,8'd18} : s = 66;
	{8'd62,8'd19} : s = 261;
	{8'd62,8'd20} : s = 259;
	{8'd62,8'd21} : s = 389;
	{8'd62,8'd22} : s = 224;
	{8'd62,8'd23} : s = 387;
	{8'd62,8'd24} : s = 368;
	{8'd62,8'd25} : s = 466;
	{8'd62,8'd26} : s = 208;
	{8'd62,8'd27} : s = 360;
	{8'd62,8'd28} : s = 356;
	{8'd62,8'd29} : s = 465;
	{8'd62,8'd30} : s = 354;
	{8'd62,8'd31} : s = 460;
	{8'd62,8'd32} : s = 458;
	{8'd62,8'd33} : s = 500;
	{8'd62,8'd34} : s = 65;
	{8'd62,8'd35} : s = 200;
	{8'd62,8'd36} : s = 196;
	{8'd62,8'd37} : s = 353;
	{8'd62,8'd38} : s = 194;
	{8'd62,8'd39} : s = 344;
	{8'd62,8'd40} : s = 340;
	{8'd62,8'd41} : s = 457;
	{8'd62,8'd42} : s = 193;
	{8'd62,8'd43} : s = 338;
	{8'd62,8'd44} : s = 337;
	{8'd62,8'd45} : s = 454;
	{8'd62,8'd46} : s = 332;
	{8'd62,8'd47} : s = 453;
	{8'd62,8'd48} : s = 451;
	{8'd62,8'd49} : s = 498;
	{8'd62,8'd50} : s = 176;
	{8'd62,8'd51} : s = 330;
	{8'd62,8'd52} : s = 329;
	{8'd62,8'd53} : s = 440;
	{8'd62,8'd54} : s = 326;
	{8'd62,8'd55} : s = 436;
	{8'd62,8'd56} : s = 434;
	{8'd62,8'd57} : s = 497;
	{8'd62,8'd58} : s = 325;
	{8'd62,8'd59} : s = 433;
	{8'd62,8'd60} : s = 428;
	{8'd62,8'd61} : s = 492;
	{8'd62,8'd62} : s = 426;
	{8'd62,8'd63} : s = 490;
	{8'd62,8'd64} : s = 489;
	{8'd62,8'd65} : s = 508;
	{8'd62,8'd66} : s = 2;
	{8'd62,8'd67} : s = 48;
	{8'd62,8'd68} : s = 40;
	{8'd62,8'd69} : s = 168;
	{8'd62,8'd70} : s = 36;
	{8'd62,8'd71} : s = 164;
	{8'd62,8'd72} : s = 162;
	{8'd62,8'd73} : s = 323;
	{8'd62,8'd74} : s = 34;
	{8'd62,8'd75} : s = 161;
	{8'd62,8'd76} : s = 152;
	{8'd62,8'd77} : s = 312;
	{8'd62,8'd78} : s = 148;
	{8'd62,8'd79} : s = 308;
	{8'd62,8'd80} : s = 306;
	{8'd62,8'd81} : s = 425;
	{8'd62,8'd82} : s = 33;
	{8'd62,8'd83} : s = 146;
	{8'd62,8'd84} : s = 145;
	{8'd62,8'd85} : s = 305;
	{8'd62,8'd86} : s = 140;
	{8'd62,8'd87} : s = 300;
	{8'd62,8'd88} : s = 298;
	{8'd62,8'd89} : s = 422;
	{8'd62,8'd90} : s = 138;
	{8'd62,8'd91} : s = 297;
	{8'd62,8'd92} : s = 294;
	{8'd62,8'd93} : s = 421;
	{8'd62,8'd94} : s = 293;
	{8'd62,8'd95} : s = 419;
	{8'd62,8'd96} : s = 412;
	{8'd62,8'd97} : s = 486;
	{8'd62,8'd98} : s = 24;
	{8'd62,8'd99} : s = 137;
	{8'd62,8'd100} : s = 134;
	{8'd62,8'd101} : s = 291;
	{8'd62,8'd102} : s = 133;
	{8'd62,8'd103} : s = 284;
	{8'd62,8'd104} : s = 282;
	{8'd62,8'd105} : s = 410;
	{8'd62,8'd106} : s = 131;
	{8'd62,8'd107} : s = 281;
	{8'd62,8'd108} : s = 278;
	{8'd62,8'd109} : s = 409;
	{8'd62,8'd110} : s = 277;
	{8'd62,8'd111} : s = 406;
	{8'd62,8'd112} : s = 405;
	{8'd62,8'd113} : s = 485;
	{8'd62,8'd114} : s = 112;
	{8'd62,8'd115} : s = 275;
	{8'd62,8'd116} : s = 270;
	{8'd62,8'd117} : s = 403;
	{8'd62,8'd118} : s = 269;
	{8'd62,8'd119} : s = 398;
	{8'd62,8'd120} : s = 397;
	{8'd62,8'd121} : s = 483;
	{8'd62,8'd122} : s = 267;
	{8'd62,8'd123} : s = 395;
	{8'd62,8'd124} : s = 391;
	{8'd62,8'd125} : s = 476;
	{8'd62,8'd126} : s = 376;
	{8'd62,8'd127} : s = 474;
	{8'd62,8'd128} : s = 473;
	{8'd62,8'd129} : s = 506;
	{8'd62,8'd130} : s = 20;
	{8'd62,8'd131} : s = 104;
	{8'd62,8'd132} : s = 100;
	{8'd62,8'd133} : s = 263;
	{8'd62,8'd134} : s = 98;
	{8'd62,8'd135} : s = 240;
	{8'd62,8'd136} : s = 232;
	{8'd62,8'd137} : s = 372;
	{8'd62,8'd138} : s = 97;
	{8'd62,8'd139} : s = 228;
	{8'd62,8'd140} : s = 226;
	{8'd62,8'd141} : s = 370;
	{8'd62,8'd142} : s = 225;
	{8'd62,8'd143} : s = 369;
	{8'd62,8'd144} : s = 364;
	{8'd62,8'd145} : s = 470;
	{8'd62,8'd146} : s = 88;
	{8'd62,8'd147} : s = 216;
	{8'd62,8'd148} : s = 212;
	{8'd62,8'd149} : s = 362;
	{8'd62,8'd150} : s = 210;
	{8'd62,8'd151} : s = 361;
	{8'd62,8'd152} : s = 358;
	{8'd62,8'd153} : s = 469;
	{8'd62,8'd154} : s = 209;
	{8'd62,8'd155} : s = 357;
	{8'd62,8'd156} : s = 355;
	{8'd62,8'd157} : s = 467;
	{8'd62,8'd158} : s = 348;
	{8'd62,8'd159} : s = 462;
	{8'd62,8'd160} : s = 461;
	{8'd62,8'd161} : s = 505;
	{8'd62,8'd162} : s = 84;
	{8'd62,8'd163} : s = 204;
	{8'd62,8'd164} : s = 202;
	{8'd62,8'd165} : s = 346;
	{8'd62,8'd166} : s = 201;
	{8'd62,8'd167} : s = 345;
	{8'd62,8'd168} : s = 342;
	{8'd62,8'd169} : s = 459;
	{8'd62,8'd170} : s = 198;
	{8'd62,8'd171} : s = 341;
	{8'd62,8'd172} : s = 339;
	{8'd62,8'd173} : s = 455;
	{8'd62,8'd174} : s = 334;
	{8'd62,8'd175} : s = 444;
	{8'd62,8'd176} : s = 442;
	{8'd62,8'd177} : s = 502;
	{8'd62,8'd178} : s = 197;
	{8'd62,8'd179} : s = 333;
	{8'd62,8'd180} : s = 331;
	{8'd62,8'd181} : s = 441;
	{8'd62,8'd182} : s = 327;
	{8'd62,8'd183} : s = 438;
	{8'd62,8'd184} : s = 437;
	{8'd62,8'd185} : s = 501;
	{8'd62,8'd186} : s = 316;
	{8'd62,8'd187} : s = 435;
	{8'd62,8'd188} : s = 430;
	{8'd62,8'd189} : s = 499;
	{8'd62,8'd190} : s = 429;
	{8'd62,8'd191} : s = 494;
	{8'd62,8'd192} : s = 493;
	{8'd62,8'd193} : s = 510;
	{8'd62,8'd194} : s = 1;
	{8'd62,8'd195} : s = 18;
	{8'd62,8'd196} : s = 17;
	{8'd62,8'd197} : s = 82;
	{8'd62,8'd198} : s = 12;
	{8'd62,8'd199} : s = 81;
	{8'd62,8'd200} : s = 76;
	{8'd62,8'd201} : s = 195;
	{8'd62,8'd202} : s = 10;
	{8'd62,8'd203} : s = 74;
	{8'd62,8'd204} : s = 73;
	{8'd62,8'd205} : s = 184;
	{8'd62,8'd206} : s = 70;
	{8'd62,8'd207} : s = 180;
	{8'd62,8'd208} : s = 178;
	{8'd62,8'd209} : s = 314;
	{8'd62,8'd210} : s = 9;
	{8'd62,8'd211} : s = 69;
	{8'd62,8'd212} : s = 67;
	{8'd62,8'd213} : s = 177;
	{8'd62,8'd214} : s = 56;
	{8'd62,8'd215} : s = 172;
	{8'd62,8'd216} : s = 170;
	{8'd62,8'd217} : s = 313;
	{8'd62,8'd218} : s = 52;
	{8'd62,8'd219} : s = 169;
	{8'd62,8'd220} : s = 166;
	{8'd62,8'd221} : s = 310;
	{8'd62,8'd222} : s = 165;
	{8'd62,8'd223} : s = 309;
	{8'd62,8'd224} : s = 307;
	{8'd62,8'd225} : s = 427;
	{8'd62,8'd226} : s = 6;
	{8'd62,8'd227} : s = 50;
	{8'd62,8'd228} : s = 49;
	{8'd62,8'd229} : s = 163;
	{8'd62,8'd230} : s = 44;
	{8'd62,8'd231} : s = 156;
	{8'd62,8'd232} : s = 154;
	{8'd62,8'd233} : s = 302;
	{8'd62,8'd234} : s = 42;
	{8'd62,8'd235} : s = 153;
	{8'd62,8'd236} : s = 150;
	{8'd62,8'd237} : s = 301;
	{8'd62,8'd238} : s = 149;
	{8'd62,8'd239} : s = 299;
	{8'd62,8'd240} : s = 295;
	{8'd62,8'd241} : s = 423;
	{8'd62,8'd242} : s = 41;
	{8'd62,8'd243} : s = 147;
	{8'd62,8'd244} : s = 142;
	{8'd62,8'd245} : s = 286;
	{8'd62,8'd246} : s = 141;
	{8'd62,8'd247} : s = 285;
	{8'd62,8'd248} : s = 283;
	{8'd62,8'd249} : s = 414;
	{8'd62,8'd250} : s = 139;
	{8'd62,8'd251} : s = 279;
	{8'd62,8'd252} : s = 271;
	{8'd62,8'd253} : s = 413;
	{8'd62,8'd254} : s = 248;
	{8'd62,8'd255} : s = 411;
	{8'd63,8'd0} : s = 504;
	{8'd63,8'd1} : s = 4;
	{8'd63,8'd2} : s = 96;
	{8'd63,8'd3} : s = 80;
	{8'd63,8'd4} : s = 274;
	{8'd63,8'd5} : s = 72;
	{8'd63,8'd6} : s = 273;
	{8'd63,8'd7} : s = 268;
	{8'd63,8'd8} : s = 396;
	{8'd63,8'd9} : s = 68;
	{8'd63,8'd10} : s = 266;
	{8'd63,8'd11} : s = 265;
	{8'd63,8'd12} : s = 394;
	{8'd63,8'd13} : s = 262;
	{8'd63,8'd14} : s = 393;
	{8'd63,8'd15} : s = 390;
	{8'd63,8'd16} : s = 468;
	{8'd63,8'd17} : s = 66;
	{8'd63,8'd18} : s = 261;
	{8'd63,8'd19} : s = 259;
	{8'd63,8'd20} : s = 389;
	{8'd63,8'd21} : s = 224;
	{8'd63,8'd22} : s = 387;
	{8'd63,8'd23} : s = 368;
	{8'd63,8'd24} : s = 466;
	{8'd63,8'd25} : s = 208;
	{8'd63,8'd26} : s = 360;
	{8'd63,8'd27} : s = 356;
	{8'd63,8'd28} : s = 465;
	{8'd63,8'd29} : s = 354;
	{8'd63,8'd30} : s = 460;
	{8'd63,8'd31} : s = 458;
	{8'd63,8'd32} : s = 500;
	{8'd63,8'd33} : s = 65;
	{8'd63,8'd34} : s = 200;
	{8'd63,8'd35} : s = 196;
	{8'd63,8'd36} : s = 353;
	{8'd63,8'd37} : s = 194;
	{8'd63,8'd38} : s = 344;
	{8'd63,8'd39} : s = 340;
	{8'd63,8'd40} : s = 457;
	{8'd63,8'd41} : s = 193;
	{8'd63,8'd42} : s = 338;
	{8'd63,8'd43} : s = 337;
	{8'd63,8'd44} : s = 454;
	{8'd63,8'd45} : s = 332;
	{8'd63,8'd46} : s = 453;
	{8'd63,8'd47} : s = 451;
	{8'd63,8'd48} : s = 498;
	{8'd63,8'd49} : s = 176;
	{8'd63,8'd50} : s = 330;
	{8'd63,8'd51} : s = 329;
	{8'd63,8'd52} : s = 440;
	{8'd63,8'd53} : s = 326;
	{8'd63,8'd54} : s = 436;
	{8'd63,8'd55} : s = 434;
	{8'd63,8'd56} : s = 497;
	{8'd63,8'd57} : s = 325;
	{8'd63,8'd58} : s = 433;
	{8'd63,8'd59} : s = 428;
	{8'd63,8'd60} : s = 492;
	{8'd63,8'd61} : s = 426;
	{8'd63,8'd62} : s = 490;
	{8'd63,8'd63} : s = 489;
	{8'd63,8'd64} : s = 508;
	{8'd63,8'd65} : s = 2;
	{8'd63,8'd66} : s = 48;
	{8'd63,8'd67} : s = 40;
	{8'd63,8'd68} : s = 168;
	{8'd63,8'd69} : s = 36;
	{8'd63,8'd70} : s = 164;
	{8'd63,8'd71} : s = 162;
	{8'd63,8'd72} : s = 323;
	{8'd63,8'd73} : s = 34;
	{8'd63,8'd74} : s = 161;
	{8'd63,8'd75} : s = 152;
	{8'd63,8'd76} : s = 312;
	{8'd63,8'd77} : s = 148;
	{8'd63,8'd78} : s = 308;
	{8'd63,8'd79} : s = 306;
	{8'd63,8'd80} : s = 425;
	{8'd63,8'd81} : s = 33;
	{8'd63,8'd82} : s = 146;
	{8'd63,8'd83} : s = 145;
	{8'd63,8'd84} : s = 305;
	{8'd63,8'd85} : s = 140;
	{8'd63,8'd86} : s = 300;
	{8'd63,8'd87} : s = 298;
	{8'd63,8'd88} : s = 422;
	{8'd63,8'd89} : s = 138;
	{8'd63,8'd90} : s = 297;
	{8'd63,8'd91} : s = 294;
	{8'd63,8'd92} : s = 421;
	{8'd63,8'd93} : s = 293;
	{8'd63,8'd94} : s = 419;
	{8'd63,8'd95} : s = 412;
	{8'd63,8'd96} : s = 486;
	{8'd63,8'd97} : s = 24;
	{8'd63,8'd98} : s = 137;
	{8'd63,8'd99} : s = 134;
	{8'd63,8'd100} : s = 291;
	{8'd63,8'd101} : s = 133;
	{8'd63,8'd102} : s = 284;
	{8'd63,8'd103} : s = 282;
	{8'd63,8'd104} : s = 410;
	{8'd63,8'd105} : s = 131;
	{8'd63,8'd106} : s = 281;
	{8'd63,8'd107} : s = 278;
	{8'd63,8'd108} : s = 409;
	{8'd63,8'd109} : s = 277;
	{8'd63,8'd110} : s = 406;
	{8'd63,8'd111} : s = 405;
	{8'd63,8'd112} : s = 485;
	{8'd63,8'd113} : s = 112;
	{8'd63,8'd114} : s = 275;
	{8'd63,8'd115} : s = 270;
	{8'd63,8'd116} : s = 403;
	{8'd63,8'd117} : s = 269;
	{8'd63,8'd118} : s = 398;
	{8'd63,8'd119} : s = 397;
	{8'd63,8'd120} : s = 483;
	{8'd63,8'd121} : s = 267;
	{8'd63,8'd122} : s = 395;
	{8'd63,8'd123} : s = 391;
	{8'd63,8'd124} : s = 476;
	{8'd63,8'd125} : s = 376;
	{8'd63,8'd126} : s = 474;
	{8'd63,8'd127} : s = 473;
	{8'd63,8'd128} : s = 506;
	{8'd63,8'd129} : s = 20;
	{8'd63,8'd130} : s = 104;
	{8'd63,8'd131} : s = 100;
	{8'd63,8'd132} : s = 263;
	{8'd63,8'd133} : s = 98;
	{8'd63,8'd134} : s = 240;
	{8'd63,8'd135} : s = 232;
	{8'd63,8'd136} : s = 372;
	{8'd63,8'd137} : s = 97;
	{8'd63,8'd138} : s = 228;
	{8'd63,8'd139} : s = 226;
	{8'd63,8'd140} : s = 370;
	{8'd63,8'd141} : s = 225;
	{8'd63,8'd142} : s = 369;
	{8'd63,8'd143} : s = 364;
	{8'd63,8'd144} : s = 470;
	{8'd63,8'd145} : s = 88;
	{8'd63,8'd146} : s = 216;
	{8'd63,8'd147} : s = 212;
	{8'd63,8'd148} : s = 362;
	{8'd63,8'd149} : s = 210;
	{8'd63,8'd150} : s = 361;
	{8'd63,8'd151} : s = 358;
	{8'd63,8'd152} : s = 469;
	{8'd63,8'd153} : s = 209;
	{8'd63,8'd154} : s = 357;
	{8'd63,8'd155} : s = 355;
	{8'd63,8'd156} : s = 467;
	{8'd63,8'd157} : s = 348;
	{8'd63,8'd158} : s = 462;
	{8'd63,8'd159} : s = 461;
	{8'd63,8'd160} : s = 505;
	{8'd63,8'd161} : s = 84;
	{8'd63,8'd162} : s = 204;
	{8'd63,8'd163} : s = 202;
	{8'd63,8'd164} : s = 346;
	{8'd63,8'd165} : s = 201;
	{8'd63,8'd166} : s = 345;
	{8'd63,8'd167} : s = 342;
	{8'd63,8'd168} : s = 459;
	{8'd63,8'd169} : s = 198;
	{8'd63,8'd170} : s = 341;
	{8'd63,8'd171} : s = 339;
	{8'd63,8'd172} : s = 455;
	{8'd63,8'd173} : s = 334;
	{8'd63,8'd174} : s = 444;
	{8'd63,8'd175} : s = 442;
	{8'd63,8'd176} : s = 502;
	{8'd63,8'd177} : s = 197;
	{8'd63,8'd178} : s = 333;
	{8'd63,8'd179} : s = 331;
	{8'd63,8'd180} : s = 441;
	{8'd63,8'd181} : s = 327;
	{8'd63,8'd182} : s = 438;
	{8'd63,8'd183} : s = 437;
	{8'd63,8'd184} : s = 501;
	{8'd63,8'd185} : s = 316;
	{8'd63,8'd186} : s = 435;
	{8'd63,8'd187} : s = 430;
	{8'd63,8'd188} : s = 499;
	{8'd63,8'd189} : s = 429;
	{8'd63,8'd190} : s = 494;
	{8'd63,8'd191} : s = 493;
	{8'd63,8'd192} : s = 510;
	{8'd63,8'd193} : s = 1;
	{8'd63,8'd194} : s = 18;
	{8'd63,8'd195} : s = 17;
	{8'd63,8'd196} : s = 82;
	{8'd63,8'd197} : s = 12;
	{8'd63,8'd198} : s = 81;
	{8'd63,8'd199} : s = 76;
	{8'd63,8'd200} : s = 195;
	{8'd63,8'd201} : s = 10;
	{8'd63,8'd202} : s = 74;
	{8'd63,8'd203} : s = 73;
	{8'd63,8'd204} : s = 184;
	{8'd63,8'd205} : s = 70;
	{8'd63,8'd206} : s = 180;
	{8'd63,8'd207} : s = 178;
	{8'd63,8'd208} : s = 314;
	{8'd63,8'd209} : s = 9;
	{8'd63,8'd210} : s = 69;
	{8'd63,8'd211} : s = 67;
	{8'd63,8'd212} : s = 177;
	{8'd63,8'd213} : s = 56;
	{8'd63,8'd214} : s = 172;
	{8'd63,8'd215} : s = 170;
	{8'd63,8'd216} : s = 313;
	{8'd63,8'd217} : s = 52;
	{8'd63,8'd218} : s = 169;
	{8'd63,8'd219} : s = 166;
	{8'd63,8'd220} : s = 310;
	{8'd63,8'd221} : s = 165;
	{8'd63,8'd222} : s = 309;
	{8'd63,8'd223} : s = 307;
	{8'd63,8'd224} : s = 427;
	{8'd63,8'd225} : s = 6;
	{8'd63,8'd226} : s = 50;
	{8'd63,8'd227} : s = 49;
	{8'd63,8'd228} : s = 163;
	{8'd63,8'd229} : s = 44;
	{8'd63,8'd230} : s = 156;
	{8'd63,8'd231} : s = 154;
	{8'd63,8'd232} : s = 302;
	{8'd63,8'd233} : s = 42;
	{8'd63,8'd234} : s = 153;
	{8'd63,8'd235} : s = 150;
	{8'd63,8'd236} : s = 301;
	{8'd63,8'd237} : s = 149;
	{8'd63,8'd238} : s = 299;
	{8'd63,8'd239} : s = 295;
	{8'd63,8'd240} : s = 423;
	{8'd63,8'd241} : s = 41;
	{8'd63,8'd242} : s = 147;
	{8'd63,8'd243} : s = 142;
	{8'd63,8'd244} : s = 286;
	{8'd63,8'd245} : s = 141;
	{8'd63,8'd246} : s = 285;
	{8'd63,8'd247} : s = 283;
	{8'd63,8'd248} : s = 414;
	{8'd63,8'd249} : s = 139;
	{8'd63,8'd250} : s = 279;
	{8'd63,8'd251} : s = 271;
	{8'd63,8'd252} : s = 413;
	{8'd63,8'd253} : s = 248;
	{8'd63,8'd254} : s = 411;
	{8'd63,8'd255} : s = 407;
	{8'd64,8'd0} : s = 4;
	{8'd64,8'd1} : s = 96;
	{8'd64,8'd2} : s = 80;
	{8'd64,8'd3} : s = 274;
	{8'd64,8'd4} : s = 72;
	{8'd64,8'd5} : s = 273;
	{8'd64,8'd6} : s = 268;
	{8'd64,8'd7} : s = 396;
	{8'd64,8'd8} : s = 68;
	{8'd64,8'd9} : s = 266;
	{8'd64,8'd10} : s = 265;
	{8'd64,8'd11} : s = 394;
	{8'd64,8'd12} : s = 262;
	{8'd64,8'd13} : s = 393;
	{8'd64,8'd14} : s = 390;
	{8'd64,8'd15} : s = 468;
	{8'd64,8'd16} : s = 66;
	{8'd64,8'd17} : s = 261;
	{8'd64,8'd18} : s = 259;
	{8'd64,8'd19} : s = 389;
	{8'd64,8'd20} : s = 224;
	{8'd64,8'd21} : s = 387;
	{8'd64,8'd22} : s = 368;
	{8'd64,8'd23} : s = 466;
	{8'd64,8'd24} : s = 208;
	{8'd64,8'd25} : s = 360;
	{8'd64,8'd26} : s = 356;
	{8'd64,8'd27} : s = 465;
	{8'd64,8'd28} : s = 354;
	{8'd64,8'd29} : s = 460;
	{8'd64,8'd30} : s = 458;
	{8'd64,8'd31} : s = 500;
	{8'd64,8'd32} : s = 65;
	{8'd64,8'd33} : s = 200;
	{8'd64,8'd34} : s = 196;
	{8'd64,8'd35} : s = 353;
	{8'd64,8'd36} : s = 194;
	{8'd64,8'd37} : s = 344;
	{8'd64,8'd38} : s = 340;
	{8'd64,8'd39} : s = 457;
	{8'd64,8'd40} : s = 193;
	{8'd64,8'd41} : s = 338;
	{8'd64,8'd42} : s = 337;
	{8'd64,8'd43} : s = 454;
	{8'd64,8'd44} : s = 332;
	{8'd64,8'd45} : s = 453;
	{8'd64,8'd46} : s = 451;
	{8'd64,8'd47} : s = 498;
	{8'd64,8'd48} : s = 176;
	{8'd64,8'd49} : s = 330;
	{8'd64,8'd50} : s = 329;
	{8'd64,8'd51} : s = 440;
	{8'd64,8'd52} : s = 326;
	{8'd64,8'd53} : s = 436;
	{8'd64,8'd54} : s = 434;
	{8'd64,8'd55} : s = 497;
	{8'd64,8'd56} : s = 325;
	{8'd64,8'd57} : s = 433;
	{8'd64,8'd58} : s = 428;
	{8'd64,8'd59} : s = 492;
	{8'd64,8'd60} : s = 426;
	{8'd64,8'd61} : s = 490;
	{8'd64,8'd62} : s = 489;
	{8'd64,8'd63} : s = 508;
	{8'd64,8'd64} : s = 2;
	{8'd64,8'd65} : s = 48;
	{8'd64,8'd66} : s = 40;
	{8'd64,8'd67} : s = 168;
	{8'd64,8'd68} : s = 36;
	{8'd64,8'd69} : s = 164;
	{8'd64,8'd70} : s = 162;
	{8'd64,8'd71} : s = 323;
	{8'd64,8'd72} : s = 34;
	{8'd64,8'd73} : s = 161;
	{8'd64,8'd74} : s = 152;
	{8'd64,8'd75} : s = 312;
	{8'd64,8'd76} : s = 148;
	{8'd64,8'd77} : s = 308;
	{8'd64,8'd78} : s = 306;
	{8'd64,8'd79} : s = 425;
	{8'd64,8'd80} : s = 33;
	{8'd64,8'd81} : s = 146;
	{8'd64,8'd82} : s = 145;
	{8'd64,8'd83} : s = 305;
	{8'd64,8'd84} : s = 140;
	{8'd64,8'd85} : s = 300;
	{8'd64,8'd86} : s = 298;
	{8'd64,8'd87} : s = 422;
	{8'd64,8'd88} : s = 138;
	{8'd64,8'd89} : s = 297;
	{8'd64,8'd90} : s = 294;
	{8'd64,8'd91} : s = 421;
	{8'd64,8'd92} : s = 293;
	{8'd64,8'd93} : s = 419;
	{8'd64,8'd94} : s = 412;
	{8'd64,8'd95} : s = 486;
	{8'd64,8'd96} : s = 24;
	{8'd64,8'd97} : s = 137;
	{8'd64,8'd98} : s = 134;
	{8'd64,8'd99} : s = 291;
	{8'd64,8'd100} : s = 133;
	{8'd64,8'd101} : s = 284;
	{8'd64,8'd102} : s = 282;
	{8'd64,8'd103} : s = 410;
	{8'd64,8'd104} : s = 131;
	{8'd64,8'd105} : s = 281;
	{8'd64,8'd106} : s = 278;
	{8'd64,8'd107} : s = 409;
	{8'd64,8'd108} : s = 277;
	{8'd64,8'd109} : s = 406;
	{8'd64,8'd110} : s = 405;
	{8'd64,8'd111} : s = 485;
	{8'd64,8'd112} : s = 112;
	{8'd64,8'd113} : s = 275;
	{8'd64,8'd114} : s = 270;
	{8'd64,8'd115} : s = 403;
	{8'd64,8'd116} : s = 269;
	{8'd64,8'd117} : s = 398;
	{8'd64,8'd118} : s = 397;
	{8'd64,8'd119} : s = 483;
	{8'd64,8'd120} : s = 267;
	{8'd64,8'd121} : s = 395;
	{8'd64,8'd122} : s = 391;
	{8'd64,8'd123} : s = 476;
	{8'd64,8'd124} : s = 376;
	{8'd64,8'd125} : s = 474;
	{8'd64,8'd126} : s = 473;
	{8'd64,8'd127} : s = 506;
	{8'd64,8'd128} : s = 20;
	{8'd64,8'd129} : s = 104;
	{8'd64,8'd130} : s = 100;
	{8'd64,8'd131} : s = 263;
	{8'd64,8'd132} : s = 98;
	{8'd64,8'd133} : s = 240;
	{8'd64,8'd134} : s = 232;
	{8'd64,8'd135} : s = 372;
	{8'd64,8'd136} : s = 97;
	{8'd64,8'd137} : s = 228;
	{8'd64,8'd138} : s = 226;
	{8'd64,8'd139} : s = 370;
	{8'd64,8'd140} : s = 225;
	{8'd64,8'd141} : s = 369;
	{8'd64,8'd142} : s = 364;
	{8'd64,8'd143} : s = 470;
	{8'd64,8'd144} : s = 88;
	{8'd64,8'd145} : s = 216;
	{8'd64,8'd146} : s = 212;
	{8'd64,8'd147} : s = 362;
	{8'd64,8'd148} : s = 210;
	{8'd64,8'd149} : s = 361;
	{8'd64,8'd150} : s = 358;
	{8'd64,8'd151} : s = 469;
	{8'd64,8'd152} : s = 209;
	{8'd64,8'd153} : s = 357;
	{8'd64,8'd154} : s = 355;
	{8'd64,8'd155} : s = 467;
	{8'd64,8'd156} : s = 348;
	{8'd64,8'd157} : s = 462;
	{8'd64,8'd158} : s = 461;
	{8'd64,8'd159} : s = 505;
	{8'd64,8'd160} : s = 84;
	{8'd64,8'd161} : s = 204;
	{8'd64,8'd162} : s = 202;
	{8'd64,8'd163} : s = 346;
	{8'd64,8'd164} : s = 201;
	{8'd64,8'd165} : s = 345;
	{8'd64,8'd166} : s = 342;
	{8'd64,8'd167} : s = 459;
	{8'd64,8'd168} : s = 198;
	{8'd64,8'd169} : s = 341;
	{8'd64,8'd170} : s = 339;
	{8'd64,8'd171} : s = 455;
	{8'd64,8'd172} : s = 334;
	{8'd64,8'd173} : s = 444;
	{8'd64,8'd174} : s = 442;
	{8'd64,8'd175} : s = 502;
	{8'd64,8'd176} : s = 197;
	{8'd64,8'd177} : s = 333;
	{8'd64,8'd178} : s = 331;
	{8'd64,8'd179} : s = 441;
	{8'd64,8'd180} : s = 327;
	{8'd64,8'd181} : s = 438;
	{8'd64,8'd182} : s = 437;
	{8'd64,8'd183} : s = 501;
	{8'd64,8'd184} : s = 316;
	{8'd64,8'd185} : s = 435;
	{8'd64,8'd186} : s = 430;
	{8'd64,8'd187} : s = 499;
	{8'd64,8'd188} : s = 429;
	{8'd64,8'd189} : s = 494;
	{8'd64,8'd190} : s = 493;
	{8'd64,8'd191} : s = 510;
	{8'd64,8'd192} : s = 1;
	{8'd64,8'd193} : s = 18;
	{8'd64,8'd194} : s = 17;
	{8'd64,8'd195} : s = 82;
	{8'd64,8'd196} : s = 12;
	{8'd64,8'd197} : s = 81;
	{8'd64,8'd198} : s = 76;
	{8'd64,8'd199} : s = 195;
	{8'd64,8'd200} : s = 10;
	{8'd64,8'd201} : s = 74;
	{8'd64,8'd202} : s = 73;
	{8'd64,8'd203} : s = 184;
	{8'd64,8'd204} : s = 70;
	{8'd64,8'd205} : s = 180;
	{8'd64,8'd206} : s = 178;
	{8'd64,8'd207} : s = 314;
	{8'd64,8'd208} : s = 9;
	{8'd64,8'd209} : s = 69;
	{8'd64,8'd210} : s = 67;
	{8'd64,8'd211} : s = 177;
	{8'd64,8'd212} : s = 56;
	{8'd64,8'd213} : s = 172;
	{8'd64,8'd214} : s = 170;
	{8'd64,8'd215} : s = 313;
	{8'd64,8'd216} : s = 52;
	{8'd64,8'd217} : s = 169;
	{8'd64,8'd218} : s = 166;
	{8'd64,8'd219} : s = 310;
	{8'd64,8'd220} : s = 165;
	{8'd64,8'd221} : s = 309;
	{8'd64,8'd222} : s = 307;
	{8'd64,8'd223} : s = 427;
	{8'd64,8'd224} : s = 6;
	{8'd64,8'd225} : s = 50;
	{8'd64,8'd226} : s = 49;
	{8'd64,8'd227} : s = 163;
	{8'd64,8'd228} : s = 44;
	{8'd64,8'd229} : s = 156;
	{8'd64,8'd230} : s = 154;
	{8'd64,8'd231} : s = 302;
	{8'd64,8'd232} : s = 42;
	{8'd64,8'd233} : s = 153;
	{8'd64,8'd234} : s = 150;
	{8'd64,8'd235} : s = 301;
	{8'd64,8'd236} : s = 149;
	{8'd64,8'd237} : s = 299;
	{8'd64,8'd238} : s = 295;
	{8'd64,8'd239} : s = 423;
	{8'd64,8'd240} : s = 41;
	{8'd64,8'd241} : s = 147;
	{8'd64,8'd242} : s = 142;
	{8'd64,8'd243} : s = 286;
	{8'd64,8'd244} : s = 141;
	{8'd64,8'd245} : s = 285;
	{8'd64,8'd246} : s = 283;
	{8'd64,8'd247} : s = 414;
	{8'd64,8'd248} : s = 139;
	{8'd64,8'd249} : s = 279;
	{8'd64,8'd250} : s = 271;
	{8'd64,8'd251} : s = 413;
	{8'd64,8'd252} : s = 248;
	{8'd64,8'd253} : s = 411;
	{8'd64,8'd254} : s = 407;
	{8'd64,8'd255} : s = 491;
	{8'd65,8'd0} : s = 96;
	{8'd65,8'd1} : s = 80;
	{8'd65,8'd2} : s = 274;
	{8'd65,8'd3} : s = 72;
	{8'd65,8'd4} : s = 273;
	{8'd65,8'd5} : s = 268;
	{8'd65,8'd6} : s = 396;
	{8'd65,8'd7} : s = 68;
	{8'd65,8'd8} : s = 266;
	{8'd65,8'd9} : s = 265;
	{8'd65,8'd10} : s = 394;
	{8'd65,8'd11} : s = 262;
	{8'd65,8'd12} : s = 393;
	{8'd65,8'd13} : s = 390;
	{8'd65,8'd14} : s = 468;
	{8'd65,8'd15} : s = 66;
	{8'd65,8'd16} : s = 261;
	{8'd65,8'd17} : s = 259;
	{8'd65,8'd18} : s = 389;
	{8'd65,8'd19} : s = 224;
	{8'd65,8'd20} : s = 387;
	{8'd65,8'd21} : s = 368;
	{8'd65,8'd22} : s = 466;
	{8'd65,8'd23} : s = 208;
	{8'd65,8'd24} : s = 360;
	{8'd65,8'd25} : s = 356;
	{8'd65,8'd26} : s = 465;
	{8'd65,8'd27} : s = 354;
	{8'd65,8'd28} : s = 460;
	{8'd65,8'd29} : s = 458;
	{8'd65,8'd30} : s = 500;
	{8'd65,8'd31} : s = 65;
	{8'd65,8'd32} : s = 200;
	{8'd65,8'd33} : s = 196;
	{8'd65,8'd34} : s = 353;
	{8'd65,8'd35} : s = 194;
	{8'd65,8'd36} : s = 344;
	{8'd65,8'd37} : s = 340;
	{8'd65,8'd38} : s = 457;
	{8'd65,8'd39} : s = 193;
	{8'd65,8'd40} : s = 338;
	{8'd65,8'd41} : s = 337;
	{8'd65,8'd42} : s = 454;
	{8'd65,8'd43} : s = 332;
	{8'd65,8'd44} : s = 453;
	{8'd65,8'd45} : s = 451;
	{8'd65,8'd46} : s = 498;
	{8'd65,8'd47} : s = 176;
	{8'd65,8'd48} : s = 330;
	{8'd65,8'd49} : s = 329;
	{8'd65,8'd50} : s = 440;
	{8'd65,8'd51} : s = 326;
	{8'd65,8'd52} : s = 436;
	{8'd65,8'd53} : s = 434;
	{8'd65,8'd54} : s = 497;
	{8'd65,8'd55} : s = 325;
	{8'd65,8'd56} : s = 433;
	{8'd65,8'd57} : s = 428;
	{8'd65,8'd58} : s = 492;
	{8'd65,8'd59} : s = 426;
	{8'd65,8'd60} : s = 490;
	{8'd65,8'd61} : s = 489;
	{8'd65,8'd62} : s = 508;
	{8'd65,8'd63} : s = 2;
	{8'd65,8'd64} : s = 48;
	{8'd65,8'd65} : s = 40;
	{8'd65,8'd66} : s = 168;
	{8'd65,8'd67} : s = 36;
	{8'd65,8'd68} : s = 164;
	{8'd65,8'd69} : s = 162;
	{8'd65,8'd70} : s = 323;
	{8'd65,8'd71} : s = 34;
	{8'd65,8'd72} : s = 161;
	{8'd65,8'd73} : s = 152;
	{8'd65,8'd74} : s = 312;
	{8'd65,8'd75} : s = 148;
	{8'd65,8'd76} : s = 308;
	{8'd65,8'd77} : s = 306;
	{8'd65,8'd78} : s = 425;
	{8'd65,8'd79} : s = 33;
	{8'd65,8'd80} : s = 146;
	{8'd65,8'd81} : s = 145;
	{8'd65,8'd82} : s = 305;
	{8'd65,8'd83} : s = 140;
	{8'd65,8'd84} : s = 300;
	{8'd65,8'd85} : s = 298;
	{8'd65,8'd86} : s = 422;
	{8'd65,8'd87} : s = 138;
	{8'd65,8'd88} : s = 297;
	{8'd65,8'd89} : s = 294;
	{8'd65,8'd90} : s = 421;
	{8'd65,8'd91} : s = 293;
	{8'd65,8'd92} : s = 419;
	{8'd65,8'd93} : s = 412;
	{8'd65,8'd94} : s = 486;
	{8'd65,8'd95} : s = 24;
	{8'd65,8'd96} : s = 137;
	{8'd65,8'd97} : s = 134;
	{8'd65,8'd98} : s = 291;
	{8'd65,8'd99} : s = 133;
	{8'd65,8'd100} : s = 284;
	{8'd65,8'd101} : s = 282;
	{8'd65,8'd102} : s = 410;
	{8'd65,8'd103} : s = 131;
	{8'd65,8'd104} : s = 281;
	{8'd65,8'd105} : s = 278;
	{8'd65,8'd106} : s = 409;
	{8'd65,8'd107} : s = 277;
	{8'd65,8'd108} : s = 406;
	{8'd65,8'd109} : s = 405;
	{8'd65,8'd110} : s = 485;
	{8'd65,8'd111} : s = 112;
	{8'd65,8'd112} : s = 275;
	{8'd65,8'd113} : s = 270;
	{8'd65,8'd114} : s = 403;
	{8'd65,8'd115} : s = 269;
	{8'd65,8'd116} : s = 398;
	{8'd65,8'd117} : s = 397;
	{8'd65,8'd118} : s = 483;
	{8'd65,8'd119} : s = 267;
	{8'd65,8'd120} : s = 395;
	{8'd65,8'd121} : s = 391;
	{8'd65,8'd122} : s = 476;
	{8'd65,8'd123} : s = 376;
	{8'd65,8'd124} : s = 474;
	{8'd65,8'd125} : s = 473;
	{8'd65,8'd126} : s = 506;
	{8'd65,8'd127} : s = 20;
	{8'd65,8'd128} : s = 104;
	{8'd65,8'd129} : s = 100;
	{8'd65,8'd130} : s = 263;
	{8'd65,8'd131} : s = 98;
	{8'd65,8'd132} : s = 240;
	{8'd65,8'd133} : s = 232;
	{8'd65,8'd134} : s = 372;
	{8'd65,8'd135} : s = 97;
	{8'd65,8'd136} : s = 228;
	{8'd65,8'd137} : s = 226;
	{8'd65,8'd138} : s = 370;
	{8'd65,8'd139} : s = 225;
	{8'd65,8'd140} : s = 369;
	{8'd65,8'd141} : s = 364;
	{8'd65,8'd142} : s = 470;
	{8'd65,8'd143} : s = 88;
	{8'd65,8'd144} : s = 216;
	{8'd65,8'd145} : s = 212;
	{8'd65,8'd146} : s = 362;
	{8'd65,8'd147} : s = 210;
	{8'd65,8'd148} : s = 361;
	{8'd65,8'd149} : s = 358;
	{8'd65,8'd150} : s = 469;
	{8'd65,8'd151} : s = 209;
	{8'd65,8'd152} : s = 357;
	{8'd65,8'd153} : s = 355;
	{8'd65,8'd154} : s = 467;
	{8'd65,8'd155} : s = 348;
	{8'd65,8'd156} : s = 462;
	{8'd65,8'd157} : s = 461;
	{8'd65,8'd158} : s = 505;
	{8'd65,8'd159} : s = 84;
	{8'd65,8'd160} : s = 204;
	{8'd65,8'd161} : s = 202;
	{8'd65,8'd162} : s = 346;
	{8'd65,8'd163} : s = 201;
	{8'd65,8'd164} : s = 345;
	{8'd65,8'd165} : s = 342;
	{8'd65,8'd166} : s = 459;
	{8'd65,8'd167} : s = 198;
	{8'd65,8'd168} : s = 341;
	{8'd65,8'd169} : s = 339;
	{8'd65,8'd170} : s = 455;
	{8'd65,8'd171} : s = 334;
	{8'd65,8'd172} : s = 444;
	{8'd65,8'd173} : s = 442;
	{8'd65,8'd174} : s = 502;
	{8'd65,8'd175} : s = 197;
	{8'd65,8'd176} : s = 333;
	{8'd65,8'd177} : s = 331;
	{8'd65,8'd178} : s = 441;
	{8'd65,8'd179} : s = 327;
	{8'd65,8'd180} : s = 438;
	{8'd65,8'd181} : s = 437;
	{8'd65,8'd182} : s = 501;
	{8'd65,8'd183} : s = 316;
	{8'd65,8'd184} : s = 435;
	{8'd65,8'd185} : s = 430;
	{8'd65,8'd186} : s = 499;
	{8'd65,8'd187} : s = 429;
	{8'd65,8'd188} : s = 494;
	{8'd65,8'd189} : s = 493;
	{8'd65,8'd190} : s = 510;
	{8'd65,8'd191} : s = 1;
	{8'd65,8'd192} : s = 18;
	{8'd65,8'd193} : s = 17;
	{8'd65,8'd194} : s = 82;
	{8'd65,8'd195} : s = 12;
	{8'd65,8'd196} : s = 81;
	{8'd65,8'd197} : s = 76;
	{8'd65,8'd198} : s = 195;
	{8'd65,8'd199} : s = 10;
	{8'd65,8'd200} : s = 74;
	{8'd65,8'd201} : s = 73;
	{8'd65,8'd202} : s = 184;
	{8'd65,8'd203} : s = 70;
	{8'd65,8'd204} : s = 180;
	{8'd65,8'd205} : s = 178;
	{8'd65,8'd206} : s = 314;
	{8'd65,8'd207} : s = 9;
	{8'd65,8'd208} : s = 69;
	{8'd65,8'd209} : s = 67;
	{8'd65,8'd210} : s = 177;
	{8'd65,8'd211} : s = 56;
	{8'd65,8'd212} : s = 172;
	{8'd65,8'd213} : s = 170;
	{8'd65,8'd214} : s = 313;
	{8'd65,8'd215} : s = 52;
	{8'd65,8'd216} : s = 169;
	{8'd65,8'd217} : s = 166;
	{8'd65,8'd218} : s = 310;
	{8'd65,8'd219} : s = 165;
	{8'd65,8'd220} : s = 309;
	{8'd65,8'd221} : s = 307;
	{8'd65,8'd222} : s = 427;
	{8'd65,8'd223} : s = 6;
	{8'd65,8'd224} : s = 50;
	{8'd65,8'd225} : s = 49;
	{8'd65,8'd226} : s = 163;
	{8'd65,8'd227} : s = 44;
	{8'd65,8'd228} : s = 156;
	{8'd65,8'd229} : s = 154;
	{8'd65,8'd230} : s = 302;
	{8'd65,8'd231} : s = 42;
	{8'd65,8'd232} : s = 153;
	{8'd65,8'd233} : s = 150;
	{8'd65,8'd234} : s = 301;
	{8'd65,8'd235} : s = 149;
	{8'd65,8'd236} : s = 299;
	{8'd65,8'd237} : s = 295;
	{8'd65,8'd238} : s = 423;
	{8'd65,8'd239} : s = 41;
	{8'd65,8'd240} : s = 147;
	{8'd65,8'd241} : s = 142;
	{8'd65,8'd242} : s = 286;
	{8'd65,8'd243} : s = 141;
	{8'd65,8'd244} : s = 285;
	{8'd65,8'd245} : s = 283;
	{8'd65,8'd246} : s = 414;
	{8'd65,8'd247} : s = 139;
	{8'd65,8'd248} : s = 279;
	{8'd65,8'd249} : s = 271;
	{8'd65,8'd250} : s = 413;
	{8'd65,8'd251} : s = 248;
	{8'd65,8'd252} : s = 411;
	{8'd65,8'd253} : s = 407;
	{8'd65,8'd254} : s = 491;
	{8'd65,8'd255} : s = 5;
	{8'd66,8'd0} : s = 80;
	{8'd66,8'd1} : s = 274;
	{8'd66,8'd2} : s = 72;
	{8'd66,8'd3} : s = 273;
	{8'd66,8'd4} : s = 268;
	{8'd66,8'd5} : s = 396;
	{8'd66,8'd6} : s = 68;
	{8'd66,8'd7} : s = 266;
	{8'd66,8'd8} : s = 265;
	{8'd66,8'd9} : s = 394;
	{8'd66,8'd10} : s = 262;
	{8'd66,8'd11} : s = 393;
	{8'd66,8'd12} : s = 390;
	{8'd66,8'd13} : s = 468;
	{8'd66,8'd14} : s = 66;
	{8'd66,8'd15} : s = 261;
	{8'd66,8'd16} : s = 259;
	{8'd66,8'd17} : s = 389;
	{8'd66,8'd18} : s = 224;
	{8'd66,8'd19} : s = 387;
	{8'd66,8'd20} : s = 368;
	{8'd66,8'd21} : s = 466;
	{8'd66,8'd22} : s = 208;
	{8'd66,8'd23} : s = 360;
	{8'd66,8'd24} : s = 356;
	{8'd66,8'd25} : s = 465;
	{8'd66,8'd26} : s = 354;
	{8'd66,8'd27} : s = 460;
	{8'd66,8'd28} : s = 458;
	{8'd66,8'd29} : s = 500;
	{8'd66,8'd30} : s = 65;
	{8'd66,8'd31} : s = 200;
	{8'd66,8'd32} : s = 196;
	{8'd66,8'd33} : s = 353;
	{8'd66,8'd34} : s = 194;
	{8'd66,8'd35} : s = 344;
	{8'd66,8'd36} : s = 340;
	{8'd66,8'd37} : s = 457;
	{8'd66,8'd38} : s = 193;
	{8'd66,8'd39} : s = 338;
	{8'd66,8'd40} : s = 337;
	{8'd66,8'd41} : s = 454;
	{8'd66,8'd42} : s = 332;
	{8'd66,8'd43} : s = 453;
	{8'd66,8'd44} : s = 451;
	{8'd66,8'd45} : s = 498;
	{8'd66,8'd46} : s = 176;
	{8'd66,8'd47} : s = 330;
	{8'd66,8'd48} : s = 329;
	{8'd66,8'd49} : s = 440;
	{8'd66,8'd50} : s = 326;
	{8'd66,8'd51} : s = 436;
	{8'd66,8'd52} : s = 434;
	{8'd66,8'd53} : s = 497;
	{8'd66,8'd54} : s = 325;
	{8'd66,8'd55} : s = 433;
	{8'd66,8'd56} : s = 428;
	{8'd66,8'd57} : s = 492;
	{8'd66,8'd58} : s = 426;
	{8'd66,8'd59} : s = 490;
	{8'd66,8'd60} : s = 489;
	{8'd66,8'd61} : s = 508;
	{8'd66,8'd62} : s = 2;
	{8'd66,8'd63} : s = 48;
	{8'd66,8'd64} : s = 40;
	{8'd66,8'd65} : s = 168;
	{8'd66,8'd66} : s = 36;
	{8'd66,8'd67} : s = 164;
	{8'd66,8'd68} : s = 162;
	{8'd66,8'd69} : s = 323;
	{8'd66,8'd70} : s = 34;
	{8'd66,8'd71} : s = 161;
	{8'd66,8'd72} : s = 152;
	{8'd66,8'd73} : s = 312;
	{8'd66,8'd74} : s = 148;
	{8'd66,8'd75} : s = 308;
	{8'd66,8'd76} : s = 306;
	{8'd66,8'd77} : s = 425;
	{8'd66,8'd78} : s = 33;
	{8'd66,8'd79} : s = 146;
	{8'd66,8'd80} : s = 145;
	{8'd66,8'd81} : s = 305;
	{8'd66,8'd82} : s = 140;
	{8'd66,8'd83} : s = 300;
	{8'd66,8'd84} : s = 298;
	{8'd66,8'd85} : s = 422;
	{8'd66,8'd86} : s = 138;
	{8'd66,8'd87} : s = 297;
	{8'd66,8'd88} : s = 294;
	{8'd66,8'd89} : s = 421;
	{8'd66,8'd90} : s = 293;
	{8'd66,8'd91} : s = 419;
	{8'd66,8'd92} : s = 412;
	{8'd66,8'd93} : s = 486;
	{8'd66,8'd94} : s = 24;
	{8'd66,8'd95} : s = 137;
	{8'd66,8'd96} : s = 134;
	{8'd66,8'd97} : s = 291;
	{8'd66,8'd98} : s = 133;
	{8'd66,8'd99} : s = 284;
	{8'd66,8'd100} : s = 282;
	{8'd66,8'd101} : s = 410;
	{8'd66,8'd102} : s = 131;
	{8'd66,8'd103} : s = 281;
	{8'd66,8'd104} : s = 278;
	{8'd66,8'd105} : s = 409;
	{8'd66,8'd106} : s = 277;
	{8'd66,8'd107} : s = 406;
	{8'd66,8'd108} : s = 405;
	{8'd66,8'd109} : s = 485;
	{8'd66,8'd110} : s = 112;
	{8'd66,8'd111} : s = 275;
	{8'd66,8'd112} : s = 270;
	{8'd66,8'd113} : s = 403;
	{8'd66,8'd114} : s = 269;
	{8'd66,8'd115} : s = 398;
	{8'd66,8'd116} : s = 397;
	{8'd66,8'd117} : s = 483;
	{8'd66,8'd118} : s = 267;
	{8'd66,8'd119} : s = 395;
	{8'd66,8'd120} : s = 391;
	{8'd66,8'd121} : s = 476;
	{8'd66,8'd122} : s = 376;
	{8'd66,8'd123} : s = 474;
	{8'd66,8'd124} : s = 473;
	{8'd66,8'd125} : s = 506;
	{8'd66,8'd126} : s = 20;
	{8'd66,8'd127} : s = 104;
	{8'd66,8'd128} : s = 100;
	{8'd66,8'd129} : s = 263;
	{8'd66,8'd130} : s = 98;
	{8'd66,8'd131} : s = 240;
	{8'd66,8'd132} : s = 232;
	{8'd66,8'd133} : s = 372;
	{8'd66,8'd134} : s = 97;
	{8'd66,8'd135} : s = 228;
	{8'd66,8'd136} : s = 226;
	{8'd66,8'd137} : s = 370;
	{8'd66,8'd138} : s = 225;
	{8'd66,8'd139} : s = 369;
	{8'd66,8'd140} : s = 364;
	{8'd66,8'd141} : s = 470;
	{8'd66,8'd142} : s = 88;
	{8'd66,8'd143} : s = 216;
	{8'd66,8'd144} : s = 212;
	{8'd66,8'd145} : s = 362;
	{8'd66,8'd146} : s = 210;
	{8'd66,8'd147} : s = 361;
	{8'd66,8'd148} : s = 358;
	{8'd66,8'd149} : s = 469;
	{8'd66,8'd150} : s = 209;
	{8'd66,8'd151} : s = 357;
	{8'd66,8'd152} : s = 355;
	{8'd66,8'd153} : s = 467;
	{8'd66,8'd154} : s = 348;
	{8'd66,8'd155} : s = 462;
	{8'd66,8'd156} : s = 461;
	{8'd66,8'd157} : s = 505;
	{8'd66,8'd158} : s = 84;
	{8'd66,8'd159} : s = 204;
	{8'd66,8'd160} : s = 202;
	{8'd66,8'd161} : s = 346;
	{8'd66,8'd162} : s = 201;
	{8'd66,8'd163} : s = 345;
	{8'd66,8'd164} : s = 342;
	{8'd66,8'd165} : s = 459;
	{8'd66,8'd166} : s = 198;
	{8'd66,8'd167} : s = 341;
	{8'd66,8'd168} : s = 339;
	{8'd66,8'd169} : s = 455;
	{8'd66,8'd170} : s = 334;
	{8'd66,8'd171} : s = 444;
	{8'd66,8'd172} : s = 442;
	{8'd66,8'd173} : s = 502;
	{8'd66,8'd174} : s = 197;
	{8'd66,8'd175} : s = 333;
	{8'd66,8'd176} : s = 331;
	{8'd66,8'd177} : s = 441;
	{8'd66,8'd178} : s = 327;
	{8'd66,8'd179} : s = 438;
	{8'd66,8'd180} : s = 437;
	{8'd66,8'd181} : s = 501;
	{8'd66,8'd182} : s = 316;
	{8'd66,8'd183} : s = 435;
	{8'd66,8'd184} : s = 430;
	{8'd66,8'd185} : s = 499;
	{8'd66,8'd186} : s = 429;
	{8'd66,8'd187} : s = 494;
	{8'd66,8'd188} : s = 493;
	{8'd66,8'd189} : s = 510;
	{8'd66,8'd190} : s = 1;
	{8'd66,8'd191} : s = 18;
	{8'd66,8'd192} : s = 17;
	{8'd66,8'd193} : s = 82;
	{8'd66,8'd194} : s = 12;
	{8'd66,8'd195} : s = 81;
	{8'd66,8'd196} : s = 76;
	{8'd66,8'd197} : s = 195;
	{8'd66,8'd198} : s = 10;
	{8'd66,8'd199} : s = 74;
	{8'd66,8'd200} : s = 73;
	{8'd66,8'd201} : s = 184;
	{8'd66,8'd202} : s = 70;
	{8'd66,8'd203} : s = 180;
	{8'd66,8'd204} : s = 178;
	{8'd66,8'd205} : s = 314;
	{8'd66,8'd206} : s = 9;
	{8'd66,8'd207} : s = 69;
	{8'd66,8'd208} : s = 67;
	{8'd66,8'd209} : s = 177;
	{8'd66,8'd210} : s = 56;
	{8'd66,8'd211} : s = 172;
	{8'd66,8'd212} : s = 170;
	{8'd66,8'd213} : s = 313;
	{8'd66,8'd214} : s = 52;
	{8'd66,8'd215} : s = 169;
	{8'd66,8'd216} : s = 166;
	{8'd66,8'd217} : s = 310;
	{8'd66,8'd218} : s = 165;
	{8'd66,8'd219} : s = 309;
	{8'd66,8'd220} : s = 307;
	{8'd66,8'd221} : s = 427;
	{8'd66,8'd222} : s = 6;
	{8'd66,8'd223} : s = 50;
	{8'd66,8'd224} : s = 49;
	{8'd66,8'd225} : s = 163;
	{8'd66,8'd226} : s = 44;
	{8'd66,8'd227} : s = 156;
	{8'd66,8'd228} : s = 154;
	{8'd66,8'd229} : s = 302;
	{8'd66,8'd230} : s = 42;
	{8'd66,8'd231} : s = 153;
	{8'd66,8'd232} : s = 150;
	{8'd66,8'd233} : s = 301;
	{8'd66,8'd234} : s = 149;
	{8'd66,8'd235} : s = 299;
	{8'd66,8'd236} : s = 295;
	{8'd66,8'd237} : s = 423;
	{8'd66,8'd238} : s = 41;
	{8'd66,8'd239} : s = 147;
	{8'd66,8'd240} : s = 142;
	{8'd66,8'd241} : s = 286;
	{8'd66,8'd242} : s = 141;
	{8'd66,8'd243} : s = 285;
	{8'd66,8'd244} : s = 283;
	{8'd66,8'd245} : s = 414;
	{8'd66,8'd246} : s = 139;
	{8'd66,8'd247} : s = 279;
	{8'd66,8'd248} : s = 271;
	{8'd66,8'd249} : s = 413;
	{8'd66,8'd250} : s = 248;
	{8'd66,8'd251} : s = 411;
	{8'd66,8'd252} : s = 407;
	{8'd66,8'd253} : s = 491;
	{8'd66,8'd254} : s = 5;
	{8'd66,8'd255} : s = 38;
	{8'd67,8'd0} : s = 274;
	{8'd67,8'd1} : s = 72;
	{8'd67,8'd2} : s = 273;
	{8'd67,8'd3} : s = 268;
	{8'd67,8'd4} : s = 396;
	{8'd67,8'd5} : s = 68;
	{8'd67,8'd6} : s = 266;
	{8'd67,8'd7} : s = 265;
	{8'd67,8'd8} : s = 394;
	{8'd67,8'd9} : s = 262;
	{8'd67,8'd10} : s = 393;
	{8'd67,8'd11} : s = 390;
	{8'd67,8'd12} : s = 468;
	{8'd67,8'd13} : s = 66;
	{8'd67,8'd14} : s = 261;
	{8'd67,8'd15} : s = 259;
	{8'd67,8'd16} : s = 389;
	{8'd67,8'd17} : s = 224;
	{8'd67,8'd18} : s = 387;
	{8'd67,8'd19} : s = 368;
	{8'd67,8'd20} : s = 466;
	{8'd67,8'd21} : s = 208;
	{8'd67,8'd22} : s = 360;
	{8'd67,8'd23} : s = 356;
	{8'd67,8'd24} : s = 465;
	{8'd67,8'd25} : s = 354;
	{8'd67,8'd26} : s = 460;
	{8'd67,8'd27} : s = 458;
	{8'd67,8'd28} : s = 500;
	{8'd67,8'd29} : s = 65;
	{8'd67,8'd30} : s = 200;
	{8'd67,8'd31} : s = 196;
	{8'd67,8'd32} : s = 353;
	{8'd67,8'd33} : s = 194;
	{8'd67,8'd34} : s = 344;
	{8'd67,8'd35} : s = 340;
	{8'd67,8'd36} : s = 457;
	{8'd67,8'd37} : s = 193;
	{8'd67,8'd38} : s = 338;
	{8'd67,8'd39} : s = 337;
	{8'd67,8'd40} : s = 454;
	{8'd67,8'd41} : s = 332;
	{8'd67,8'd42} : s = 453;
	{8'd67,8'd43} : s = 451;
	{8'd67,8'd44} : s = 498;
	{8'd67,8'd45} : s = 176;
	{8'd67,8'd46} : s = 330;
	{8'd67,8'd47} : s = 329;
	{8'd67,8'd48} : s = 440;
	{8'd67,8'd49} : s = 326;
	{8'd67,8'd50} : s = 436;
	{8'd67,8'd51} : s = 434;
	{8'd67,8'd52} : s = 497;
	{8'd67,8'd53} : s = 325;
	{8'd67,8'd54} : s = 433;
	{8'd67,8'd55} : s = 428;
	{8'd67,8'd56} : s = 492;
	{8'd67,8'd57} : s = 426;
	{8'd67,8'd58} : s = 490;
	{8'd67,8'd59} : s = 489;
	{8'd67,8'd60} : s = 508;
	{8'd67,8'd61} : s = 2;
	{8'd67,8'd62} : s = 48;
	{8'd67,8'd63} : s = 40;
	{8'd67,8'd64} : s = 168;
	{8'd67,8'd65} : s = 36;
	{8'd67,8'd66} : s = 164;
	{8'd67,8'd67} : s = 162;
	{8'd67,8'd68} : s = 323;
	{8'd67,8'd69} : s = 34;
	{8'd67,8'd70} : s = 161;
	{8'd67,8'd71} : s = 152;
	{8'd67,8'd72} : s = 312;
	{8'd67,8'd73} : s = 148;
	{8'd67,8'd74} : s = 308;
	{8'd67,8'd75} : s = 306;
	{8'd67,8'd76} : s = 425;
	{8'd67,8'd77} : s = 33;
	{8'd67,8'd78} : s = 146;
	{8'd67,8'd79} : s = 145;
	{8'd67,8'd80} : s = 305;
	{8'd67,8'd81} : s = 140;
	{8'd67,8'd82} : s = 300;
	{8'd67,8'd83} : s = 298;
	{8'd67,8'd84} : s = 422;
	{8'd67,8'd85} : s = 138;
	{8'd67,8'd86} : s = 297;
	{8'd67,8'd87} : s = 294;
	{8'd67,8'd88} : s = 421;
	{8'd67,8'd89} : s = 293;
	{8'd67,8'd90} : s = 419;
	{8'd67,8'd91} : s = 412;
	{8'd67,8'd92} : s = 486;
	{8'd67,8'd93} : s = 24;
	{8'd67,8'd94} : s = 137;
	{8'd67,8'd95} : s = 134;
	{8'd67,8'd96} : s = 291;
	{8'd67,8'd97} : s = 133;
	{8'd67,8'd98} : s = 284;
	{8'd67,8'd99} : s = 282;
	{8'd67,8'd100} : s = 410;
	{8'd67,8'd101} : s = 131;
	{8'd67,8'd102} : s = 281;
	{8'd67,8'd103} : s = 278;
	{8'd67,8'd104} : s = 409;
	{8'd67,8'd105} : s = 277;
	{8'd67,8'd106} : s = 406;
	{8'd67,8'd107} : s = 405;
	{8'd67,8'd108} : s = 485;
	{8'd67,8'd109} : s = 112;
	{8'd67,8'd110} : s = 275;
	{8'd67,8'd111} : s = 270;
	{8'd67,8'd112} : s = 403;
	{8'd67,8'd113} : s = 269;
	{8'd67,8'd114} : s = 398;
	{8'd67,8'd115} : s = 397;
	{8'd67,8'd116} : s = 483;
	{8'd67,8'd117} : s = 267;
	{8'd67,8'd118} : s = 395;
	{8'd67,8'd119} : s = 391;
	{8'd67,8'd120} : s = 476;
	{8'd67,8'd121} : s = 376;
	{8'd67,8'd122} : s = 474;
	{8'd67,8'd123} : s = 473;
	{8'd67,8'd124} : s = 506;
	{8'd67,8'd125} : s = 20;
	{8'd67,8'd126} : s = 104;
	{8'd67,8'd127} : s = 100;
	{8'd67,8'd128} : s = 263;
	{8'd67,8'd129} : s = 98;
	{8'd67,8'd130} : s = 240;
	{8'd67,8'd131} : s = 232;
	{8'd67,8'd132} : s = 372;
	{8'd67,8'd133} : s = 97;
	{8'd67,8'd134} : s = 228;
	{8'd67,8'd135} : s = 226;
	{8'd67,8'd136} : s = 370;
	{8'd67,8'd137} : s = 225;
	{8'd67,8'd138} : s = 369;
	{8'd67,8'd139} : s = 364;
	{8'd67,8'd140} : s = 470;
	{8'd67,8'd141} : s = 88;
	{8'd67,8'd142} : s = 216;
	{8'd67,8'd143} : s = 212;
	{8'd67,8'd144} : s = 362;
	{8'd67,8'd145} : s = 210;
	{8'd67,8'd146} : s = 361;
	{8'd67,8'd147} : s = 358;
	{8'd67,8'd148} : s = 469;
	{8'd67,8'd149} : s = 209;
	{8'd67,8'd150} : s = 357;
	{8'd67,8'd151} : s = 355;
	{8'd67,8'd152} : s = 467;
	{8'd67,8'd153} : s = 348;
	{8'd67,8'd154} : s = 462;
	{8'd67,8'd155} : s = 461;
	{8'd67,8'd156} : s = 505;
	{8'd67,8'd157} : s = 84;
	{8'd67,8'd158} : s = 204;
	{8'd67,8'd159} : s = 202;
	{8'd67,8'd160} : s = 346;
	{8'd67,8'd161} : s = 201;
	{8'd67,8'd162} : s = 345;
	{8'd67,8'd163} : s = 342;
	{8'd67,8'd164} : s = 459;
	{8'd67,8'd165} : s = 198;
	{8'd67,8'd166} : s = 341;
	{8'd67,8'd167} : s = 339;
	{8'd67,8'd168} : s = 455;
	{8'd67,8'd169} : s = 334;
	{8'd67,8'd170} : s = 444;
	{8'd67,8'd171} : s = 442;
	{8'd67,8'd172} : s = 502;
	{8'd67,8'd173} : s = 197;
	{8'd67,8'd174} : s = 333;
	{8'd67,8'd175} : s = 331;
	{8'd67,8'd176} : s = 441;
	{8'd67,8'd177} : s = 327;
	{8'd67,8'd178} : s = 438;
	{8'd67,8'd179} : s = 437;
	{8'd67,8'd180} : s = 501;
	{8'd67,8'd181} : s = 316;
	{8'd67,8'd182} : s = 435;
	{8'd67,8'd183} : s = 430;
	{8'd67,8'd184} : s = 499;
	{8'd67,8'd185} : s = 429;
	{8'd67,8'd186} : s = 494;
	{8'd67,8'd187} : s = 493;
	{8'd67,8'd188} : s = 510;
	{8'd67,8'd189} : s = 1;
	{8'd67,8'd190} : s = 18;
	{8'd67,8'd191} : s = 17;
	{8'd67,8'd192} : s = 82;
	{8'd67,8'd193} : s = 12;
	{8'd67,8'd194} : s = 81;
	{8'd67,8'd195} : s = 76;
	{8'd67,8'd196} : s = 195;
	{8'd67,8'd197} : s = 10;
	{8'd67,8'd198} : s = 74;
	{8'd67,8'd199} : s = 73;
	{8'd67,8'd200} : s = 184;
	{8'd67,8'd201} : s = 70;
	{8'd67,8'd202} : s = 180;
	{8'd67,8'd203} : s = 178;
	{8'd67,8'd204} : s = 314;
	{8'd67,8'd205} : s = 9;
	{8'd67,8'd206} : s = 69;
	{8'd67,8'd207} : s = 67;
	{8'd67,8'd208} : s = 177;
	{8'd67,8'd209} : s = 56;
	{8'd67,8'd210} : s = 172;
	{8'd67,8'd211} : s = 170;
	{8'd67,8'd212} : s = 313;
	{8'd67,8'd213} : s = 52;
	{8'd67,8'd214} : s = 169;
	{8'd67,8'd215} : s = 166;
	{8'd67,8'd216} : s = 310;
	{8'd67,8'd217} : s = 165;
	{8'd67,8'd218} : s = 309;
	{8'd67,8'd219} : s = 307;
	{8'd67,8'd220} : s = 427;
	{8'd67,8'd221} : s = 6;
	{8'd67,8'd222} : s = 50;
	{8'd67,8'd223} : s = 49;
	{8'd67,8'd224} : s = 163;
	{8'd67,8'd225} : s = 44;
	{8'd67,8'd226} : s = 156;
	{8'd67,8'd227} : s = 154;
	{8'd67,8'd228} : s = 302;
	{8'd67,8'd229} : s = 42;
	{8'd67,8'd230} : s = 153;
	{8'd67,8'd231} : s = 150;
	{8'd67,8'd232} : s = 301;
	{8'd67,8'd233} : s = 149;
	{8'd67,8'd234} : s = 299;
	{8'd67,8'd235} : s = 295;
	{8'd67,8'd236} : s = 423;
	{8'd67,8'd237} : s = 41;
	{8'd67,8'd238} : s = 147;
	{8'd67,8'd239} : s = 142;
	{8'd67,8'd240} : s = 286;
	{8'd67,8'd241} : s = 141;
	{8'd67,8'd242} : s = 285;
	{8'd67,8'd243} : s = 283;
	{8'd67,8'd244} : s = 414;
	{8'd67,8'd245} : s = 139;
	{8'd67,8'd246} : s = 279;
	{8'd67,8'd247} : s = 271;
	{8'd67,8'd248} : s = 413;
	{8'd67,8'd249} : s = 248;
	{8'd67,8'd250} : s = 411;
	{8'd67,8'd251} : s = 407;
	{8'd67,8'd252} : s = 491;
	{8'd67,8'd253} : s = 5;
	{8'd67,8'd254} : s = 38;
	{8'd67,8'd255} : s = 37;
	{8'd68,8'd0} : s = 72;
	{8'd68,8'd1} : s = 273;
	{8'd68,8'd2} : s = 268;
	{8'd68,8'd3} : s = 396;
	{8'd68,8'd4} : s = 68;
	{8'd68,8'd5} : s = 266;
	{8'd68,8'd6} : s = 265;
	{8'd68,8'd7} : s = 394;
	{8'd68,8'd8} : s = 262;
	{8'd68,8'd9} : s = 393;
	{8'd68,8'd10} : s = 390;
	{8'd68,8'd11} : s = 468;
	{8'd68,8'd12} : s = 66;
	{8'd68,8'd13} : s = 261;
	{8'd68,8'd14} : s = 259;
	{8'd68,8'd15} : s = 389;
	{8'd68,8'd16} : s = 224;
	{8'd68,8'd17} : s = 387;
	{8'd68,8'd18} : s = 368;
	{8'd68,8'd19} : s = 466;
	{8'd68,8'd20} : s = 208;
	{8'd68,8'd21} : s = 360;
	{8'd68,8'd22} : s = 356;
	{8'd68,8'd23} : s = 465;
	{8'd68,8'd24} : s = 354;
	{8'd68,8'd25} : s = 460;
	{8'd68,8'd26} : s = 458;
	{8'd68,8'd27} : s = 500;
	{8'd68,8'd28} : s = 65;
	{8'd68,8'd29} : s = 200;
	{8'd68,8'd30} : s = 196;
	{8'd68,8'd31} : s = 353;
	{8'd68,8'd32} : s = 194;
	{8'd68,8'd33} : s = 344;
	{8'd68,8'd34} : s = 340;
	{8'd68,8'd35} : s = 457;
	{8'd68,8'd36} : s = 193;
	{8'd68,8'd37} : s = 338;
	{8'd68,8'd38} : s = 337;
	{8'd68,8'd39} : s = 454;
	{8'd68,8'd40} : s = 332;
	{8'd68,8'd41} : s = 453;
	{8'd68,8'd42} : s = 451;
	{8'd68,8'd43} : s = 498;
	{8'd68,8'd44} : s = 176;
	{8'd68,8'd45} : s = 330;
	{8'd68,8'd46} : s = 329;
	{8'd68,8'd47} : s = 440;
	{8'd68,8'd48} : s = 326;
	{8'd68,8'd49} : s = 436;
	{8'd68,8'd50} : s = 434;
	{8'd68,8'd51} : s = 497;
	{8'd68,8'd52} : s = 325;
	{8'd68,8'd53} : s = 433;
	{8'd68,8'd54} : s = 428;
	{8'd68,8'd55} : s = 492;
	{8'd68,8'd56} : s = 426;
	{8'd68,8'd57} : s = 490;
	{8'd68,8'd58} : s = 489;
	{8'd68,8'd59} : s = 508;
	{8'd68,8'd60} : s = 2;
	{8'd68,8'd61} : s = 48;
	{8'd68,8'd62} : s = 40;
	{8'd68,8'd63} : s = 168;
	{8'd68,8'd64} : s = 36;
	{8'd68,8'd65} : s = 164;
	{8'd68,8'd66} : s = 162;
	{8'd68,8'd67} : s = 323;
	{8'd68,8'd68} : s = 34;
	{8'd68,8'd69} : s = 161;
	{8'd68,8'd70} : s = 152;
	{8'd68,8'd71} : s = 312;
	{8'd68,8'd72} : s = 148;
	{8'd68,8'd73} : s = 308;
	{8'd68,8'd74} : s = 306;
	{8'd68,8'd75} : s = 425;
	{8'd68,8'd76} : s = 33;
	{8'd68,8'd77} : s = 146;
	{8'd68,8'd78} : s = 145;
	{8'd68,8'd79} : s = 305;
	{8'd68,8'd80} : s = 140;
	{8'd68,8'd81} : s = 300;
	{8'd68,8'd82} : s = 298;
	{8'd68,8'd83} : s = 422;
	{8'd68,8'd84} : s = 138;
	{8'd68,8'd85} : s = 297;
	{8'd68,8'd86} : s = 294;
	{8'd68,8'd87} : s = 421;
	{8'd68,8'd88} : s = 293;
	{8'd68,8'd89} : s = 419;
	{8'd68,8'd90} : s = 412;
	{8'd68,8'd91} : s = 486;
	{8'd68,8'd92} : s = 24;
	{8'd68,8'd93} : s = 137;
	{8'd68,8'd94} : s = 134;
	{8'd68,8'd95} : s = 291;
	{8'd68,8'd96} : s = 133;
	{8'd68,8'd97} : s = 284;
	{8'd68,8'd98} : s = 282;
	{8'd68,8'd99} : s = 410;
	{8'd68,8'd100} : s = 131;
	{8'd68,8'd101} : s = 281;
	{8'd68,8'd102} : s = 278;
	{8'd68,8'd103} : s = 409;
	{8'd68,8'd104} : s = 277;
	{8'd68,8'd105} : s = 406;
	{8'd68,8'd106} : s = 405;
	{8'd68,8'd107} : s = 485;
	{8'd68,8'd108} : s = 112;
	{8'd68,8'd109} : s = 275;
	{8'd68,8'd110} : s = 270;
	{8'd68,8'd111} : s = 403;
	{8'd68,8'd112} : s = 269;
	{8'd68,8'd113} : s = 398;
	{8'd68,8'd114} : s = 397;
	{8'd68,8'd115} : s = 483;
	{8'd68,8'd116} : s = 267;
	{8'd68,8'd117} : s = 395;
	{8'd68,8'd118} : s = 391;
	{8'd68,8'd119} : s = 476;
	{8'd68,8'd120} : s = 376;
	{8'd68,8'd121} : s = 474;
	{8'd68,8'd122} : s = 473;
	{8'd68,8'd123} : s = 506;
	{8'd68,8'd124} : s = 20;
	{8'd68,8'd125} : s = 104;
	{8'd68,8'd126} : s = 100;
	{8'd68,8'd127} : s = 263;
	{8'd68,8'd128} : s = 98;
	{8'd68,8'd129} : s = 240;
	{8'd68,8'd130} : s = 232;
	{8'd68,8'd131} : s = 372;
	{8'd68,8'd132} : s = 97;
	{8'd68,8'd133} : s = 228;
	{8'd68,8'd134} : s = 226;
	{8'd68,8'd135} : s = 370;
	{8'd68,8'd136} : s = 225;
	{8'd68,8'd137} : s = 369;
	{8'd68,8'd138} : s = 364;
	{8'd68,8'd139} : s = 470;
	{8'd68,8'd140} : s = 88;
	{8'd68,8'd141} : s = 216;
	{8'd68,8'd142} : s = 212;
	{8'd68,8'd143} : s = 362;
	{8'd68,8'd144} : s = 210;
	{8'd68,8'd145} : s = 361;
	{8'd68,8'd146} : s = 358;
	{8'd68,8'd147} : s = 469;
	{8'd68,8'd148} : s = 209;
	{8'd68,8'd149} : s = 357;
	{8'd68,8'd150} : s = 355;
	{8'd68,8'd151} : s = 467;
	{8'd68,8'd152} : s = 348;
	{8'd68,8'd153} : s = 462;
	{8'd68,8'd154} : s = 461;
	{8'd68,8'd155} : s = 505;
	{8'd68,8'd156} : s = 84;
	{8'd68,8'd157} : s = 204;
	{8'd68,8'd158} : s = 202;
	{8'd68,8'd159} : s = 346;
	{8'd68,8'd160} : s = 201;
	{8'd68,8'd161} : s = 345;
	{8'd68,8'd162} : s = 342;
	{8'd68,8'd163} : s = 459;
	{8'd68,8'd164} : s = 198;
	{8'd68,8'd165} : s = 341;
	{8'd68,8'd166} : s = 339;
	{8'd68,8'd167} : s = 455;
	{8'd68,8'd168} : s = 334;
	{8'd68,8'd169} : s = 444;
	{8'd68,8'd170} : s = 442;
	{8'd68,8'd171} : s = 502;
	{8'd68,8'd172} : s = 197;
	{8'd68,8'd173} : s = 333;
	{8'd68,8'd174} : s = 331;
	{8'd68,8'd175} : s = 441;
	{8'd68,8'd176} : s = 327;
	{8'd68,8'd177} : s = 438;
	{8'd68,8'd178} : s = 437;
	{8'd68,8'd179} : s = 501;
	{8'd68,8'd180} : s = 316;
	{8'd68,8'd181} : s = 435;
	{8'd68,8'd182} : s = 430;
	{8'd68,8'd183} : s = 499;
	{8'd68,8'd184} : s = 429;
	{8'd68,8'd185} : s = 494;
	{8'd68,8'd186} : s = 493;
	{8'd68,8'd187} : s = 510;
	{8'd68,8'd188} : s = 1;
	{8'd68,8'd189} : s = 18;
	{8'd68,8'd190} : s = 17;
	{8'd68,8'd191} : s = 82;
	{8'd68,8'd192} : s = 12;
	{8'd68,8'd193} : s = 81;
	{8'd68,8'd194} : s = 76;
	{8'd68,8'd195} : s = 195;
	{8'd68,8'd196} : s = 10;
	{8'd68,8'd197} : s = 74;
	{8'd68,8'd198} : s = 73;
	{8'd68,8'd199} : s = 184;
	{8'd68,8'd200} : s = 70;
	{8'd68,8'd201} : s = 180;
	{8'd68,8'd202} : s = 178;
	{8'd68,8'd203} : s = 314;
	{8'd68,8'd204} : s = 9;
	{8'd68,8'd205} : s = 69;
	{8'd68,8'd206} : s = 67;
	{8'd68,8'd207} : s = 177;
	{8'd68,8'd208} : s = 56;
	{8'd68,8'd209} : s = 172;
	{8'd68,8'd210} : s = 170;
	{8'd68,8'd211} : s = 313;
	{8'd68,8'd212} : s = 52;
	{8'd68,8'd213} : s = 169;
	{8'd68,8'd214} : s = 166;
	{8'd68,8'd215} : s = 310;
	{8'd68,8'd216} : s = 165;
	{8'd68,8'd217} : s = 309;
	{8'd68,8'd218} : s = 307;
	{8'd68,8'd219} : s = 427;
	{8'd68,8'd220} : s = 6;
	{8'd68,8'd221} : s = 50;
	{8'd68,8'd222} : s = 49;
	{8'd68,8'd223} : s = 163;
	{8'd68,8'd224} : s = 44;
	{8'd68,8'd225} : s = 156;
	{8'd68,8'd226} : s = 154;
	{8'd68,8'd227} : s = 302;
	{8'd68,8'd228} : s = 42;
	{8'd68,8'd229} : s = 153;
	{8'd68,8'd230} : s = 150;
	{8'd68,8'd231} : s = 301;
	{8'd68,8'd232} : s = 149;
	{8'd68,8'd233} : s = 299;
	{8'd68,8'd234} : s = 295;
	{8'd68,8'd235} : s = 423;
	{8'd68,8'd236} : s = 41;
	{8'd68,8'd237} : s = 147;
	{8'd68,8'd238} : s = 142;
	{8'd68,8'd239} : s = 286;
	{8'd68,8'd240} : s = 141;
	{8'd68,8'd241} : s = 285;
	{8'd68,8'd242} : s = 283;
	{8'd68,8'd243} : s = 414;
	{8'd68,8'd244} : s = 139;
	{8'd68,8'd245} : s = 279;
	{8'd68,8'd246} : s = 271;
	{8'd68,8'd247} : s = 413;
	{8'd68,8'd248} : s = 248;
	{8'd68,8'd249} : s = 411;
	{8'd68,8'd250} : s = 407;
	{8'd68,8'd251} : s = 491;
	{8'd68,8'd252} : s = 5;
	{8'd68,8'd253} : s = 38;
	{8'd68,8'd254} : s = 37;
	{8'd68,8'd255} : s = 135;
	{8'd69,8'd0} : s = 273;
	{8'd69,8'd1} : s = 268;
	{8'd69,8'd2} : s = 396;
	{8'd69,8'd3} : s = 68;
	{8'd69,8'd4} : s = 266;
	{8'd69,8'd5} : s = 265;
	{8'd69,8'd6} : s = 394;
	{8'd69,8'd7} : s = 262;
	{8'd69,8'd8} : s = 393;
	{8'd69,8'd9} : s = 390;
	{8'd69,8'd10} : s = 468;
	{8'd69,8'd11} : s = 66;
	{8'd69,8'd12} : s = 261;
	{8'd69,8'd13} : s = 259;
	{8'd69,8'd14} : s = 389;
	{8'd69,8'd15} : s = 224;
	{8'd69,8'd16} : s = 387;
	{8'd69,8'd17} : s = 368;
	{8'd69,8'd18} : s = 466;
	{8'd69,8'd19} : s = 208;
	{8'd69,8'd20} : s = 360;
	{8'd69,8'd21} : s = 356;
	{8'd69,8'd22} : s = 465;
	{8'd69,8'd23} : s = 354;
	{8'd69,8'd24} : s = 460;
	{8'd69,8'd25} : s = 458;
	{8'd69,8'd26} : s = 500;
	{8'd69,8'd27} : s = 65;
	{8'd69,8'd28} : s = 200;
	{8'd69,8'd29} : s = 196;
	{8'd69,8'd30} : s = 353;
	{8'd69,8'd31} : s = 194;
	{8'd69,8'd32} : s = 344;
	{8'd69,8'd33} : s = 340;
	{8'd69,8'd34} : s = 457;
	{8'd69,8'd35} : s = 193;
	{8'd69,8'd36} : s = 338;
	{8'd69,8'd37} : s = 337;
	{8'd69,8'd38} : s = 454;
	{8'd69,8'd39} : s = 332;
	{8'd69,8'd40} : s = 453;
	{8'd69,8'd41} : s = 451;
	{8'd69,8'd42} : s = 498;
	{8'd69,8'd43} : s = 176;
	{8'd69,8'd44} : s = 330;
	{8'd69,8'd45} : s = 329;
	{8'd69,8'd46} : s = 440;
	{8'd69,8'd47} : s = 326;
	{8'd69,8'd48} : s = 436;
	{8'd69,8'd49} : s = 434;
	{8'd69,8'd50} : s = 497;
	{8'd69,8'd51} : s = 325;
	{8'd69,8'd52} : s = 433;
	{8'd69,8'd53} : s = 428;
	{8'd69,8'd54} : s = 492;
	{8'd69,8'd55} : s = 426;
	{8'd69,8'd56} : s = 490;
	{8'd69,8'd57} : s = 489;
	{8'd69,8'd58} : s = 508;
	{8'd69,8'd59} : s = 2;
	{8'd69,8'd60} : s = 48;
	{8'd69,8'd61} : s = 40;
	{8'd69,8'd62} : s = 168;
	{8'd69,8'd63} : s = 36;
	{8'd69,8'd64} : s = 164;
	{8'd69,8'd65} : s = 162;
	{8'd69,8'd66} : s = 323;
	{8'd69,8'd67} : s = 34;
	{8'd69,8'd68} : s = 161;
	{8'd69,8'd69} : s = 152;
	{8'd69,8'd70} : s = 312;
	{8'd69,8'd71} : s = 148;
	{8'd69,8'd72} : s = 308;
	{8'd69,8'd73} : s = 306;
	{8'd69,8'd74} : s = 425;
	{8'd69,8'd75} : s = 33;
	{8'd69,8'd76} : s = 146;
	{8'd69,8'd77} : s = 145;
	{8'd69,8'd78} : s = 305;
	{8'd69,8'd79} : s = 140;
	{8'd69,8'd80} : s = 300;
	{8'd69,8'd81} : s = 298;
	{8'd69,8'd82} : s = 422;
	{8'd69,8'd83} : s = 138;
	{8'd69,8'd84} : s = 297;
	{8'd69,8'd85} : s = 294;
	{8'd69,8'd86} : s = 421;
	{8'd69,8'd87} : s = 293;
	{8'd69,8'd88} : s = 419;
	{8'd69,8'd89} : s = 412;
	{8'd69,8'd90} : s = 486;
	{8'd69,8'd91} : s = 24;
	{8'd69,8'd92} : s = 137;
	{8'd69,8'd93} : s = 134;
	{8'd69,8'd94} : s = 291;
	{8'd69,8'd95} : s = 133;
	{8'd69,8'd96} : s = 284;
	{8'd69,8'd97} : s = 282;
	{8'd69,8'd98} : s = 410;
	{8'd69,8'd99} : s = 131;
	{8'd69,8'd100} : s = 281;
	{8'd69,8'd101} : s = 278;
	{8'd69,8'd102} : s = 409;
	{8'd69,8'd103} : s = 277;
	{8'd69,8'd104} : s = 406;
	{8'd69,8'd105} : s = 405;
	{8'd69,8'd106} : s = 485;
	{8'd69,8'd107} : s = 112;
	{8'd69,8'd108} : s = 275;
	{8'd69,8'd109} : s = 270;
	{8'd69,8'd110} : s = 403;
	{8'd69,8'd111} : s = 269;
	{8'd69,8'd112} : s = 398;
	{8'd69,8'd113} : s = 397;
	{8'd69,8'd114} : s = 483;
	{8'd69,8'd115} : s = 267;
	{8'd69,8'd116} : s = 395;
	{8'd69,8'd117} : s = 391;
	{8'd69,8'd118} : s = 476;
	{8'd69,8'd119} : s = 376;
	{8'd69,8'd120} : s = 474;
	{8'd69,8'd121} : s = 473;
	{8'd69,8'd122} : s = 506;
	{8'd69,8'd123} : s = 20;
	{8'd69,8'd124} : s = 104;
	{8'd69,8'd125} : s = 100;
	{8'd69,8'd126} : s = 263;
	{8'd69,8'd127} : s = 98;
	{8'd69,8'd128} : s = 240;
	{8'd69,8'd129} : s = 232;
	{8'd69,8'd130} : s = 372;
	{8'd69,8'd131} : s = 97;
	{8'd69,8'd132} : s = 228;
	{8'd69,8'd133} : s = 226;
	{8'd69,8'd134} : s = 370;
	{8'd69,8'd135} : s = 225;
	{8'd69,8'd136} : s = 369;
	{8'd69,8'd137} : s = 364;
	{8'd69,8'd138} : s = 470;
	{8'd69,8'd139} : s = 88;
	{8'd69,8'd140} : s = 216;
	{8'd69,8'd141} : s = 212;
	{8'd69,8'd142} : s = 362;
	{8'd69,8'd143} : s = 210;
	{8'd69,8'd144} : s = 361;
	{8'd69,8'd145} : s = 358;
	{8'd69,8'd146} : s = 469;
	{8'd69,8'd147} : s = 209;
	{8'd69,8'd148} : s = 357;
	{8'd69,8'd149} : s = 355;
	{8'd69,8'd150} : s = 467;
	{8'd69,8'd151} : s = 348;
	{8'd69,8'd152} : s = 462;
	{8'd69,8'd153} : s = 461;
	{8'd69,8'd154} : s = 505;
	{8'd69,8'd155} : s = 84;
	{8'd69,8'd156} : s = 204;
	{8'd69,8'd157} : s = 202;
	{8'd69,8'd158} : s = 346;
	{8'd69,8'd159} : s = 201;
	{8'd69,8'd160} : s = 345;
	{8'd69,8'd161} : s = 342;
	{8'd69,8'd162} : s = 459;
	{8'd69,8'd163} : s = 198;
	{8'd69,8'd164} : s = 341;
	{8'd69,8'd165} : s = 339;
	{8'd69,8'd166} : s = 455;
	{8'd69,8'd167} : s = 334;
	{8'd69,8'd168} : s = 444;
	{8'd69,8'd169} : s = 442;
	{8'd69,8'd170} : s = 502;
	{8'd69,8'd171} : s = 197;
	{8'd69,8'd172} : s = 333;
	{8'd69,8'd173} : s = 331;
	{8'd69,8'd174} : s = 441;
	{8'd69,8'd175} : s = 327;
	{8'd69,8'd176} : s = 438;
	{8'd69,8'd177} : s = 437;
	{8'd69,8'd178} : s = 501;
	{8'd69,8'd179} : s = 316;
	{8'd69,8'd180} : s = 435;
	{8'd69,8'd181} : s = 430;
	{8'd69,8'd182} : s = 499;
	{8'd69,8'd183} : s = 429;
	{8'd69,8'd184} : s = 494;
	{8'd69,8'd185} : s = 493;
	{8'd69,8'd186} : s = 510;
	{8'd69,8'd187} : s = 1;
	{8'd69,8'd188} : s = 18;
	{8'd69,8'd189} : s = 17;
	{8'd69,8'd190} : s = 82;
	{8'd69,8'd191} : s = 12;
	{8'd69,8'd192} : s = 81;
	{8'd69,8'd193} : s = 76;
	{8'd69,8'd194} : s = 195;
	{8'd69,8'd195} : s = 10;
	{8'd69,8'd196} : s = 74;
	{8'd69,8'd197} : s = 73;
	{8'd69,8'd198} : s = 184;
	{8'd69,8'd199} : s = 70;
	{8'd69,8'd200} : s = 180;
	{8'd69,8'd201} : s = 178;
	{8'd69,8'd202} : s = 314;
	{8'd69,8'd203} : s = 9;
	{8'd69,8'd204} : s = 69;
	{8'd69,8'd205} : s = 67;
	{8'd69,8'd206} : s = 177;
	{8'd69,8'd207} : s = 56;
	{8'd69,8'd208} : s = 172;
	{8'd69,8'd209} : s = 170;
	{8'd69,8'd210} : s = 313;
	{8'd69,8'd211} : s = 52;
	{8'd69,8'd212} : s = 169;
	{8'd69,8'd213} : s = 166;
	{8'd69,8'd214} : s = 310;
	{8'd69,8'd215} : s = 165;
	{8'd69,8'd216} : s = 309;
	{8'd69,8'd217} : s = 307;
	{8'd69,8'd218} : s = 427;
	{8'd69,8'd219} : s = 6;
	{8'd69,8'd220} : s = 50;
	{8'd69,8'd221} : s = 49;
	{8'd69,8'd222} : s = 163;
	{8'd69,8'd223} : s = 44;
	{8'd69,8'd224} : s = 156;
	{8'd69,8'd225} : s = 154;
	{8'd69,8'd226} : s = 302;
	{8'd69,8'd227} : s = 42;
	{8'd69,8'd228} : s = 153;
	{8'd69,8'd229} : s = 150;
	{8'd69,8'd230} : s = 301;
	{8'd69,8'd231} : s = 149;
	{8'd69,8'd232} : s = 299;
	{8'd69,8'd233} : s = 295;
	{8'd69,8'd234} : s = 423;
	{8'd69,8'd235} : s = 41;
	{8'd69,8'd236} : s = 147;
	{8'd69,8'd237} : s = 142;
	{8'd69,8'd238} : s = 286;
	{8'd69,8'd239} : s = 141;
	{8'd69,8'd240} : s = 285;
	{8'd69,8'd241} : s = 283;
	{8'd69,8'd242} : s = 414;
	{8'd69,8'd243} : s = 139;
	{8'd69,8'd244} : s = 279;
	{8'd69,8'd245} : s = 271;
	{8'd69,8'd246} : s = 413;
	{8'd69,8'd247} : s = 248;
	{8'd69,8'd248} : s = 411;
	{8'd69,8'd249} : s = 407;
	{8'd69,8'd250} : s = 491;
	{8'd69,8'd251} : s = 5;
	{8'd69,8'd252} : s = 38;
	{8'd69,8'd253} : s = 37;
	{8'd69,8'd254} : s = 135;
	{8'd69,8'd255} : s = 35;
	{8'd70,8'd0} : s = 268;
	{8'd70,8'd1} : s = 396;
	{8'd70,8'd2} : s = 68;
	{8'd70,8'd3} : s = 266;
	{8'd70,8'd4} : s = 265;
	{8'd70,8'd5} : s = 394;
	{8'd70,8'd6} : s = 262;
	{8'd70,8'd7} : s = 393;
	{8'd70,8'd8} : s = 390;
	{8'd70,8'd9} : s = 468;
	{8'd70,8'd10} : s = 66;
	{8'd70,8'd11} : s = 261;
	{8'd70,8'd12} : s = 259;
	{8'd70,8'd13} : s = 389;
	{8'd70,8'd14} : s = 224;
	{8'd70,8'd15} : s = 387;
	{8'd70,8'd16} : s = 368;
	{8'd70,8'd17} : s = 466;
	{8'd70,8'd18} : s = 208;
	{8'd70,8'd19} : s = 360;
	{8'd70,8'd20} : s = 356;
	{8'd70,8'd21} : s = 465;
	{8'd70,8'd22} : s = 354;
	{8'd70,8'd23} : s = 460;
	{8'd70,8'd24} : s = 458;
	{8'd70,8'd25} : s = 500;
	{8'd70,8'd26} : s = 65;
	{8'd70,8'd27} : s = 200;
	{8'd70,8'd28} : s = 196;
	{8'd70,8'd29} : s = 353;
	{8'd70,8'd30} : s = 194;
	{8'd70,8'd31} : s = 344;
	{8'd70,8'd32} : s = 340;
	{8'd70,8'd33} : s = 457;
	{8'd70,8'd34} : s = 193;
	{8'd70,8'd35} : s = 338;
	{8'd70,8'd36} : s = 337;
	{8'd70,8'd37} : s = 454;
	{8'd70,8'd38} : s = 332;
	{8'd70,8'd39} : s = 453;
	{8'd70,8'd40} : s = 451;
	{8'd70,8'd41} : s = 498;
	{8'd70,8'd42} : s = 176;
	{8'd70,8'd43} : s = 330;
	{8'd70,8'd44} : s = 329;
	{8'd70,8'd45} : s = 440;
	{8'd70,8'd46} : s = 326;
	{8'd70,8'd47} : s = 436;
	{8'd70,8'd48} : s = 434;
	{8'd70,8'd49} : s = 497;
	{8'd70,8'd50} : s = 325;
	{8'd70,8'd51} : s = 433;
	{8'd70,8'd52} : s = 428;
	{8'd70,8'd53} : s = 492;
	{8'd70,8'd54} : s = 426;
	{8'd70,8'd55} : s = 490;
	{8'd70,8'd56} : s = 489;
	{8'd70,8'd57} : s = 508;
	{8'd70,8'd58} : s = 2;
	{8'd70,8'd59} : s = 48;
	{8'd70,8'd60} : s = 40;
	{8'd70,8'd61} : s = 168;
	{8'd70,8'd62} : s = 36;
	{8'd70,8'd63} : s = 164;
	{8'd70,8'd64} : s = 162;
	{8'd70,8'd65} : s = 323;
	{8'd70,8'd66} : s = 34;
	{8'd70,8'd67} : s = 161;
	{8'd70,8'd68} : s = 152;
	{8'd70,8'd69} : s = 312;
	{8'd70,8'd70} : s = 148;
	{8'd70,8'd71} : s = 308;
	{8'd70,8'd72} : s = 306;
	{8'd70,8'd73} : s = 425;
	{8'd70,8'd74} : s = 33;
	{8'd70,8'd75} : s = 146;
	{8'd70,8'd76} : s = 145;
	{8'd70,8'd77} : s = 305;
	{8'd70,8'd78} : s = 140;
	{8'd70,8'd79} : s = 300;
	{8'd70,8'd80} : s = 298;
	{8'd70,8'd81} : s = 422;
	{8'd70,8'd82} : s = 138;
	{8'd70,8'd83} : s = 297;
	{8'd70,8'd84} : s = 294;
	{8'd70,8'd85} : s = 421;
	{8'd70,8'd86} : s = 293;
	{8'd70,8'd87} : s = 419;
	{8'd70,8'd88} : s = 412;
	{8'd70,8'd89} : s = 486;
	{8'd70,8'd90} : s = 24;
	{8'd70,8'd91} : s = 137;
	{8'd70,8'd92} : s = 134;
	{8'd70,8'd93} : s = 291;
	{8'd70,8'd94} : s = 133;
	{8'd70,8'd95} : s = 284;
	{8'd70,8'd96} : s = 282;
	{8'd70,8'd97} : s = 410;
	{8'd70,8'd98} : s = 131;
	{8'd70,8'd99} : s = 281;
	{8'd70,8'd100} : s = 278;
	{8'd70,8'd101} : s = 409;
	{8'd70,8'd102} : s = 277;
	{8'd70,8'd103} : s = 406;
	{8'd70,8'd104} : s = 405;
	{8'd70,8'd105} : s = 485;
	{8'd70,8'd106} : s = 112;
	{8'd70,8'd107} : s = 275;
	{8'd70,8'd108} : s = 270;
	{8'd70,8'd109} : s = 403;
	{8'd70,8'd110} : s = 269;
	{8'd70,8'd111} : s = 398;
	{8'd70,8'd112} : s = 397;
	{8'd70,8'd113} : s = 483;
	{8'd70,8'd114} : s = 267;
	{8'd70,8'd115} : s = 395;
	{8'd70,8'd116} : s = 391;
	{8'd70,8'd117} : s = 476;
	{8'd70,8'd118} : s = 376;
	{8'd70,8'd119} : s = 474;
	{8'd70,8'd120} : s = 473;
	{8'd70,8'd121} : s = 506;
	{8'd70,8'd122} : s = 20;
	{8'd70,8'd123} : s = 104;
	{8'd70,8'd124} : s = 100;
	{8'd70,8'd125} : s = 263;
	{8'd70,8'd126} : s = 98;
	{8'd70,8'd127} : s = 240;
	{8'd70,8'd128} : s = 232;
	{8'd70,8'd129} : s = 372;
	{8'd70,8'd130} : s = 97;
	{8'd70,8'd131} : s = 228;
	{8'd70,8'd132} : s = 226;
	{8'd70,8'd133} : s = 370;
	{8'd70,8'd134} : s = 225;
	{8'd70,8'd135} : s = 369;
	{8'd70,8'd136} : s = 364;
	{8'd70,8'd137} : s = 470;
	{8'd70,8'd138} : s = 88;
	{8'd70,8'd139} : s = 216;
	{8'd70,8'd140} : s = 212;
	{8'd70,8'd141} : s = 362;
	{8'd70,8'd142} : s = 210;
	{8'd70,8'd143} : s = 361;
	{8'd70,8'd144} : s = 358;
	{8'd70,8'd145} : s = 469;
	{8'd70,8'd146} : s = 209;
	{8'd70,8'd147} : s = 357;
	{8'd70,8'd148} : s = 355;
	{8'd70,8'd149} : s = 467;
	{8'd70,8'd150} : s = 348;
	{8'd70,8'd151} : s = 462;
	{8'd70,8'd152} : s = 461;
	{8'd70,8'd153} : s = 505;
	{8'd70,8'd154} : s = 84;
	{8'd70,8'd155} : s = 204;
	{8'd70,8'd156} : s = 202;
	{8'd70,8'd157} : s = 346;
	{8'd70,8'd158} : s = 201;
	{8'd70,8'd159} : s = 345;
	{8'd70,8'd160} : s = 342;
	{8'd70,8'd161} : s = 459;
	{8'd70,8'd162} : s = 198;
	{8'd70,8'd163} : s = 341;
	{8'd70,8'd164} : s = 339;
	{8'd70,8'd165} : s = 455;
	{8'd70,8'd166} : s = 334;
	{8'd70,8'd167} : s = 444;
	{8'd70,8'd168} : s = 442;
	{8'd70,8'd169} : s = 502;
	{8'd70,8'd170} : s = 197;
	{8'd70,8'd171} : s = 333;
	{8'd70,8'd172} : s = 331;
	{8'd70,8'd173} : s = 441;
	{8'd70,8'd174} : s = 327;
	{8'd70,8'd175} : s = 438;
	{8'd70,8'd176} : s = 437;
	{8'd70,8'd177} : s = 501;
	{8'd70,8'd178} : s = 316;
	{8'd70,8'd179} : s = 435;
	{8'd70,8'd180} : s = 430;
	{8'd70,8'd181} : s = 499;
	{8'd70,8'd182} : s = 429;
	{8'd70,8'd183} : s = 494;
	{8'd70,8'd184} : s = 493;
	{8'd70,8'd185} : s = 510;
	{8'd70,8'd186} : s = 1;
	{8'd70,8'd187} : s = 18;
	{8'd70,8'd188} : s = 17;
	{8'd70,8'd189} : s = 82;
	{8'd70,8'd190} : s = 12;
	{8'd70,8'd191} : s = 81;
	{8'd70,8'd192} : s = 76;
	{8'd70,8'd193} : s = 195;
	{8'd70,8'd194} : s = 10;
	{8'd70,8'd195} : s = 74;
	{8'd70,8'd196} : s = 73;
	{8'd70,8'd197} : s = 184;
	{8'd70,8'd198} : s = 70;
	{8'd70,8'd199} : s = 180;
	{8'd70,8'd200} : s = 178;
	{8'd70,8'd201} : s = 314;
	{8'd70,8'd202} : s = 9;
	{8'd70,8'd203} : s = 69;
	{8'd70,8'd204} : s = 67;
	{8'd70,8'd205} : s = 177;
	{8'd70,8'd206} : s = 56;
	{8'd70,8'd207} : s = 172;
	{8'd70,8'd208} : s = 170;
	{8'd70,8'd209} : s = 313;
	{8'd70,8'd210} : s = 52;
	{8'd70,8'd211} : s = 169;
	{8'd70,8'd212} : s = 166;
	{8'd70,8'd213} : s = 310;
	{8'd70,8'd214} : s = 165;
	{8'd70,8'd215} : s = 309;
	{8'd70,8'd216} : s = 307;
	{8'd70,8'd217} : s = 427;
	{8'd70,8'd218} : s = 6;
	{8'd70,8'd219} : s = 50;
	{8'd70,8'd220} : s = 49;
	{8'd70,8'd221} : s = 163;
	{8'd70,8'd222} : s = 44;
	{8'd70,8'd223} : s = 156;
	{8'd70,8'd224} : s = 154;
	{8'd70,8'd225} : s = 302;
	{8'd70,8'd226} : s = 42;
	{8'd70,8'd227} : s = 153;
	{8'd70,8'd228} : s = 150;
	{8'd70,8'd229} : s = 301;
	{8'd70,8'd230} : s = 149;
	{8'd70,8'd231} : s = 299;
	{8'd70,8'd232} : s = 295;
	{8'd70,8'd233} : s = 423;
	{8'd70,8'd234} : s = 41;
	{8'd70,8'd235} : s = 147;
	{8'd70,8'd236} : s = 142;
	{8'd70,8'd237} : s = 286;
	{8'd70,8'd238} : s = 141;
	{8'd70,8'd239} : s = 285;
	{8'd70,8'd240} : s = 283;
	{8'd70,8'd241} : s = 414;
	{8'd70,8'd242} : s = 139;
	{8'd70,8'd243} : s = 279;
	{8'd70,8'd244} : s = 271;
	{8'd70,8'd245} : s = 413;
	{8'd70,8'd246} : s = 248;
	{8'd70,8'd247} : s = 411;
	{8'd70,8'd248} : s = 407;
	{8'd70,8'd249} : s = 491;
	{8'd70,8'd250} : s = 5;
	{8'd70,8'd251} : s = 38;
	{8'd70,8'd252} : s = 37;
	{8'd70,8'd253} : s = 135;
	{8'd70,8'd254} : s = 35;
	{8'd70,8'd255} : s = 120;
	{8'd71,8'd0} : s = 396;
	{8'd71,8'd1} : s = 68;
	{8'd71,8'd2} : s = 266;
	{8'd71,8'd3} : s = 265;
	{8'd71,8'd4} : s = 394;
	{8'd71,8'd5} : s = 262;
	{8'd71,8'd6} : s = 393;
	{8'd71,8'd7} : s = 390;
	{8'd71,8'd8} : s = 468;
	{8'd71,8'd9} : s = 66;
	{8'd71,8'd10} : s = 261;
	{8'd71,8'd11} : s = 259;
	{8'd71,8'd12} : s = 389;
	{8'd71,8'd13} : s = 224;
	{8'd71,8'd14} : s = 387;
	{8'd71,8'd15} : s = 368;
	{8'd71,8'd16} : s = 466;
	{8'd71,8'd17} : s = 208;
	{8'd71,8'd18} : s = 360;
	{8'd71,8'd19} : s = 356;
	{8'd71,8'd20} : s = 465;
	{8'd71,8'd21} : s = 354;
	{8'd71,8'd22} : s = 460;
	{8'd71,8'd23} : s = 458;
	{8'd71,8'd24} : s = 500;
	{8'd71,8'd25} : s = 65;
	{8'd71,8'd26} : s = 200;
	{8'd71,8'd27} : s = 196;
	{8'd71,8'd28} : s = 353;
	{8'd71,8'd29} : s = 194;
	{8'd71,8'd30} : s = 344;
	{8'd71,8'd31} : s = 340;
	{8'd71,8'd32} : s = 457;
	{8'd71,8'd33} : s = 193;
	{8'd71,8'd34} : s = 338;
	{8'd71,8'd35} : s = 337;
	{8'd71,8'd36} : s = 454;
	{8'd71,8'd37} : s = 332;
	{8'd71,8'd38} : s = 453;
	{8'd71,8'd39} : s = 451;
	{8'd71,8'd40} : s = 498;
	{8'd71,8'd41} : s = 176;
	{8'd71,8'd42} : s = 330;
	{8'd71,8'd43} : s = 329;
	{8'd71,8'd44} : s = 440;
	{8'd71,8'd45} : s = 326;
	{8'd71,8'd46} : s = 436;
	{8'd71,8'd47} : s = 434;
	{8'd71,8'd48} : s = 497;
	{8'd71,8'd49} : s = 325;
	{8'd71,8'd50} : s = 433;
	{8'd71,8'd51} : s = 428;
	{8'd71,8'd52} : s = 492;
	{8'd71,8'd53} : s = 426;
	{8'd71,8'd54} : s = 490;
	{8'd71,8'd55} : s = 489;
	{8'd71,8'd56} : s = 508;
	{8'd71,8'd57} : s = 2;
	{8'd71,8'd58} : s = 48;
	{8'd71,8'd59} : s = 40;
	{8'd71,8'd60} : s = 168;
	{8'd71,8'd61} : s = 36;
	{8'd71,8'd62} : s = 164;
	{8'd71,8'd63} : s = 162;
	{8'd71,8'd64} : s = 323;
	{8'd71,8'd65} : s = 34;
	{8'd71,8'd66} : s = 161;
	{8'd71,8'd67} : s = 152;
	{8'd71,8'd68} : s = 312;
	{8'd71,8'd69} : s = 148;
	{8'd71,8'd70} : s = 308;
	{8'd71,8'd71} : s = 306;
	{8'd71,8'd72} : s = 425;
	{8'd71,8'd73} : s = 33;
	{8'd71,8'd74} : s = 146;
	{8'd71,8'd75} : s = 145;
	{8'd71,8'd76} : s = 305;
	{8'd71,8'd77} : s = 140;
	{8'd71,8'd78} : s = 300;
	{8'd71,8'd79} : s = 298;
	{8'd71,8'd80} : s = 422;
	{8'd71,8'd81} : s = 138;
	{8'd71,8'd82} : s = 297;
	{8'd71,8'd83} : s = 294;
	{8'd71,8'd84} : s = 421;
	{8'd71,8'd85} : s = 293;
	{8'd71,8'd86} : s = 419;
	{8'd71,8'd87} : s = 412;
	{8'd71,8'd88} : s = 486;
	{8'd71,8'd89} : s = 24;
	{8'd71,8'd90} : s = 137;
	{8'd71,8'd91} : s = 134;
	{8'd71,8'd92} : s = 291;
	{8'd71,8'd93} : s = 133;
	{8'd71,8'd94} : s = 284;
	{8'd71,8'd95} : s = 282;
	{8'd71,8'd96} : s = 410;
	{8'd71,8'd97} : s = 131;
	{8'd71,8'd98} : s = 281;
	{8'd71,8'd99} : s = 278;
	{8'd71,8'd100} : s = 409;
	{8'd71,8'd101} : s = 277;
	{8'd71,8'd102} : s = 406;
	{8'd71,8'd103} : s = 405;
	{8'd71,8'd104} : s = 485;
	{8'd71,8'd105} : s = 112;
	{8'd71,8'd106} : s = 275;
	{8'd71,8'd107} : s = 270;
	{8'd71,8'd108} : s = 403;
	{8'd71,8'd109} : s = 269;
	{8'd71,8'd110} : s = 398;
	{8'd71,8'd111} : s = 397;
	{8'd71,8'd112} : s = 483;
	{8'd71,8'd113} : s = 267;
	{8'd71,8'd114} : s = 395;
	{8'd71,8'd115} : s = 391;
	{8'd71,8'd116} : s = 476;
	{8'd71,8'd117} : s = 376;
	{8'd71,8'd118} : s = 474;
	{8'd71,8'd119} : s = 473;
	{8'd71,8'd120} : s = 506;
	{8'd71,8'd121} : s = 20;
	{8'd71,8'd122} : s = 104;
	{8'd71,8'd123} : s = 100;
	{8'd71,8'd124} : s = 263;
	{8'd71,8'd125} : s = 98;
	{8'd71,8'd126} : s = 240;
	{8'd71,8'd127} : s = 232;
	{8'd71,8'd128} : s = 372;
	{8'd71,8'd129} : s = 97;
	{8'd71,8'd130} : s = 228;
	{8'd71,8'd131} : s = 226;
	{8'd71,8'd132} : s = 370;
	{8'd71,8'd133} : s = 225;
	{8'd71,8'd134} : s = 369;
	{8'd71,8'd135} : s = 364;
	{8'd71,8'd136} : s = 470;
	{8'd71,8'd137} : s = 88;
	{8'd71,8'd138} : s = 216;
	{8'd71,8'd139} : s = 212;
	{8'd71,8'd140} : s = 362;
	{8'd71,8'd141} : s = 210;
	{8'd71,8'd142} : s = 361;
	{8'd71,8'd143} : s = 358;
	{8'd71,8'd144} : s = 469;
	{8'd71,8'd145} : s = 209;
	{8'd71,8'd146} : s = 357;
	{8'd71,8'd147} : s = 355;
	{8'd71,8'd148} : s = 467;
	{8'd71,8'd149} : s = 348;
	{8'd71,8'd150} : s = 462;
	{8'd71,8'd151} : s = 461;
	{8'd71,8'd152} : s = 505;
	{8'd71,8'd153} : s = 84;
	{8'd71,8'd154} : s = 204;
	{8'd71,8'd155} : s = 202;
	{8'd71,8'd156} : s = 346;
	{8'd71,8'd157} : s = 201;
	{8'd71,8'd158} : s = 345;
	{8'd71,8'd159} : s = 342;
	{8'd71,8'd160} : s = 459;
	{8'd71,8'd161} : s = 198;
	{8'd71,8'd162} : s = 341;
	{8'd71,8'd163} : s = 339;
	{8'd71,8'd164} : s = 455;
	{8'd71,8'd165} : s = 334;
	{8'd71,8'd166} : s = 444;
	{8'd71,8'd167} : s = 442;
	{8'd71,8'd168} : s = 502;
	{8'd71,8'd169} : s = 197;
	{8'd71,8'd170} : s = 333;
	{8'd71,8'd171} : s = 331;
	{8'd71,8'd172} : s = 441;
	{8'd71,8'd173} : s = 327;
	{8'd71,8'd174} : s = 438;
	{8'd71,8'd175} : s = 437;
	{8'd71,8'd176} : s = 501;
	{8'd71,8'd177} : s = 316;
	{8'd71,8'd178} : s = 435;
	{8'd71,8'd179} : s = 430;
	{8'd71,8'd180} : s = 499;
	{8'd71,8'd181} : s = 429;
	{8'd71,8'd182} : s = 494;
	{8'd71,8'd183} : s = 493;
	{8'd71,8'd184} : s = 510;
	{8'd71,8'd185} : s = 1;
	{8'd71,8'd186} : s = 18;
	{8'd71,8'd187} : s = 17;
	{8'd71,8'd188} : s = 82;
	{8'd71,8'd189} : s = 12;
	{8'd71,8'd190} : s = 81;
	{8'd71,8'd191} : s = 76;
	{8'd71,8'd192} : s = 195;
	{8'd71,8'd193} : s = 10;
	{8'd71,8'd194} : s = 74;
	{8'd71,8'd195} : s = 73;
	{8'd71,8'd196} : s = 184;
	{8'd71,8'd197} : s = 70;
	{8'd71,8'd198} : s = 180;
	{8'd71,8'd199} : s = 178;
	{8'd71,8'd200} : s = 314;
	{8'd71,8'd201} : s = 9;
	{8'd71,8'd202} : s = 69;
	{8'd71,8'd203} : s = 67;
	{8'd71,8'd204} : s = 177;
	{8'd71,8'd205} : s = 56;
	{8'd71,8'd206} : s = 172;
	{8'd71,8'd207} : s = 170;
	{8'd71,8'd208} : s = 313;
	{8'd71,8'd209} : s = 52;
	{8'd71,8'd210} : s = 169;
	{8'd71,8'd211} : s = 166;
	{8'd71,8'd212} : s = 310;
	{8'd71,8'd213} : s = 165;
	{8'd71,8'd214} : s = 309;
	{8'd71,8'd215} : s = 307;
	{8'd71,8'd216} : s = 427;
	{8'd71,8'd217} : s = 6;
	{8'd71,8'd218} : s = 50;
	{8'd71,8'd219} : s = 49;
	{8'd71,8'd220} : s = 163;
	{8'd71,8'd221} : s = 44;
	{8'd71,8'd222} : s = 156;
	{8'd71,8'd223} : s = 154;
	{8'd71,8'd224} : s = 302;
	{8'd71,8'd225} : s = 42;
	{8'd71,8'd226} : s = 153;
	{8'd71,8'd227} : s = 150;
	{8'd71,8'd228} : s = 301;
	{8'd71,8'd229} : s = 149;
	{8'd71,8'd230} : s = 299;
	{8'd71,8'd231} : s = 295;
	{8'd71,8'd232} : s = 423;
	{8'd71,8'd233} : s = 41;
	{8'd71,8'd234} : s = 147;
	{8'd71,8'd235} : s = 142;
	{8'd71,8'd236} : s = 286;
	{8'd71,8'd237} : s = 141;
	{8'd71,8'd238} : s = 285;
	{8'd71,8'd239} : s = 283;
	{8'd71,8'd240} : s = 414;
	{8'd71,8'd241} : s = 139;
	{8'd71,8'd242} : s = 279;
	{8'd71,8'd243} : s = 271;
	{8'd71,8'd244} : s = 413;
	{8'd71,8'd245} : s = 248;
	{8'd71,8'd246} : s = 411;
	{8'd71,8'd247} : s = 407;
	{8'd71,8'd248} : s = 491;
	{8'd71,8'd249} : s = 5;
	{8'd71,8'd250} : s = 38;
	{8'd71,8'd251} : s = 37;
	{8'd71,8'd252} : s = 135;
	{8'd71,8'd253} : s = 35;
	{8'd71,8'd254} : s = 120;
	{8'd71,8'd255} : s = 116;
	{8'd72,8'd0} : s = 68;
	{8'd72,8'd1} : s = 266;
	{8'd72,8'd2} : s = 265;
	{8'd72,8'd3} : s = 394;
	{8'd72,8'd4} : s = 262;
	{8'd72,8'd5} : s = 393;
	{8'd72,8'd6} : s = 390;
	{8'd72,8'd7} : s = 468;
	{8'd72,8'd8} : s = 66;
	{8'd72,8'd9} : s = 261;
	{8'd72,8'd10} : s = 259;
	{8'd72,8'd11} : s = 389;
	{8'd72,8'd12} : s = 224;
	{8'd72,8'd13} : s = 387;
	{8'd72,8'd14} : s = 368;
	{8'd72,8'd15} : s = 466;
	{8'd72,8'd16} : s = 208;
	{8'd72,8'd17} : s = 360;
	{8'd72,8'd18} : s = 356;
	{8'd72,8'd19} : s = 465;
	{8'd72,8'd20} : s = 354;
	{8'd72,8'd21} : s = 460;
	{8'd72,8'd22} : s = 458;
	{8'd72,8'd23} : s = 500;
	{8'd72,8'd24} : s = 65;
	{8'd72,8'd25} : s = 200;
	{8'd72,8'd26} : s = 196;
	{8'd72,8'd27} : s = 353;
	{8'd72,8'd28} : s = 194;
	{8'd72,8'd29} : s = 344;
	{8'd72,8'd30} : s = 340;
	{8'd72,8'd31} : s = 457;
	{8'd72,8'd32} : s = 193;
	{8'd72,8'd33} : s = 338;
	{8'd72,8'd34} : s = 337;
	{8'd72,8'd35} : s = 454;
	{8'd72,8'd36} : s = 332;
	{8'd72,8'd37} : s = 453;
	{8'd72,8'd38} : s = 451;
	{8'd72,8'd39} : s = 498;
	{8'd72,8'd40} : s = 176;
	{8'd72,8'd41} : s = 330;
	{8'd72,8'd42} : s = 329;
	{8'd72,8'd43} : s = 440;
	{8'd72,8'd44} : s = 326;
	{8'd72,8'd45} : s = 436;
	{8'd72,8'd46} : s = 434;
	{8'd72,8'd47} : s = 497;
	{8'd72,8'd48} : s = 325;
	{8'd72,8'd49} : s = 433;
	{8'd72,8'd50} : s = 428;
	{8'd72,8'd51} : s = 492;
	{8'd72,8'd52} : s = 426;
	{8'd72,8'd53} : s = 490;
	{8'd72,8'd54} : s = 489;
	{8'd72,8'd55} : s = 508;
	{8'd72,8'd56} : s = 2;
	{8'd72,8'd57} : s = 48;
	{8'd72,8'd58} : s = 40;
	{8'd72,8'd59} : s = 168;
	{8'd72,8'd60} : s = 36;
	{8'd72,8'd61} : s = 164;
	{8'd72,8'd62} : s = 162;
	{8'd72,8'd63} : s = 323;
	{8'd72,8'd64} : s = 34;
	{8'd72,8'd65} : s = 161;
	{8'd72,8'd66} : s = 152;
	{8'd72,8'd67} : s = 312;
	{8'd72,8'd68} : s = 148;
	{8'd72,8'd69} : s = 308;
	{8'd72,8'd70} : s = 306;
	{8'd72,8'd71} : s = 425;
	{8'd72,8'd72} : s = 33;
	{8'd72,8'd73} : s = 146;
	{8'd72,8'd74} : s = 145;
	{8'd72,8'd75} : s = 305;
	{8'd72,8'd76} : s = 140;
	{8'd72,8'd77} : s = 300;
	{8'd72,8'd78} : s = 298;
	{8'd72,8'd79} : s = 422;
	{8'd72,8'd80} : s = 138;
	{8'd72,8'd81} : s = 297;
	{8'd72,8'd82} : s = 294;
	{8'd72,8'd83} : s = 421;
	{8'd72,8'd84} : s = 293;
	{8'd72,8'd85} : s = 419;
	{8'd72,8'd86} : s = 412;
	{8'd72,8'd87} : s = 486;
	{8'd72,8'd88} : s = 24;
	{8'd72,8'd89} : s = 137;
	{8'd72,8'd90} : s = 134;
	{8'd72,8'd91} : s = 291;
	{8'd72,8'd92} : s = 133;
	{8'd72,8'd93} : s = 284;
	{8'd72,8'd94} : s = 282;
	{8'd72,8'd95} : s = 410;
	{8'd72,8'd96} : s = 131;
	{8'd72,8'd97} : s = 281;
	{8'd72,8'd98} : s = 278;
	{8'd72,8'd99} : s = 409;
	{8'd72,8'd100} : s = 277;
	{8'd72,8'd101} : s = 406;
	{8'd72,8'd102} : s = 405;
	{8'd72,8'd103} : s = 485;
	{8'd72,8'd104} : s = 112;
	{8'd72,8'd105} : s = 275;
	{8'd72,8'd106} : s = 270;
	{8'd72,8'd107} : s = 403;
	{8'd72,8'd108} : s = 269;
	{8'd72,8'd109} : s = 398;
	{8'd72,8'd110} : s = 397;
	{8'd72,8'd111} : s = 483;
	{8'd72,8'd112} : s = 267;
	{8'd72,8'd113} : s = 395;
	{8'd72,8'd114} : s = 391;
	{8'd72,8'd115} : s = 476;
	{8'd72,8'd116} : s = 376;
	{8'd72,8'd117} : s = 474;
	{8'd72,8'd118} : s = 473;
	{8'd72,8'd119} : s = 506;
	{8'd72,8'd120} : s = 20;
	{8'd72,8'd121} : s = 104;
	{8'd72,8'd122} : s = 100;
	{8'd72,8'd123} : s = 263;
	{8'd72,8'd124} : s = 98;
	{8'd72,8'd125} : s = 240;
	{8'd72,8'd126} : s = 232;
	{8'd72,8'd127} : s = 372;
	{8'd72,8'd128} : s = 97;
	{8'd72,8'd129} : s = 228;
	{8'd72,8'd130} : s = 226;
	{8'd72,8'd131} : s = 370;
	{8'd72,8'd132} : s = 225;
	{8'd72,8'd133} : s = 369;
	{8'd72,8'd134} : s = 364;
	{8'd72,8'd135} : s = 470;
	{8'd72,8'd136} : s = 88;
	{8'd72,8'd137} : s = 216;
	{8'd72,8'd138} : s = 212;
	{8'd72,8'd139} : s = 362;
	{8'd72,8'd140} : s = 210;
	{8'd72,8'd141} : s = 361;
	{8'd72,8'd142} : s = 358;
	{8'd72,8'd143} : s = 469;
	{8'd72,8'd144} : s = 209;
	{8'd72,8'd145} : s = 357;
	{8'd72,8'd146} : s = 355;
	{8'd72,8'd147} : s = 467;
	{8'd72,8'd148} : s = 348;
	{8'd72,8'd149} : s = 462;
	{8'd72,8'd150} : s = 461;
	{8'd72,8'd151} : s = 505;
	{8'd72,8'd152} : s = 84;
	{8'd72,8'd153} : s = 204;
	{8'd72,8'd154} : s = 202;
	{8'd72,8'd155} : s = 346;
	{8'd72,8'd156} : s = 201;
	{8'd72,8'd157} : s = 345;
	{8'd72,8'd158} : s = 342;
	{8'd72,8'd159} : s = 459;
	{8'd72,8'd160} : s = 198;
	{8'd72,8'd161} : s = 341;
	{8'd72,8'd162} : s = 339;
	{8'd72,8'd163} : s = 455;
	{8'd72,8'd164} : s = 334;
	{8'd72,8'd165} : s = 444;
	{8'd72,8'd166} : s = 442;
	{8'd72,8'd167} : s = 502;
	{8'd72,8'd168} : s = 197;
	{8'd72,8'd169} : s = 333;
	{8'd72,8'd170} : s = 331;
	{8'd72,8'd171} : s = 441;
	{8'd72,8'd172} : s = 327;
	{8'd72,8'd173} : s = 438;
	{8'd72,8'd174} : s = 437;
	{8'd72,8'd175} : s = 501;
	{8'd72,8'd176} : s = 316;
	{8'd72,8'd177} : s = 435;
	{8'd72,8'd178} : s = 430;
	{8'd72,8'd179} : s = 499;
	{8'd72,8'd180} : s = 429;
	{8'd72,8'd181} : s = 494;
	{8'd72,8'd182} : s = 493;
	{8'd72,8'd183} : s = 510;
	{8'd72,8'd184} : s = 1;
	{8'd72,8'd185} : s = 18;
	{8'd72,8'd186} : s = 17;
	{8'd72,8'd187} : s = 82;
	{8'd72,8'd188} : s = 12;
	{8'd72,8'd189} : s = 81;
	{8'd72,8'd190} : s = 76;
	{8'd72,8'd191} : s = 195;
	{8'd72,8'd192} : s = 10;
	{8'd72,8'd193} : s = 74;
	{8'd72,8'd194} : s = 73;
	{8'd72,8'd195} : s = 184;
	{8'd72,8'd196} : s = 70;
	{8'd72,8'd197} : s = 180;
	{8'd72,8'd198} : s = 178;
	{8'd72,8'd199} : s = 314;
	{8'd72,8'd200} : s = 9;
	{8'd72,8'd201} : s = 69;
	{8'd72,8'd202} : s = 67;
	{8'd72,8'd203} : s = 177;
	{8'd72,8'd204} : s = 56;
	{8'd72,8'd205} : s = 172;
	{8'd72,8'd206} : s = 170;
	{8'd72,8'd207} : s = 313;
	{8'd72,8'd208} : s = 52;
	{8'd72,8'd209} : s = 169;
	{8'd72,8'd210} : s = 166;
	{8'd72,8'd211} : s = 310;
	{8'd72,8'd212} : s = 165;
	{8'd72,8'd213} : s = 309;
	{8'd72,8'd214} : s = 307;
	{8'd72,8'd215} : s = 427;
	{8'd72,8'd216} : s = 6;
	{8'd72,8'd217} : s = 50;
	{8'd72,8'd218} : s = 49;
	{8'd72,8'd219} : s = 163;
	{8'd72,8'd220} : s = 44;
	{8'd72,8'd221} : s = 156;
	{8'd72,8'd222} : s = 154;
	{8'd72,8'd223} : s = 302;
	{8'd72,8'd224} : s = 42;
	{8'd72,8'd225} : s = 153;
	{8'd72,8'd226} : s = 150;
	{8'd72,8'd227} : s = 301;
	{8'd72,8'd228} : s = 149;
	{8'd72,8'd229} : s = 299;
	{8'd72,8'd230} : s = 295;
	{8'd72,8'd231} : s = 423;
	{8'd72,8'd232} : s = 41;
	{8'd72,8'd233} : s = 147;
	{8'd72,8'd234} : s = 142;
	{8'd72,8'd235} : s = 286;
	{8'd72,8'd236} : s = 141;
	{8'd72,8'd237} : s = 285;
	{8'd72,8'd238} : s = 283;
	{8'd72,8'd239} : s = 414;
	{8'd72,8'd240} : s = 139;
	{8'd72,8'd241} : s = 279;
	{8'd72,8'd242} : s = 271;
	{8'd72,8'd243} : s = 413;
	{8'd72,8'd244} : s = 248;
	{8'd72,8'd245} : s = 411;
	{8'd72,8'd246} : s = 407;
	{8'd72,8'd247} : s = 491;
	{8'd72,8'd248} : s = 5;
	{8'd72,8'd249} : s = 38;
	{8'd72,8'd250} : s = 37;
	{8'd72,8'd251} : s = 135;
	{8'd72,8'd252} : s = 35;
	{8'd72,8'd253} : s = 120;
	{8'd72,8'd254} : s = 116;
	{8'd72,8'd255} : s = 244;
	{8'd73,8'd0} : s = 266;
	{8'd73,8'd1} : s = 265;
	{8'd73,8'd2} : s = 394;
	{8'd73,8'd3} : s = 262;
	{8'd73,8'd4} : s = 393;
	{8'd73,8'd5} : s = 390;
	{8'd73,8'd6} : s = 468;
	{8'd73,8'd7} : s = 66;
	{8'd73,8'd8} : s = 261;
	{8'd73,8'd9} : s = 259;
	{8'd73,8'd10} : s = 389;
	{8'd73,8'd11} : s = 224;
	{8'd73,8'd12} : s = 387;
	{8'd73,8'd13} : s = 368;
	{8'd73,8'd14} : s = 466;
	{8'd73,8'd15} : s = 208;
	{8'd73,8'd16} : s = 360;
	{8'd73,8'd17} : s = 356;
	{8'd73,8'd18} : s = 465;
	{8'd73,8'd19} : s = 354;
	{8'd73,8'd20} : s = 460;
	{8'd73,8'd21} : s = 458;
	{8'd73,8'd22} : s = 500;
	{8'd73,8'd23} : s = 65;
	{8'd73,8'd24} : s = 200;
	{8'd73,8'd25} : s = 196;
	{8'd73,8'd26} : s = 353;
	{8'd73,8'd27} : s = 194;
	{8'd73,8'd28} : s = 344;
	{8'd73,8'd29} : s = 340;
	{8'd73,8'd30} : s = 457;
	{8'd73,8'd31} : s = 193;
	{8'd73,8'd32} : s = 338;
	{8'd73,8'd33} : s = 337;
	{8'd73,8'd34} : s = 454;
	{8'd73,8'd35} : s = 332;
	{8'd73,8'd36} : s = 453;
	{8'd73,8'd37} : s = 451;
	{8'd73,8'd38} : s = 498;
	{8'd73,8'd39} : s = 176;
	{8'd73,8'd40} : s = 330;
	{8'd73,8'd41} : s = 329;
	{8'd73,8'd42} : s = 440;
	{8'd73,8'd43} : s = 326;
	{8'd73,8'd44} : s = 436;
	{8'd73,8'd45} : s = 434;
	{8'd73,8'd46} : s = 497;
	{8'd73,8'd47} : s = 325;
	{8'd73,8'd48} : s = 433;
	{8'd73,8'd49} : s = 428;
	{8'd73,8'd50} : s = 492;
	{8'd73,8'd51} : s = 426;
	{8'd73,8'd52} : s = 490;
	{8'd73,8'd53} : s = 489;
	{8'd73,8'd54} : s = 508;
	{8'd73,8'd55} : s = 2;
	{8'd73,8'd56} : s = 48;
	{8'd73,8'd57} : s = 40;
	{8'd73,8'd58} : s = 168;
	{8'd73,8'd59} : s = 36;
	{8'd73,8'd60} : s = 164;
	{8'd73,8'd61} : s = 162;
	{8'd73,8'd62} : s = 323;
	{8'd73,8'd63} : s = 34;
	{8'd73,8'd64} : s = 161;
	{8'd73,8'd65} : s = 152;
	{8'd73,8'd66} : s = 312;
	{8'd73,8'd67} : s = 148;
	{8'd73,8'd68} : s = 308;
	{8'd73,8'd69} : s = 306;
	{8'd73,8'd70} : s = 425;
	{8'd73,8'd71} : s = 33;
	{8'd73,8'd72} : s = 146;
	{8'd73,8'd73} : s = 145;
	{8'd73,8'd74} : s = 305;
	{8'd73,8'd75} : s = 140;
	{8'd73,8'd76} : s = 300;
	{8'd73,8'd77} : s = 298;
	{8'd73,8'd78} : s = 422;
	{8'd73,8'd79} : s = 138;
	{8'd73,8'd80} : s = 297;
	{8'd73,8'd81} : s = 294;
	{8'd73,8'd82} : s = 421;
	{8'd73,8'd83} : s = 293;
	{8'd73,8'd84} : s = 419;
	{8'd73,8'd85} : s = 412;
	{8'd73,8'd86} : s = 486;
	{8'd73,8'd87} : s = 24;
	{8'd73,8'd88} : s = 137;
	{8'd73,8'd89} : s = 134;
	{8'd73,8'd90} : s = 291;
	{8'd73,8'd91} : s = 133;
	{8'd73,8'd92} : s = 284;
	{8'd73,8'd93} : s = 282;
	{8'd73,8'd94} : s = 410;
	{8'd73,8'd95} : s = 131;
	{8'd73,8'd96} : s = 281;
	{8'd73,8'd97} : s = 278;
	{8'd73,8'd98} : s = 409;
	{8'd73,8'd99} : s = 277;
	{8'd73,8'd100} : s = 406;
	{8'd73,8'd101} : s = 405;
	{8'd73,8'd102} : s = 485;
	{8'd73,8'd103} : s = 112;
	{8'd73,8'd104} : s = 275;
	{8'd73,8'd105} : s = 270;
	{8'd73,8'd106} : s = 403;
	{8'd73,8'd107} : s = 269;
	{8'd73,8'd108} : s = 398;
	{8'd73,8'd109} : s = 397;
	{8'd73,8'd110} : s = 483;
	{8'd73,8'd111} : s = 267;
	{8'd73,8'd112} : s = 395;
	{8'd73,8'd113} : s = 391;
	{8'd73,8'd114} : s = 476;
	{8'd73,8'd115} : s = 376;
	{8'd73,8'd116} : s = 474;
	{8'd73,8'd117} : s = 473;
	{8'd73,8'd118} : s = 506;
	{8'd73,8'd119} : s = 20;
	{8'd73,8'd120} : s = 104;
	{8'd73,8'd121} : s = 100;
	{8'd73,8'd122} : s = 263;
	{8'd73,8'd123} : s = 98;
	{8'd73,8'd124} : s = 240;
	{8'd73,8'd125} : s = 232;
	{8'd73,8'd126} : s = 372;
	{8'd73,8'd127} : s = 97;
	{8'd73,8'd128} : s = 228;
	{8'd73,8'd129} : s = 226;
	{8'd73,8'd130} : s = 370;
	{8'd73,8'd131} : s = 225;
	{8'd73,8'd132} : s = 369;
	{8'd73,8'd133} : s = 364;
	{8'd73,8'd134} : s = 470;
	{8'd73,8'd135} : s = 88;
	{8'd73,8'd136} : s = 216;
	{8'd73,8'd137} : s = 212;
	{8'd73,8'd138} : s = 362;
	{8'd73,8'd139} : s = 210;
	{8'd73,8'd140} : s = 361;
	{8'd73,8'd141} : s = 358;
	{8'd73,8'd142} : s = 469;
	{8'd73,8'd143} : s = 209;
	{8'd73,8'd144} : s = 357;
	{8'd73,8'd145} : s = 355;
	{8'd73,8'd146} : s = 467;
	{8'd73,8'd147} : s = 348;
	{8'd73,8'd148} : s = 462;
	{8'd73,8'd149} : s = 461;
	{8'd73,8'd150} : s = 505;
	{8'd73,8'd151} : s = 84;
	{8'd73,8'd152} : s = 204;
	{8'd73,8'd153} : s = 202;
	{8'd73,8'd154} : s = 346;
	{8'd73,8'd155} : s = 201;
	{8'd73,8'd156} : s = 345;
	{8'd73,8'd157} : s = 342;
	{8'd73,8'd158} : s = 459;
	{8'd73,8'd159} : s = 198;
	{8'd73,8'd160} : s = 341;
	{8'd73,8'd161} : s = 339;
	{8'd73,8'd162} : s = 455;
	{8'd73,8'd163} : s = 334;
	{8'd73,8'd164} : s = 444;
	{8'd73,8'd165} : s = 442;
	{8'd73,8'd166} : s = 502;
	{8'd73,8'd167} : s = 197;
	{8'd73,8'd168} : s = 333;
	{8'd73,8'd169} : s = 331;
	{8'd73,8'd170} : s = 441;
	{8'd73,8'd171} : s = 327;
	{8'd73,8'd172} : s = 438;
	{8'd73,8'd173} : s = 437;
	{8'd73,8'd174} : s = 501;
	{8'd73,8'd175} : s = 316;
	{8'd73,8'd176} : s = 435;
	{8'd73,8'd177} : s = 430;
	{8'd73,8'd178} : s = 499;
	{8'd73,8'd179} : s = 429;
	{8'd73,8'd180} : s = 494;
	{8'd73,8'd181} : s = 493;
	{8'd73,8'd182} : s = 510;
	{8'd73,8'd183} : s = 1;
	{8'd73,8'd184} : s = 18;
	{8'd73,8'd185} : s = 17;
	{8'd73,8'd186} : s = 82;
	{8'd73,8'd187} : s = 12;
	{8'd73,8'd188} : s = 81;
	{8'd73,8'd189} : s = 76;
	{8'd73,8'd190} : s = 195;
	{8'd73,8'd191} : s = 10;
	{8'd73,8'd192} : s = 74;
	{8'd73,8'd193} : s = 73;
	{8'd73,8'd194} : s = 184;
	{8'd73,8'd195} : s = 70;
	{8'd73,8'd196} : s = 180;
	{8'd73,8'd197} : s = 178;
	{8'd73,8'd198} : s = 314;
	{8'd73,8'd199} : s = 9;
	{8'd73,8'd200} : s = 69;
	{8'd73,8'd201} : s = 67;
	{8'd73,8'd202} : s = 177;
	{8'd73,8'd203} : s = 56;
	{8'd73,8'd204} : s = 172;
	{8'd73,8'd205} : s = 170;
	{8'd73,8'd206} : s = 313;
	{8'd73,8'd207} : s = 52;
	{8'd73,8'd208} : s = 169;
	{8'd73,8'd209} : s = 166;
	{8'd73,8'd210} : s = 310;
	{8'd73,8'd211} : s = 165;
	{8'd73,8'd212} : s = 309;
	{8'd73,8'd213} : s = 307;
	{8'd73,8'd214} : s = 427;
	{8'd73,8'd215} : s = 6;
	{8'd73,8'd216} : s = 50;
	{8'd73,8'd217} : s = 49;
	{8'd73,8'd218} : s = 163;
	{8'd73,8'd219} : s = 44;
	{8'd73,8'd220} : s = 156;
	{8'd73,8'd221} : s = 154;
	{8'd73,8'd222} : s = 302;
	{8'd73,8'd223} : s = 42;
	{8'd73,8'd224} : s = 153;
	{8'd73,8'd225} : s = 150;
	{8'd73,8'd226} : s = 301;
	{8'd73,8'd227} : s = 149;
	{8'd73,8'd228} : s = 299;
	{8'd73,8'd229} : s = 295;
	{8'd73,8'd230} : s = 423;
	{8'd73,8'd231} : s = 41;
	{8'd73,8'd232} : s = 147;
	{8'd73,8'd233} : s = 142;
	{8'd73,8'd234} : s = 286;
	{8'd73,8'd235} : s = 141;
	{8'd73,8'd236} : s = 285;
	{8'd73,8'd237} : s = 283;
	{8'd73,8'd238} : s = 414;
	{8'd73,8'd239} : s = 139;
	{8'd73,8'd240} : s = 279;
	{8'd73,8'd241} : s = 271;
	{8'd73,8'd242} : s = 413;
	{8'd73,8'd243} : s = 248;
	{8'd73,8'd244} : s = 411;
	{8'd73,8'd245} : s = 407;
	{8'd73,8'd246} : s = 491;
	{8'd73,8'd247} : s = 5;
	{8'd73,8'd248} : s = 38;
	{8'd73,8'd249} : s = 37;
	{8'd73,8'd250} : s = 135;
	{8'd73,8'd251} : s = 35;
	{8'd73,8'd252} : s = 120;
	{8'd73,8'd253} : s = 116;
	{8'd73,8'd254} : s = 244;
	{8'd73,8'd255} : s = 28;
	{8'd74,8'd0} : s = 265;
	{8'd74,8'd1} : s = 394;
	{8'd74,8'd2} : s = 262;
	{8'd74,8'd3} : s = 393;
	{8'd74,8'd4} : s = 390;
	{8'd74,8'd5} : s = 468;
	{8'd74,8'd6} : s = 66;
	{8'd74,8'd7} : s = 261;
	{8'd74,8'd8} : s = 259;
	{8'd74,8'd9} : s = 389;
	{8'd74,8'd10} : s = 224;
	{8'd74,8'd11} : s = 387;
	{8'd74,8'd12} : s = 368;
	{8'd74,8'd13} : s = 466;
	{8'd74,8'd14} : s = 208;
	{8'd74,8'd15} : s = 360;
	{8'd74,8'd16} : s = 356;
	{8'd74,8'd17} : s = 465;
	{8'd74,8'd18} : s = 354;
	{8'd74,8'd19} : s = 460;
	{8'd74,8'd20} : s = 458;
	{8'd74,8'd21} : s = 500;
	{8'd74,8'd22} : s = 65;
	{8'd74,8'd23} : s = 200;
	{8'd74,8'd24} : s = 196;
	{8'd74,8'd25} : s = 353;
	{8'd74,8'd26} : s = 194;
	{8'd74,8'd27} : s = 344;
	{8'd74,8'd28} : s = 340;
	{8'd74,8'd29} : s = 457;
	{8'd74,8'd30} : s = 193;
	{8'd74,8'd31} : s = 338;
	{8'd74,8'd32} : s = 337;
	{8'd74,8'd33} : s = 454;
	{8'd74,8'd34} : s = 332;
	{8'd74,8'd35} : s = 453;
	{8'd74,8'd36} : s = 451;
	{8'd74,8'd37} : s = 498;
	{8'd74,8'd38} : s = 176;
	{8'd74,8'd39} : s = 330;
	{8'd74,8'd40} : s = 329;
	{8'd74,8'd41} : s = 440;
	{8'd74,8'd42} : s = 326;
	{8'd74,8'd43} : s = 436;
	{8'd74,8'd44} : s = 434;
	{8'd74,8'd45} : s = 497;
	{8'd74,8'd46} : s = 325;
	{8'd74,8'd47} : s = 433;
	{8'd74,8'd48} : s = 428;
	{8'd74,8'd49} : s = 492;
	{8'd74,8'd50} : s = 426;
	{8'd74,8'd51} : s = 490;
	{8'd74,8'd52} : s = 489;
	{8'd74,8'd53} : s = 508;
	{8'd74,8'd54} : s = 2;
	{8'd74,8'd55} : s = 48;
	{8'd74,8'd56} : s = 40;
	{8'd74,8'd57} : s = 168;
	{8'd74,8'd58} : s = 36;
	{8'd74,8'd59} : s = 164;
	{8'd74,8'd60} : s = 162;
	{8'd74,8'd61} : s = 323;
	{8'd74,8'd62} : s = 34;
	{8'd74,8'd63} : s = 161;
	{8'd74,8'd64} : s = 152;
	{8'd74,8'd65} : s = 312;
	{8'd74,8'd66} : s = 148;
	{8'd74,8'd67} : s = 308;
	{8'd74,8'd68} : s = 306;
	{8'd74,8'd69} : s = 425;
	{8'd74,8'd70} : s = 33;
	{8'd74,8'd71} : s = 146;
	{8'd74,8'd72} : s = 145;
	{8'd74,8'd73} : s = 305;
	{8'd74,8'd74} : s = 140;
	{8'd74,8'd75} : s = 300;
	{8'd74,8'd76} : s = 298;
	{8'd74,8'd77} : s = 422;
	{8'd74,8'd78} : s = 138;
	{8'd74,8'd79} : s = 297;
	{8'd74,8'd80} : s = 294;
	{8'd74,8'd81} : s = 421;
	{8'd74,8'd82} : s = 293;
	{8'd74,8'd83} : s = 419;
	{8'd74,8'd84} : s = 412;
	{8'd74,8'd85} : s = 486;
	{8'd74,8'd86} : s = 24;
	{8'd74,8'd87} : s = 137;
	{8'd74,8'd88} : s = 134;
	{8'd74,8'd89} : s = 291;
	{8'd74,8'd90} : s = 133;
	{8'd74,8'd91} : s = 284;
	{8'd74,8'd92} : s = 282;
	{8'd74,8'd93} : s = 410;
	{8'd74,8'd94} : s = 131;
	{8'd74,8'd95} : s = 281;
	{8'd74,8'd96} : s = 278;
	{8'd74,8'd97} : s = 409;
	{8'd74,8'd98} : s = 277;
	{8'd74,8'd99} : s = 406;
	{8'd74,8'd100} : s = 405;
	{8'd74,8'd101} : s = 485;
	{8'd74,8'd102} : s = 112;
	{8'd74,8'd103} : s = 275;
	{8'd74,8'd104} : s = 270;
	{8'd74,8'd105} : s = 403;
	{8'd74,8'd106} : s = 269;
	{8'd74,8'd107} : s = 398;
	{8'd74,8'd108} : s = 397;
	{8'd74,8'd109} : s = 483;
	{8'd74,8'd110} : s = 267;
	{8'd74,8'd111} : s = 395;
	{8'd74,8'd112} : s = 391;
	{8'd74,8'd113} : s = 476;
	{8'd74,8'd114} : s = 376;
	{8'd74,8'd115} : s = 474;
	{8'd74,8'd116} : s = 473;
	{8'd74,8'd117} : s = 506;
	{8'd74,8'd118} : s = 20;
	{8'd74,8'd119} : s = 104;
	{8'd74,8'd120} : s = 100;
	{8'd74,8'd121} : s = 263;
	{8'd74,8'd122} : s = 98;
	{8'd74,8'd123} : s = 240;
	{8'd74,8'd124} : s = 232;
	{8'd74,8'd125} : s = 372;
	{8'd74,8'd126} : s = 97;
	{8'd74,8'd127} : s = 228;
	{8'd74,8'd128} : s = 226;
	{8'd74,8'd129} : s = 370;
	{8'd74,8'd130} : s = 225;
	{8'd74,8'd131} : s = 369;
	{8'd74,8'd132} : s = 364;
	{8'd74,8'd133} : s = 470;
	{8'd74,8'd134} : s = 88;
	{8'd74,8'd135} : s = 216;
	{8'd74,8'd136} : s = 212;
	{8'd74,8'd137} : s = 362;
	{8'd74,8'd138} : s = 210;
	{8'd74,8'd139} : s = 361;
	{8'd74,8'd140} : s = 358;
	{8'd74,8'd141} : s = 469;
	{8'd74,8'd142} : s = 209;
	{8'd74,8'd143} : s = 357;
	{8'd74,8'd144} : s = 355;
	{8'd74,8'd145} : s = 467;
	{8'd74,8'd146} : s = 348;
	{8'd74,8'd147} : s = 462;
	{8'd74,8'd148} : s = 461;
	{8'd74,8'd149} : s = 505;
	{8'd74,8'd150} : s = 84;
	{8'd74,8'd151} : s = 204;
	{8'd74,8'd152} : s = 202;
	{8'd74,8'd153} : s = 346;
	{8'd74,8'd154} : s = 201;
	{8'd74,8'd155} : s = 345;
	{8'd74,8'd156} : s = 342;
	{8'd74,8'd157} : s = 459;
	{8'd74,8'd158} : s = 198;
	{8'd74,8'd159} : s = 341;
	{8'd74,8'd160} : s = 339;
	{8'd74,8'd161} : s = 455;
	{8'd74,8'd162} : s = 334;
	{8'd74,8'd163} : s = 444;
	{8'd74,8'd164} : s = 442;
	{8'd74,8'd165} : s = 502;
	{8'd74,8'd166} : s = 197;
	{8'd74,8'd167} : s = 333;
	{8'd74,8'd168} : s = 331;
	{8'd74,8'd169} : s = 441;
	{8'd74,8'd170} : s = 327;
	{8'd74,8'd171} : s = 438;
	{8'd74,8'd172} : s = 437;
	{8'd74,8'd173} : s = 501;
	{8'd74,8'd174} : s = 316;
	{8'd74,8'd175} : s = 435;
	{8'd74,8'd176} : s = 430;
	{8'd74,8'd177} : s = 499;
	{8'd74,8'd178} : s = 429;
	{8'd74,8'd179} : s = 494;
	{8'd74,8'd180} : s = 493;
	{8'd74,8'd181} : s = 510;
	{8'd74,8'd182} : s = 1;
	{8'd74,8'd183} : s = 18;
	{8'd74,8'd184} : s = 17;
	{8'd74,8'd185} : s = 82;
	{8'd74,8'd186} : s = 12;
	{8'd74,8'd187} : s = 81;
	{8'd74,8'd188} : s = 76;
	{8'd74,8'd189} : s = 195;
	{8'd74,8'd190} : s = 10;
	{8'd74,8'd191} : s = 74;
	{8'd74,8'd192} : s = 73;
	{8'd74,8'd193} : s = 184;
	{8'd74,8'd194} : s = 70;
	{8'd74,8'd195} : s = 180;
	{8'd74,8'd196} : s = 178;
	{8'd74,8'd197} : s = 314;
	{8'd74,8'd198} : s = 9;
	{8'd74,8'd199} : s = 69;
	{8'd74,8'd200} : s = 67;
	{8'd74,8'd201} : s = 177;
	{8'd74,8'd202} : s = 56;
	{8'd74,8'd203} : s = 172;
	{8'd74,8'd204} : s = 170;
	{8'd74,8'd205} : s = 313;
	{8'd74,8'd206} : s = 52;
	{8'd74,8'd207} : s = 169;
	{8'd74,8'd208} : s = 166;
	{8'd74,8'd209} : s = 310;
	{8'd74,8'd210} : s = 165;
	{8'd74,8'd211} : s = 309;
	{8'd74,8'd212} : s = 307;
	{8'd74,8'd213} : s = 427;
	{8'd74,8'd214} : s = 6;
	{8'd74,8'd215} : s = 50;
	{8'd74,8'd216} : s = 49;
	{8'd74,8'd217} : s = 163;
	{8'd74,8'd218} : s = 44;
	{8'd74,8'd219} : s = 156;
	{8'd74,8'd220} : s = 154;
	{8'd74,8'd221} : s = 302;
	{8'd74,8'd222} : s = 42;
	{8'd74,8'd223} : s = 153;
	{8'd74,8'd224} : s = 150;
	{8'd74,8'd225} : s = 301;
	{8'd74,8'd226} : s = 149;
	{8'd74,8'd227} : s = 299;
	{8'd74,8'd228} : s = 295;
	{8'd74,8'd229} : s = 423;
	{8'd74,8'd230} : s = 41;
	{8'd74,8'd231} : s = 147;
	{8'd74,8'd232} : s = 142;
	{8'd74,8'd233} : s = 286;
	{8'd74,8'd234} : s = 141;
	{8'd74,8'd235} : s = 285;
	{8'd74,8'd236} : s = 283;
	{8'd74,8'd237} : s = 414;
	{8'd74,8'd238} : s = 139;
	{8'd74,8'd239} : s = 279;
	{8'd74,8'd240} : s = 271;
	{8'd74,8'd241} : s = 413;
	{8'd74,8'd242} : s = 248;
	{8'd74,8'd243} : s = 411;
	{8'd74,8'd244} : s = 407;
	{8'd74,8'd245} : s = 491;
	{8'd74,8'd246} : s = 5;
	{8'd74,8'd247} : s = 38;
	{8'd74,8'd248} : s = 37;
	{8'd74,8'd249} : s = 135;
	{8'd74,8'd250} : s = 35;
	{8'd74,8'd251} : s = 120;
	{8'd74,8'd252} : s = 116;
	{8'd74,8'd253} : s = 244;
	{8'd74,8'd254} : s = 28;
	{8'd74,8'd255} : s = 114;
	{8'd75,8'd0} : s = 394;
	{8'd75,8'd1} : s = 262;
	{8'd75,8'd2} : s = 393;
	{8'd75,8'd3} : s = 390;
	{8'd75,8'd4} : s = 468;
	{8'd75,8'd5} : s = 66;
	{8'd75,8'd6} : s = 261;
	{8'd75,8'd7} : s = 259;
	{8'd75,8'd8} : s = 389;
	{8'd75,8'd9} : s = 224;
	{8'd75,8'd10} : s = 387;
	{8'd75,8'd11} : s = 368;
	{8'd75,8'd12} : s = 466;
	{8'd75,8'd13} : s = 208;
	{8'd75,8'd14} : s = 360;
	{8'd75,8'd15} : s = 356;
	{8'd75,8'd16} : s = 465;
	{8'd75,8'd17} : s = 354;
	{8'd75,8'd18} : s = 460;
	{8'd75,8'd19} : s = 458;
	{8'd75,8'd20} : s = 500;
	{8'd75,8'd21} : s = 65;
	{8'd75,8'd22} : s = 200;
	{8'd75,8'd23} : s = 196;
	{8'd75,8'd24} : s = 353;
	{8'd75,8'd25} : s = 194;
	{8'd75,8'd26} : s = 344;
	{8'd75,8'd27} : s = 340;
	{8'd75,8'd28} : s = 457;
	{8'd75,8'd29} : s = 193;
	{8'd75,8'd30} : s = 338;
	{8'd75,8'd31} : s = 337;
	{8'd75,8'd32} : s = 454;
	{8'd75,8'd33} : s = 332;
	{8'd75,8'd34} : s = 453;
	{8'd75,8'd35} : s = 451;
	{8'd75,8'd36} : s = 498;
	{8'd75,8'd37} : s = 176;
	{8'd75,8'd38} : s = 330;
	{8'd75,8'd39} : s = 329;
	{8'd75,8'd40} : s = 440;
	{8'd75,8'd41} : s = 326;
	{8'd75,8'd42} : s = 436;
	{8'd75,8'd43} : s = 434;
	{8'd75,8'd44} : s = 497;
	{8'd75,8'd45} : s = 325;
	{8'd75,8'd46} : s = 433;
	{8'd75,8'd47} : s = 428;
	{8'd75,8'd48} : s = 492;
	{8'd75,8'd49} : s = 426;
	{8'd75,8'd50} : s = 490;
	{8'd75,8'd51} : s = 489;
	{8'd75,8'd52} : s = 508;
	{8'd75,8'd53} : s = 2;
	{8'd75,8'd54} : s = 48;
	{8'd75,8'd55} : s = 40;
	{8'd75,8'd56} : s = 168;
	{8'd75,8'd57} : s = 36;
	{8'd75,8'd58} : s = 164;
	{8'd75,8'd59} : s = 162;
	{8'd75,8'd60} : s = 323;
	{8'd75,8'd61} : s = 34;
	{8'd75,8'd62} : s = 161;
	{8'd75,8'd63} : s = 152;
	{8'd75,8'd64} : s = 312;
	{8'd75,8'd65} : s = 148;
	{8'd75,8'd66} : s = 308;
	{8'd75,8'd67} : s = 306;
	{8'd75,8'd68} : s = 425;
	{8'd75,8'd69} : s = 33;
	{8'd75,8'd70} : s = 146;
	{8'd75,8'd71} : s = 145;
	{8'd75,8'd72} : s = 305;
	{8'd75,8'd73} : s = 140;
	{8'd75,8'd74} : s = 300;
	{8'd75,8'd75} : s = 298;
	{8'd75,8'd76} : s = 422;
	{8'd75,8'd77} : s = 138;
	{8'd75,8'd78} : s = 297;
	{8'd75,8'd79} : s = 294;
	{8'd75,8'd80} : s = 421;
	{8'd75,8'd81} : s = 293;
	{8'd75,8'd82} : s = 419;
	{8'd75,8'd83} : s = 412;
	{8'd75,8'd84} : s = 486;
	{8'd75,8'd85} : s = 24;
	{8'd75,8'd86} : s = 137;
	{8'd75,8'd87} : s = 134;
	{8'd75,8'd88} : s = 291;
	{8'd75,8'd89} : s = 133;
	{8'd75,8'd90} : s = 284;
	{8'd75,8'd91} : s = 282;
	{8'd75,8'd92} : s = 410;
	{8'd75,8'd93} : s = 131;
	{8'd75,8'd94} : s = 281;
	{8'd75,8'd95} : s = 278;
	{8'd75,8'd96} : s = 409;
	{8'd75,8'd97} : s = 277;
	{8'd75,8'd98} : s = 406;
	{8'd75,8'd99} : s = 405;
	{8'd75,8'd100} : s = 485;
	{8'd75,8'd101} : s = 112;
	{8'd75,8'd102} : s = 275;
	{8'd75,8'd103} : s = 270;
	{8'd75,8'd104} : s = 403;
	{8'd75,8'd105} : s = 269;
	{8'd75,8'd106} : s = 398;
	{8'd75,8'd107} : s = 397;
	{8'd75,8'd108} : s = 483;
	{8'd75,8'd109} : s = 267;
	{8'd75,8'd110} : s = 395;
	{8'd75,8'd111} : s = 391;
	{8'd75,8'd112} : s = 476;
	{8'd75,8'd113} : s = 376;
	{8'd75,8'd114} : s = 474;
	{8'd75,8'd115} : s = 473;
	{8'd75,8'd116} : s = 506;
	{8'd75,8'd117} : s = 20;
	{8'd75,8'd118} : s = 104;
	{8'd75,8'd119} : s = 100;
	{8'd75,8'd120} : s = 263;
	{8'd75,8'd121} : s = 98;
	{8'd75,8'd122} : s = 240;
	{8'd75,8'd123} : s = 232;
	{8'd75,8'd124} : s = 372;
	{8'd75,8'd125} : s = 97;
	{8'd75,8'd126} : s = 228;
	{8'd75,8'd127} : s = 226;
	{8'd75,8'd128} : s = 370;
	{8'd75,8'd129} : s = 225;
	{8'd75,8'd130} : s = 369;
	{8'd75,8'd131} : s = 364;
	{8'd75,8'd132} : s = 470;
	{8'd75,8'd133} : s = 88;
	{8'd75,8'd134} : s = 216;
	{8'd75,8'd135} : s = 212;
	{8'd75,8'd136} : s = 362;
	{8'd75,8'd137} : s = 210;
	{8'd75,8'd138} : s = 361;
	{8'd75,8'd139} : s = 358;
	{8'd75,8'd140} : s = 469;
	{8'd75,8'd141} : s = 209;
	{8'd75,8'd142} : s = 357;
	{8'd75,8'd143} : s = 355;
	{8'd75,8'd144} : s = 467;
	{8'd75,8'd145} : s = 348;
	{8'd75,8'd146} : s = 462;
	{8'd75,8'd147} : s = 461;
	{8'd75,8'd148} : s = 505;
	{8'd75,8'd149} : s = 84;
	{8'd75,8'd150} : s = 204;
	{8'd75,8'd151} : s = 202;
	{8'd75,8'd152} : s = 346;
	{8'd75,8'd153} : s = 201;
	{8'd75,8'd154} : s = 345;
	{8'd75,8'd155} : s = 342;
	{8'd75,8'd156} : s = 459;
	{8'd75,8'd157} : s = 198;
	{8'd75,8'd158} : s = 341;
	{8'd75,8'd159} : s = 339;
	{8'd75,8'd160} : s = 455;
	{8'd75,8'd161} : s = 334;
	{8'd75,8'd162} : s = 444;
	{8'd75,8'd163} : s = 442;
	{8'd75,8'd164} : s = 502;
	{8'd75,8'd165} : s = 197;
	{8'd75,8'd166} : s = 333;
	{8'd75,8'd167} : s = 331;
	{8'd75,8'd168} : s = 441;
	{8'd75,8'd169} : s = 327;
	{8'd75,8'd170} : s = 438;
	{8'd75,8'd171} : s = 437;
	{8'd75,8'd172} : s = 501;
	{8'd75,8'd173} : s = 316;
	{8'd75,8'd174} : s = 435;
	{8'd75,8'd175} : s = 430;
	{8'd75,8'd176} : s = 499;
	{8'd75,8'd177} : s = 429;
	{8'd75,8'd178} : s = 494;
	{8'd75,8'd179} : s = 493;
	{8'd75,8'd180} : s = 510;
	{8'd75,8'd181} : s = 1;
	{8'd75,8'd182} : s = 18;
	{8'd75,8'd183} : s = 17;
	{8'd75,8'd184} : s = 82;
	{8'd75,8'd185} : s = 12;
	{8'd75,8'd186} : s = 81;
	{8'd75,8'd187} : s = 76;
	{8'd75,8'd188} : s = 195;
	{8'd75,8'd189} : s = 10;
	{8'd75,8'd190} : s = 74;
	{8'd75,8'd191} : s = 73;
	{8'd75,8'd192} : s = 184;
	{8'd75,8'd193} : s = 70;
	{8'd75,8'd194} : s = 180;
	{8'd75,8'd195} : s = 178;
	{8'd75,8'd196} : s = 314;
	{8'd75,8'd197} : s = 9;
	{8'd75,8'd198} : s = 69;
	{8'd75,8'd199} : s = 67;
	{8'd75,8'd200} : s = 177;
	{8'd75,8'd201} : s = 56;
	{8'd75,8'd202} : s = 172;
	{8'd75,8'd203} : s = 170;
	{8'd75,8'd204} : s = 313;
	{8'd75,8'd205} : s = 52;
	{8'd75,8'd206} : s = 169;
	{8'd75,8'd207} : s = 166;
	{8'd75,8'd208} : s = 310;
	{8'd75,8'd209} : s = 165;
	{8'd75,8'd210} : s = 309;
	{8'd75,8'd211} : s = 307;
	{8'd75,8'd212} : s = 427;
	{8'd75,8'd213} : s = 6;
	{8'd75,8'd214} : s = 50;
	{8'd75,8'd215} : s = 49;
	{8'd75,8'd216} : s = 163;
	{8'd75,8'd217} : s = 44;
	{8'd75,8'd218} : s = 156;
	{8'd75,8'd219} : s = 154;
	{8'd75,8'd220} : s = 302;
	{8'd75,8'd221} : s = 42;
	{8'd75,8'd222} : s = 153;
	{8'd75,8'd223} : s = 150;
	{8'd75,8'd224} : s = 301;
	{8'd75,8'd225} : s = 149;
	{8'd75,8'd226} : s = 299;
	{8'd75,8'd227} : s = 295;
	{8'd75,8'd228} : s = 423;
	{8'd75,8'd229} : s = 41;
	{8'd75,8'd230} : s = 147;
	{8'd75,8'd231} : s = 142;
	{8'd75,8'd232} : s = 286;
	{8'd75,8'd233} : s = 141;
	{8'd75,8'd234} : s = 285;
	{8'd75,8'd235} : s = 283;
	{8'd75,8'd236} : s = 414;
	{8'd75,8'd237} : s = 139;
	{8'd75,8'd238} : s = 279;
	{8'd75,8'd239} : s = 271;
	{8'd75,8'd240} : s = 413;
	{8'd75,8'd241} : s = 248;
	{8'd75,8'd242} : s = 411;
	{8'd75,8'd243} : s = 407;
	{8'd75,8'd244} : s = 491;
	{8'd75,8'd245} : s = 5;
	{8'd75,8'd246} : s = 38;
	{8'd75,8'd247} : s = 37;
	{8'd75,8'd248} : s = 135;
	{8'd75,8'd249} : s = 35;
	{8'd75,8'd250} : s = 120;
	{8'd75,8'd251} : s = 116;
	{8'd75,8'd252} : s = 244;
	{8'd75,8'd253} : s = 28;
	{8'd75,8'd254} : s = 114;
	{8'd75,8'd255} : s = 113;
	{8'd76,8'd0} : s = 262;
	{8'd76,8'd1} : s = 393;
	{8'd76,8'd2} : s = 390;
	{8'd76,8'd3} : s = 468;
	{8'd76,8'd4} : s = 66;
	{8'd76,8'd5} : s = 261;
	{8'd76,8'd6} : s = 259;
	{8'd76,8'd7} : s = 389;
	{8'd76,8'd8} : s = 224;
	{8'd76,8'd9} : s = 387;
	{8'd76,8'd10} : s = 368;
	{8'd76,8'd11} : s = 466;
	{8'd76,8'd12} : s = 208;
	{8'd76,8'd13} : s = 360;
	{8'd76,8'd14} : s = 356;
	{8'd76,8'd15} : s = 465;
	{8'd76,8'd16} : s = 354;
	{8'd76,8'd17} : s = 460;
	{8'd76,8'd18} : s = 458;
	{8'd76,8'd19} : s = 500;
	{8'd76,8'd20} : s = 65;
	{8'd76,8'd21} : s = 200;
	{8'd76,8'd22} : s = 196;
	{8'd76,8'd23} : s = 353;
	{8'd76,8'd24} : s = 194;
	{8'd76,8'd25} : s = 344;
	{8'd76,8'd26} : s = 340;
	{8'd76,8'd27} : s = 457;
	{8'd76,8'd28} : s = 193;
	{8'd76,8'd29} : s = 338;
	{8'd76,8'd30} : s = 337;
	{8'd76,8'd31} : s = 454;
	{8'd76,8'd32} : s = 332;
	{8'd76,8'd33} : s = 453;
	{8'd76,8'd34} : s = 451;
	{8'd76,8'd35} : s = 498;
	{8'd76,8'd36} : s = 176;
	{8'd76,8'd37} : s = 330;
	{8'd76,8'd38} : s = 329;
	{8'd76,8'd39} : s = 440;
	{8'd76,8'd40} : s = 326;
	{8'd76,8'd41} : s = 436;
	{8'd76,8'd42} : s = 434;
	{8'd76,8'd43} : s = 497;
	{8'd76,8'd44} : s = 325;
	{8'd76,8'd45} : s = 433;
	{8'd76,8'd46} : s = 428;
	{8'd76,8'd47} : s = 492;
	{8'd76,8'd48} : s = 426;
	{8'd76,8'd49} : s = 490;
	{8'd76,8'd50} : s = 489;
	{8'd76,8'd51} : s = 508;
	{8'd76,8'd52} : s = 2;
	{8'd76,8'd53} : s = 48;
	{8'd76,8'd54} : s = 40;
	{8'd76,8'd55} : s = 168;
	{8'd76,8'd56} : s = 36;
	{8'd76,8'd57} : s = 164;
	{8'd76,8'd58} : s = 162;
	{8'd76,8'd59} : s = 323;
	{8'd76,8'd60} : s = 34;
	{8'd76,8'd61} : s = 161;
	{8'd76,8'd62} : s = 152;
	{8'd76,8'd63} : s = 312;
	{8'd76,8'd64} : s = 148;
	{8'd76,8'd65} : s = 308;
	{8'd76,8'd66} : s = 306;
	{8'd76,8'd67} : s = 425;
	{8'd76,8'd68} : s = 33;
	{8'd76,8'd69} : s = 146;
	{8'd76,8'd70} : s = 145;
	{8'd76,8'd71} : s = 305;
	{8'd76,8'd72} : s = 140;
	{8'd76,8'd73} : s = 300;
	{8'd76,8'd74} : s = 298;
	{8'd76,8'd75} : s = 422;
	{8'd76,8'd76} : s = 138;
	{8'd76,8'd77} : s = 297;
	{8'd76,8'd78} : s = 294;
	{8'd76,8'd79} : s = 421;
	{8'd76,8'd80} : s = 293;
	{8'd76,8'd81} : s = 419;
	{8'd76,8'd82} : s = 412;
	{8'd76,8'd83} : s = 486;
	{8'd76,8'd84} : s = 24;
	{8'd76,8'd85} : s = 137;
	{8'd76,8'd86} : s = 134;
	{8'd76,8'd87} : s = 291;
	{8'd76,8'd88} : s = 133;
	{8'd76,8'd89} : s = 284;
	{8'd76,8'd90} : s = 282;
	{8'd76,8'd91} : s = 410;
	{8'd76,8'd92} : s = 131;
	{8'd76,8'd93} : s = 281;
	{8'd76,8'd94} : s = 278;
	{8'd76,8'd95} : s = 409;
	{8'd76,8'd96} : s = 277;
	{8'd76,8'd97} : s = 406;
	{8'd76,8'd98} : s = 405;
	{8'd76,8'd99} : s = 485;
	{8'd76,8'd100} : s = 112;
	{8'd76,8'd101} : s = 275;
	{8'd76,8'd102} : s = 270;
	{8'd76,8'd103} : s = 403;
	{8'd76,8'd104} : s = 269;
	{8'd76,8'd105} : s = 398;
	{8'd76,8'd106} : s = 397;
	{8'd76,8'd107} : s = 483;
	{8'd76,8'd108} : s = 267;
	{8'd76,8'd109} : s = 395;
	{8'd76,8'd110} : s = 391;
	{8'd76,8'd111} : s = 476;
	{8'd76,8'd112} : s = 376;
	{8'd76,8'd113} : s = 474;
	{8'd76,8'd114} : s = 473;
	{8'd76,8'd115} : s = 506;
	{8'd76,8'd116} : s = 20;
	{8'd76,8'd117} : s = 104;
	{8'd76,8'd118} : s = 100;
	{8'd76,8'd119} : s = 263;
	{8'd76,8'd120} : s = 98;
	{8'd76,8'd121} : s = 240;
	{8'd76,8'd122} : s = 232;
	{8'd76,8'd123} : s = 372;
	{8'd76,8'd124} : s = 97;
	{8'd76,8'd125} : s = 228;
	{8'd76,8'd126} : s = 226;
	{8'd76,8'd127} : s = 370;
	{8'd76,8'd128} : s = 225;
	{8'd76,8'd129} : s = 369;
	{8'd76,8'd130} : s = 364;
	{8'd76,8'd131} : s = 470;
	{8'd76,8'd132} : s = 88;
	{8'd76,8'd133} : s = 216;
	{8'd76,8'd134} : s = 212;
	{8'd76,8'd135} : s = 362;
	{8'd76,8'd136} : s = 210;
	{8'd76,8'd137} : s = 361;
	{8'd76,8'd138} : s = 358;
	{8'd76,8'd139} : s = 469;
	{8'd76,8'd140} : s = 209;
	{8'd76,8'd141} : s = 357;
	{8'd76,8'd142} : s = 355;
	{8'd76,8'd143} : s = 467;
	{8'd76,8'd144} : s = 348;
	{8'd76,8'd145} : s = 462;
	{8'd76,8'd146} : s = 461;
	{8'd76,8'd147} : s = 505;
	{8'd76,8'd148} : s = 84;
	{8'd76,8'd149} : s = 204;
	{8'd76,8'd150} : s = 202;
	{8'd76,8'd151} : s = 346;
	{8'd76,8'd152} : s = 201;
	{8'd76,8'd153} : s = 345;
	{8'd76,8'd154} : s = 342;
	{8'd76,8'd155} : s = 459;
	{8'd76,8'd156} : s = 198;
	{8'd76,8'd157} : s = 341;
	{8'd76,8'd158} : s = 339;
	{8'd76,8'd159} : s = 455;
	{8'd76,8'd160} : s = 334;
	{8'd76,8'd161} : s = 444;
	{8'd76,8'd162} : s = 442;
	{8'd76,8'd163} : s = 502;
	{8'd76,8'd164} : s = 197;
	{8'd76,8'd165} : s = 333;
	{8'd76,8'd166} : s = 331;
	{8'd76,8'd167} : s = 441;
	{8'd76,8'd168} : s = 327;
	{8'd76,8'd169} : s = 438;
	{8'd76,8'd170} : s = 437;
	{8'd76,8'd171} : s = 501;
	{8'd76,8'd172} : s = 316;
	{8'd76,8'd173} : s = 435;
	{8'd76,8'd174} : s = 430;
	{8'd76,8'd175} : s = 499;
	{8'd76,8'd176} : s = 429;
	{8'd76,8'd177} : s = 494;
	{8'd76,8'd178} : s = 493;
	{8'd76,8'd179} : s = 510;
	{8'd76,8'd180} : s = 1;
	{8'd76,8'd181} : s = 18;
	{8'd76,8'd182} : s = 17;
	{8'd76,8'd183} : s = 82;
	{8'd76,8'd184} : s = 12;
	{8'd76,8'd185} : s = 81;
	{8'd76,8'd186} : s = 76;
	{8'd76,8'd187} : s = 195;
	{8'd76,8'd188} : s = 10;
	{8'd76,8'd189} : s = 74;
	{8'd76,8'd190} : s = 73;
	{8'd76,8'd191} : s = 184;
	{8'd76,8'd192} : s = 70;
	{8'd76,8'd193} : s = 180;
	{8'd76,8'd194} : s = 178;
	{8'd76,8'd195} : s = 314;
	{8'd76,8'd196} : s = 9;
	{8'd76,8'd197} : s = 69;
	{8'd76,8'd198} : s = 67;
	{8'd76,8'd199} : s = 177;
	{8'd76,8'd200} : s = 56;
	{8'd76,8'd201} : s = 172;
	{8'd76,8'd202} : s = 170;
	{8'd76,8'd203} : s = 313;
	{8'd76,8'd204} : s = 52;
	{8'd76,8'd205} : s = 169;
	{8'd76,8'd206} : s = 166;
	{8'd76,8'd207} : s = 310;
	{8'd76,8'd208} : s = 165;
	{8'd76,8'd209} : s = 309;
	{8'd76,8'd210} : s = 307;
	{8'd76,8'd211} : s = 427;
	{8'd76,8'd212} : s = 6;
	{8'd76,8'd213} : s = 50;
	{8'd76,8'd214} : s = 49;
	{8'd76,8'd215} : s = 163;
	{8'd76,8'd216} : s = 44;
	{8'd76,8'd217} : s = 156;
	{8'd76,8'd218} : s = 154;
	{8'd76,8'd219} : s = 302;
	{8'd76,8'd220} : s = 42;
	{8'd76,8'd221} : s = 153;
	{8'd76,8'd222} : s = 150;
	{8'd76,8'd223} : s = 301;
	{8'd76,8'd224} : s = 149;
	{8'd76,8'd225} : s = 299;
	{8'd76,8'd226} : s = 295;
	{8'd76,8'd227} : s = 423;
	{8'd76,8'd228} : s = 41;
	{8'd76,8'd229} : s = 147;
	{8'd76,8'd230} : s = 142;
	{8'd76,8'd231} : s = 286;
	{8'd76,8'd232} : s = 141;
	{8'd76,8'd233} : s = 285;
	{8'd76,8'd234} : s = 283;
	{8'd76,8'd235} : s = 414;
	{8'd76,8'd236} : s = 139;
	{8'd76,8'd237} : s = 279;
	{8'd76,8'd238} : s = 271;
	{8'd76,8'd239} : s = 413;
	{8'd76,8'd240} : s = 248;
	{8'd76,8'd241} : s = 411;
	{8'd76,8'd242} : s = 407;
	{8'd76,8'd243} : s = 491;
	{8'd76,8'd244} : s = 5;
	{8'd76,8'd245} : s = 38;
	{8'd76,8'd246} : s = 37;
	{8'd76,8'd247} : s = 135;
	{8'd76,8'd248} : s = 35;
	{8'd76,8'd249} : s = 120;
	{8'd76,8'd250} : s = 116;
	{8'd76,8'd251} : s = 244;
	{8'd76,8'd252} : s = 28;
	{8'd76,8'd253} : s = 114;
	{8'd76,8'd254} : s = 113;
	{8'd76,8'd255} : s = 242;
	{8'd77,8'd0} : s = 393;
	{8'd77,8'd1} : s = 390;
	{8'd77,8'd2} : s = 468;
	{8'd77,8'd3} : s = 66;
	{8'd77,8'd4} : s = 261;
	{8'd77,8'd5} : s = 259;
	{8'd77,8'd6} : s = 389;
	{8'd77,8'd7} : s = 224;
	{8'd77,8'd8} : s = 387;
	{8'd77,8'd9} : s = 368;
	{8'd77,8'd10} : s = 466;
	{8'd77,8'd11} : s = 208;
	{8'd77,8'd12} : s = 360;
	{8'd77,8'd13} : s = 356;
	{8'd77,8'd14} : s = 465;
	{8'd77,8'd15} : s = 354;
	{8'd77,8'd16} : s = 460;
	{8'd77,8'd17} : s = 458;
	{8'd77,8'd18} : s = 500;
	{8'd77,8'd19} : s = 65;
	{8'd77,8'd20} : s = 200;
	{8'd77,8'd21} : s = 196;
	{8'd77,8'd22} : s = 353;
	{8'd77,8'd23} : s = 194;
	{8'd77,8'd24} : s = 344;
	{8'd77,8'd25} : s = 340;
	{8'd77,8'd26} : s = 457;
	{8'd77,8'd27} : s = 193;
	{8'd77,8'd28} : s = 338;
	{8'd77,8'd29} : s = 337;
	{8'd77,8'd30} : s = 454;
	{8'd77,8'd31} : s = 332;
	{8'd77,8'd32} : s = 453;
	{8'd77,8'd33} : s = 451;
	{8'd77,8'd34} : s = 498;
	{8'd77,8'd35} : s = 176;
	{8'd77,8'd36} : s = 330;
	{8'd77,8'd37} : s = 329;
	{8'd77,8'd38} : s = 440;
	{8'd77,8'd39} : s = 326;
	{8'd77,8'd40} : s = 436;
	{8'd77,8'd41} : s = 434;
	{8'd77,8'd42} : s = 497;
	{8'd77,8'd43} : s = 325;
	{8'd77,8'd44} : s = 433;
	{8'd77,8'd45} : s = 428;
	{8'd77,8'd46} : s = 492;
	{8'd77,8'd47} : s = 426;
	{8'd77,8'd48} : s = 490;
	{8'd77,8'd49} : s = 489;
	{8'd77,8'd50} : s = 508;
	{8'd77,8'd51} : s = 2;
	{8'd77,8'd52} : s = 48;
	{8'd77,8'd53} : s = 40;
	{8'd77,8'd54} : s = 168;
	{8'd77,8'd55} : s = 36;
	{8'd77,8'd56} : s = 164;
	{8'd77,8'd57} : s = 162;
	{8'd77,8'd58} : s = 323;
	{8'd77,8'd59} : s = 34;
	{8'd77,8'd60} : s = 161;
	{8'd77,8'd61} : s = 152;
	{8'd77,8'd62} : s = 312;
	{8'd77,8'd63} : s = 148;
	{8'd77,8'd64} : s = 308;
	{8'd77,8'd65} : s = 306;
	{8'd77,8'd66} : s = 425;
	{8'd77,8'd67} : s = 33;
	{8'd77,8'd68} : s = 146;
	{8'd77,8'd69} : s = 145;
	{8'd77,8'd70} : s = 305;
	{8'd77,8'd71} : s = 140;
	{8'd77,8'd72} : s = 300;
	{8'd77,8'd73} : s = 298;
	{8'd77,8'd74} : s = 422;
	{8'd77,8'd75} : s = 138;
	{8'd77,8'd76} : s = 297;
	{8'd77,8'd77} : s = 294;
	{8'd77,8'd78} : s = 421;
	{8'd77,8'd79} : s = 293;
	{8'd77,8'd80} : s = 419;
	{8'd77,8'd81} : s = 412;
	{8'd77,8'd82} : s = 486;
	{8'd77,8'd83} : s = 24;
	{8'd77,8'd84} : s = 137;
	{8'd77,8'd85} : s = 134;
	{8'd77,8'd86} : s = 291;
	{8'd77,8'd87} : s = 133;
	{8'd77,8'd88} : s = 284;
	{8'd77,8'd89} : s = 282;
	{8'd77,8'd90} : s = 410;
	{8'd77,8'd91} : s = 131;
	{8'd77,8'd92} : s = 281;
	{8'd77,8'd93} : s = 278;
	{8'd77,8'd94} : s = 409;
	{8'd77,8'd95} : s = 277;
	{8'd77,8'd96} : s = 406;
	{8'd77,8'd97} : s = 405;
	{8'd77,8'd98} : s = 485;
	{8'd77,8'd99} : s = 112;
	{8'd77,8'd100} : s = 275;
	{8'd77,8'd101} : s = 270;
	{8'd77,8'd102} : s = 403;
	{8'd77,8'd103} : s = 269;
	{8'd77,8'd104} : s = 398;
	{8'd77,8'd105} : s = 397;
	{8'd77,8'd106} : s = 483;
	{8'd77,8'd107} : s = 267;
	{8'd77,8'd108} : s = 395;
	{8'd77,8'd109} : s = 391;
	{8'd77,8'd110} : s = 476;
	{8'd77,8'd111} : s = 376;
	{8'd77,8'd112} : s = 474;
	{8'd77,8'd113} : s = 473;
	{8'd77,8'd114} : s = 506;
	{8'd77,8'd115} : s = 20;
	{8'd77,8'd116} : s = 104;
	{8'd77,8'd117} : s = 100;
	{8'd77,8'd118} : s = 263;
	{8'd77,8'd119} : s = 98;
	{8'd77,8'd120} : s = 240;
	{8'd77,8'd121} : s = 232;
	{8'd77,8'd122} : s = 372;
	{8'd77,8'd123} : s = 97;
	{8'd77,8'd124} : s = 228;
	{8'd77,8'd125} : s = 226;
	{8'd77,8'd126} : s = 370;
	{8'd77,8'd127} : s = 225;
	{8'd77,8'd128} : s = 369;
	{8'd77,8'd129} : s = 364;
	{8'd77,8'd130} : s = 470;
	{8'd77,8'd131} : s = 88;
	{8'd77,8'd132} : s = 216;
	{8'd77,8'd133} : s = 212;
	{8'd77,8'd134} : s = 362;
	{8'd77,8'd135} : s = 210;
	{8'd77,8'd136} : s = 361;
	{8'd77,8'd137} : s = 358;
	{8'd77,8'd138} : s = 469;
	{8'd77,8'd139} : s = 209;
	{8'd77,8'd140} : s = 357;
	{8'd77,8'd141} : s = 355;
	{8'd77,8'd142} : s = 467;
	{8'd77,8'd143} : s = 348;
	{8'd77,8'd144} : s = 462;
	{8'd77,8'd145} : s = 461;
	{8'd77,8'd146} : s = 505;
	{8'd77,8'd147} : s = 84;
	{8'd77,8'd148} : s = 204;
	{8'd77,8'd149} : s = 202;
	{8'd77,8'd150} : s = 346;
	{8'd77,8'd151} : s = 201;
	{8'd77,8'd152} : s = 345;
	{8'd77,8'd153} : s = 342;
	{8'd77,8'd154} : s = 459;
	{8'd77,8'd155} : s = 198;
	{8'd77,8'd156} : s = 341;
	{8'd77,8'd157} : s = 339;
	{8'd77,8'd158} : s = 455;
	{8'd77,8'd159} : s = 334;
	{8'd77,8'd160} : s = 444;
	{8'd77,8'd161} : s = 442;
	{8'd77,8'd162} : s = 502;
	{8'd77,8'd163} : s = 197;
	{8'd77,8'd164} : s = 333;
	{8'd77,8'd165} : s = 331;
	{8'd77,8'd166} : s = 441;
	{8'd77,8'd167} : s = 327;
	{8'd77,8'd168} : s = 438;
	{8'd77,8'd169} : s = 437;
	{8'd77,8'd170} : s = 501;
	{8'd77,8'd171} : s = 316;
	{8'd77,8'd172} : s = 435;
	{8'd77,8'd173} : s = 430;
	{8'd77,8'd174} : s = 499;
	{8'd77,8'd175} : s = 429;
	{8'd77,8'd176} : s = 494;
	{8'd77,8'd177} : s = 493;
	{8'd77,8'd178} : s = 510;
	{8'd77,8'd179} : s = 1;
	{8'd77,8'd180} : s = 18;
	{8'd77,8'd181} : s = 17;
	{8'd77,8'd182} : s = 82;
	{8'd77,8'd183} : s = 12;
	{8'd77,8'd184} : s = 81;
	{8'd77,8'd185} : s = 76;
	{8'd77,8'd186} : s = 195;
	{8'd77,8'd187} : s = 10;
	{8'd77,8'd188} : s = 74;
	{8'd77,8'd189} : s = 73;
	{8'd77,8'd190} : s = 184;
	{8'd77,8'd191} : s = 70;
	{8'd77,8'd192} : s = 180;
	{8'd77,8'd193} : s = 178;
	{8'd77,8'd194} : s = 314;
	{8'd77,8'd195} : s = 9;
	{8'd77,8'd196} : s = 69;
	{8'd77,8'd197} : s = 67;
	{8'd77,8'd198} : s = 177;
	{8'd77,8'd199} : s = 56;
	{8'd77,8'd200} : s = 172;
	{8'd77,8'd201} : s = 170;
	{8'd77,8'd202} : s = 313;
	{8'd77,8'd203} : s = 52;
	{8'd77,8'd204} : s = 169;
	{8'd77,8'd205} : s = 166;
	{8'd77,8'd206} : s = 310;
	{8'd77,8'd207} : s = 165;
	{8'd77,8'd208} : s = 309;
	{8'd77,8'd209} : s = 307;
	{8'd77,8'd210} : s = 427;
	{8'd77,8'd211} : s = 6;
	{8'd77,8'd212} : s = 50;
	{8'd77,8'd213} : s = 49;
	{8'd77,8'd214} : s = 163;
	{8'd77,8'd215} : s = 44;
	{8'd77,8'd216} : s = 156;
	{8'd77,8'd217} : s = 154;
	{8'd77,8'd218} : s = 302;
	{8'd77,8'd219} : s = 42;
	{8'd77,8'd220} : s = 153;
	{8'd77,8'd221} : s = 150;
	{8'd77,8'd222} : s = 301;
	{8'd77,8'd223} : s = 149;
	{8'd77,8'd224} : s = 299;
	{8'd77,8'd225} : s = 295;
	{8'd77,8'd226} : s = 423;
	{8'd77,8'd227} : s = 41;
	{8'd77,8'd228} : s = 147;
	{8'd77,8'd229} : s = 142;
	{8'd77,8'd230} : s = 286;
	{8'd77,8'd231} : s = 141;
	{8'd77,8'd232} : s = 285;
	{8'd77,8'd233} : s = 283;
	{8'd77,8'd234} : s = 414;
	{8'd77,8'd235} : s = 139;
	{8'd77,8'd236} : s = 279;
	{8'd77,8'd237} : s = 271;
	{8'd77,8'd238} : s = 413;
	{8'd77,8'd239} : s = 248;
	{8'd77,8'd240} : s = 411;
	{8'd77,8'd241} : s = 407;
	{8'd77,8'd242} : s = 491;
	{8'd77,8'd243} : s = 5;
	{8'd77,8'd244} : s = 38;
	{8'd77,8'd245} : s = 37;
	{8'd77,8'd246} : s = 135;
	{8'd77,8'd247} : s = 35;
	{8'd77,8'd248} : s = 120;
	{8'd77,8'd249} : s = 116;
	{8'd77,8'd250} : s = 244;
	{8'd77,8'd251} : s = 28;
	{8'd77,8'd252} : s = 114;
	{8'd77,8'd253} : s = 113;
	{8'd77,8'd254} : s = 242;
	{8'd77,8'd255} : s = 108;
	{8'd78,8'd0} : s = 390;
	{8'd78,8'd1} : s = 468;
	{8'd78,8'd2} : s = 66;
	{8'd78,8'd3} : s = 261;
	{8'd78,8'd4} : s = 259;
	{8'd78,8'd5} : s = 389;
	{8'd78,8'd6} : s = 224;
	{8'd78,8'd7} : s = 387;
	{8'd78,8'd8} : s = 368;
	{8'd78,8'd9} : s = 466;
	{8'd78,8'd10} : s = 208;
	{8'd78,8'd11} : s = 360;
	{8'd78,8'd12} : s = 356;
	{8'd78,8'd13} : s = 465;
	{8'd78,8'd14} : s = 354;
	{8'd78,8'd15} : s = 460;
	{8'd78,8'd16} : s = 458;
	{8'd78,8'd17} : s = 500;
	{8'd78,8'd18} : s = 65;
	{8'd78,8'd19} : s = 200;
	{8'd78,8'd20} : s = 196;
	{8'd78,8'd21} : s = 353;
	{8'd78,8'd22} : s = 194;
	{8'd78,8'd23} : s = 344;
	{8'd78,8'd24} : s = 340;
	{8'd78,8'd25} : s = 457;
	{8'd78,8'd26} : s = 193;
	{8'd78,8'd27} : s = 338;
	{8'd78,8'd28} : s = 337;
	{8'd78,8'd29} : s = 454;
	{8'd78,8'd30} : s = 332;
	{8'd78,8'd31} : s = 453;
	{8'd78,8'd32} : s = 451;
	{8'd78,8'd33} : s = 498;
	{8'd78,8'd34} : s = 176;
	{8'd78,8'd35} : s = 330;
	{8'd78,8'd36} : s = 329;
	{8'd78,8'd37} : s = 440;
	{8'd78,8'd38} : s = 326;
	{8'd78,8'd39} : s = 436;
	{8'd78,8'd40} : s = 434;
	{8'd78,8'd41} : s = 497;
	{8'd78,8'd42} : s = 325;
	{8'd78,8'd43} : s = 433;
	{8'd78,8'd44} : s = 428;
	{8'd78,8'd45} : s = 492;
	{8'd78,8'd46} : s = 426;
	{8'd78,8'd47} : s = 490;
	{8'd78,8'd48} : s = 489;
	{8'd78,8'd49} : s = 508;
	{8'd78,8'd50} : s = 2;
	{8'd78,8'd51} : s = 48;
	{8'd78,8'd52} : s = 40;
	{8'd78,8'd53} : s = 168;
	{8'd78,8'd54} : s = 36;
	{8'd78,8'd55} : s = 164;
	{8'd78,8'd56} : s = 162;
	{8'd78,8'd57} : s = 323;
	{8'd78,8'd58} : s = 34;
	{8'd78,8'd59} : s = 161;
	{8'd78,8'd60} : s = 152;
	{8'd78,8'd61} : s = 312;
	{8'd78,8'd62} : s = 148;
	{8'd78,8'd63} : s = 308;
	{8'd78,8'd64} : s = 306;
	{8'd78,8'd65} : s = 425;
	{8'd78,8'd66} : s = 33;
	{8'd78,8'd67} : s = 146;
	{8'd78,8'd68} : s = 145;
	{8'd78,8'd69} : s = 305;
	{8'd78,8'd70} : s = 140;
	{8'd78,8'd71} : s = 300;
	{8'd78,8'd72} : s = 298;
	{8'd78,8'd73} : s = 422;
	{8'd78,8'd74} : s = 138;
	{8'd78,8'd75} : s = 297;
	{8'd78,8'd76} : s = 294;
	{8'd78,8'd77} : s = 421;
	{8'd78,8'd78} : s = 293;
	{8'd78,8'd79} : s = 419;
	{8'd78,8'd80} : s = 412;
	{8'd78,8'd81} : s = 486;
	{8'd78,8'd82} : s = 24;
	{8'd78,8'd83} : s = 137;
	{8'd78,8'd84} : s = 134;
	{8'd78,8'd85} : s = 291;
	{8'd78,8'd86} : s = 133;
	{8'd78,8'd87} : s = 284;
	{8'd78,8'd88} : s = 282;
	{8'd78,8'd89} : s = 410;
	{8'd78,8'd90} : s = 131;
	{8'd78,8'd91} : s = 281;
	{8'd78,8'd92} : s = 278;
	{8'd78,8'd93} : s = 409;
	{8'd78,8'd94} : s = 277;
	{8'd78,8'd95} : s = 406;
	{8'd78,8'd96} : s = 405;
	{8'd78,8'd97} : s = 485;
	{8'd78,8'd98} : s = 112;
	{8'd78,8'd99} : s = 275;
	{8'd78,8'd100} : s = 270;
	{8'd78,8'd101} : s = 403;
	{8'd78,8'd102} : s = 269;
	{8'd78,8'd103} : s = 398;
	{8'd78,8'd104} : s = 397;
	{8'd78,8'd105} : s = 483;
	{8'd78,8'd106} : s = 267;
	{8'd78,8'd107} : s = 395;
	{8'd78,8'd108} : s = 391;
	{8'd78,8'd109} : s = 476;
	{8'd78,8'd110} : s = 376;
	{8'd78,8'd111} : s = 474;
	{8'd78,8'd112} : s = 473;
	{8'd78,8'd113} : s = 506;
	{8'd78,8'd114} : s = 20;
	{8'd78,8'd115} : s = 104;
	{8'd78,8'd116} : s = 100;
	{8'd78,8'd117} : s = 263;
	{8'd78,8'd118} : s = 98;
	{8'd78,8'd119} : s = 240;
	{8'd78,8'd120} : s = 232;
	{8'd78,8'd121} : s = 372;
	{8'd78,8'd122} : s = 97;
	{8'd78,8'd123} : s = 228;
	{8'd78,8'd124} : s = 226;
	{8'd78,8'd125} : s = 370;
	{8'd78,8'd126} : s = 225;
	{8'd78,8'd127} : s = 369;
	{8'd78,8'd128} : s = 364;
	{8'd78,8'd129} : s = 470;
	{8'd78,8'd130} : s = 88;
	{8'd78,8'd131} : s = 216;
	{8'd78,8'd132} : s = 212;
	{8'd78,8'd133} : s = 362;
	{8'd78,8'd134} : s = 210;
	{8'd78,8'd135} : s = 361;
	{8'd78,8'd136} : s = 358;
	{8'd78,8'd137} : s = 469;
	{8'd78,8'd138} : s = 209;
	{8'd78,8'd139} : s = 357;
	{8'd78,8'd140} : s = 355;
	{8'd78,8'd141} : s = 467;
	{8'd78,8'd142} : s = 348;
	{8'd78,8'd143} : s = 462;
	{8'd78,8'd144} : s = 461;
	{8'd78,8'd145} : s = 505;
	{8'd78,8'd146} : s = 84;
	{8'd78,8'd147} : s = 204;
	{8'd78,8'd148} : s = 202;
	{8'd78,8'd149} : s = 346;
	{8'd78,8'd150} : s = 201;
	{8'd78,8'd151} : s = 345;
	{8'd78,8'd152} : s = 342;
	{8'd78,8'd153} : s = 459;
	{8'd78,8'd154} : s = 198;
	{8'd78,8'd155} : s = 341;
	{8'd78,8'd156} : s = 339;
	{8'd78,8'd157} : s = 455;
	{8'd78,8'd158} : s = 334;
	{8'd78,8'd159} : s = 444;
	{8'd78,8'd160} : s = 442;
	{8'd78,8'd161} : s = 502;
	{8'd78,8'd162} : s = 197;
	{8'd78,8'd163} : s = 333;
	{8'd78,8'd164} : s = 331;
	{8'd78,8'd165} : s = 441;
	{8'd78,8'd166} : s = 327;
	{8'd78,8'd167} : s = 438;
	{8'd78,8'd168} : s = 437;
	{8'd78,8'd169} : s = 501;
	{8'd78,8'd170} : s = 316;
	{8'd78,8'd171} : s = 435;
	{8'd78,8'd172} : s = 430;
	{8'd78,8'd173} : s = 499;
	{8'd78,8'd174} : s = 429;
	{8'd78,8'd175} : s = 494;
	{8'd78,8'd176} : s = 493;
	{8'd78,8'd177} : s = 510;
	{8'd78,8'd178} : s = 1;
	{8'd78,8'd179} : s = 18;
	{8'd78,8'd180} : s = 17;
	{8'd78,8'd181} : s = 82;
	{8'd78,8'd182} : s = 12;
	{8'd78,8'd183} : s = 81;
	{8'd78,8'd184} : s = 76;
	{8'd78,8'd185} : s = 195;
	{8'd78,8'd186} : s = 10;
	{8'd78,8'd187} : s = 74;
	{8'd78,8'd188} : s = 73;
	{8'd78,8'd189} : s = 184;
	{8'd78,8'd190} : s = 70;
	{8'd78,8'd191} : s = 180;
	{8'd78,8'd192} : s = 178;
	{8'd78,8'd193} : s = 314;
	{8'd78,8'd194} : s = 9;
	{8'd78,8'd195} : s = 69;
	{8'd78,8'd196} : s = 67;
	{8'd78,8'd197} : s = 177;
	{8'd78,8'd198} : s = 56;
	{8'd78,8'd199} : s = 172;
	{8'd78,8'd200} : s = 170;
	{8'd78,8'd201} : s = 313;
	{8'd78,8'd202} : s = 52;
	{8'd78,8'd203} : s = 169;
	{8'd78,8'd204} : s = 166;
	{8'd78,8'd205} : s = 310;
	{8'd78,8'd206} : s = 165;
	{8'd78,8'd207} : s = 309;
	{8'd78,8'd208} : s = 307;
	{8'd78,8'd209} : s = 427;
	{8'd78,8'd210} : s = 6;
	{8'd78,8'd211} : s = 50;
	{8'd78,8'd212} : s = 49;
	{8'd78,8'd213} : s = 163;
	{8'd78,8'd214} : s = 44;
	{8'd78,8'd215} : s = 156;
	{8'd78,8'd216} : s = 154;
	{8'd78,8'd217} : s = 302;
	{8'd78,8'd218} : s = 42;
	{8'd78,8'd219} : s = 153;
	{8'd78,8'd220} : s = 150;
	{8'd78,8'd221} : s = 301;
	{8'd78,8'd222} : s = 149;
	{8'd78,8'd223} : s = 299;
	{8'd78,8'd224} : s = 295;
	{8'd78,8'd225} : s = 423;
	{8'd78,8'd226} : s = 41;
	{8'd78,8'd227} : s = 147;
	{8'd78,8'd228} : s = 142;
	{8'd78,8'd229} : s = 286;
	{8'd78,8'd230} : s = 141;
	{8'd78,8'd231} : s = 285;
	{8'd78,8'd232} : s = 283;
	{8'd78,8'd233} : s = 414;
	{8'd78,8'd234} : s = 139;
	{8'd78,8'd235} : s = 279;
	{8'd78,8'd236} : s = 271;
	{8'd78,8'd237} : s = 413;
	{8'd78,8'd238} : s = 248;
	{8'd78,8'd239} : s = 411;
	{8'd78,8'd240} : s = 407;
	{8'd78,8'd241} : s = 491;
	{8'd78,8'd242} : s = 5;
	{8'd78,8'd243} : s = 38;
	{8'd78,8'd244} : s = 37;
	{8'd78,8'd245} : s = 135;
	{8'd78,8'd246} : s = 35;
	{8'd78,8'd247} : s = 120;
	{8'd78,8'd248} : s = 116;
	{8'd78,8'd249} : s = 244;
	{8'd78,8'd250} : s = 28;
	{8'd78,8'd251} : s = 114;
	{8'd78,8'd252} : s = 113;
	{8'd78,8'd253} : s = 242;
	{8'd78,8'd254} : s = 108;
	{8'd78,8'd255} : s = 241;
	{8'd79,8'd0} : s = 468;
	{8'd79,8'd1} : s = 66;
	{8'd79,8'd2} : s = 261;
	{8'd79,8'd3} : s = 259;
	{8'd79,8'd4} : s = 389;
	{8'd79,8'd5} : s = 224;
	{8'd79,8'd6} : s = 387;
	{8'd79,8'd7} : s = 368;
	{8'd79,8'd8} : s = 466;
	{8'd79,8'd9} : s = 208;
	{8'd79,8'd10} : s = 360;
	{8'd79,8'd11} : s = 356;
	{8'd79,8'd12} : s = 465;
	{8'd79,8'd13} : s = 354;
	{8'd79,8'd14} : s = 460;
	{8'd79,8'd15} : s = 458;
	{8'd79,8'd16} : s = 500;
	{8'd79,8'd17} : s = 65;
	{8'd79,8'd18} : s = 200;
	{8'd79,8'd19} : s = 196;
	{8'd79,8'd20} : s = 353;
	{8'd79,8'd21} : s = 194;
	{8'd79,8'd22} : s = 344;
	{8'd79,8'd23} : s = 340;
	{8'd79,8'd24} : s = 457;
	{8'd79,8'd25} : s = 193;
	{8'd79,8'd26} : s = 338;
	{8'd79,8'd27} : s = 337;
	{8'd79,8'd28} : s = 454;
	{8'd79,8'd29} : s = 332;
	{8'd79,8'd30} : s = 453;
	{8'd79,8'd31} : s = 451;
	{8'd79,8'd32} : s = 498;
	{8'd79,8'd33} : s = 176;
	{8'd79,8'd34} : s = 330;
	{8'd79,8'd35} : s = 329;
	{8'd79,8'd36} : s = 440;
	{8'd79,8'd37} : s = 326;
	{8'd79,8'd38} : s = 436;
	{8'd79,8'd39} : s = 434;
	{8'd79,8'd40} : s = 497;
	{8'd79,8'd41} : s = 325;
	{8'd79,8'd42} : s = 433;
	{8'd79,8'd43} : s = 428;
	{8'd79,8'd44} : s = 492;
	{8'd79,8'd45} : s = 426;
	{8'd79,8'd46} : s = 490;
	{8'd79,8'd47} : s = 489;
	{8'd79,8'd48} : s = 508;
	{8'd79,8'd49} : s = 2;
	{8'd79,8'd50} : s = 48;
	{8'd79,8'd51} : s = 40;
	{8'd79,8'd52} : s = 168;
	{8'd79,8'd53} : s = 36;
	{8'd79,8'd54} : s = 164;
	{8'd79,8'd55} : s = 162;
	{8'd79,8'd56} : s = 323;
	{8'd79,8'd57} : s = 34;
	{8'd79,8'd58} : s = 161;
	{8'd79,8'd59} : s = 152;
	{8'd79,8'd60} : s = 312;
	{8'd79,8'd61} : s = 148;
	{8'd79,8'd62} : s = 308;
	{8'd79,8'd63} : s = 306;
	{8'd79,8'd64} : s = 425;
	{8'd79,8'd65} : s = 33;
	{8'd79,8'd66} : s = 146;
	{8'd79,8'd67} : s = 145;
	{8'd79,8'd68} : s = 305;
	{8'd79,8'd69} : s = 140;
	{8'd79,8'd70} : s = 300;
	{8'd79,8'd71} : s = 298;
	{8'd79,8'd72} : s = 422;
	{8'd79,8'd73} : s = 138;
	{8'd79,8'd74} : s = 297;
	{8'd79,8'd75} : s = 294;
	{8'd79,8'd76} : s = 421;
	{8'd79,8'd77} : s = 293;
	{8'd79,8'd78} : s = 419;
	{8'd79,8'd79} : s = 412;
	{8'd79,8'd80} : s = 486;
	{8'd79,8'd81} : s = 24;
	{8'd79,8'd82} : s = 137;
	{8'd79,8'd83} : s = 134;
	{8'd79,8'd84} : s = 291;
	{8'd79,8'd85} : s = 133;
	{8'd79,8'd86} : s = 284;
	{8'd79,8'd87} : s = 282;
	{8'd79,8'd88} : s = 410;
	{8'd79,8'd89} : s = 131;
	{8'd79,8'd90} : s = 281;
	{8'd79,8'd91} : s = 278;
	{8'd79,8'd92} : s = 409;
	{8'd79,8'd93} : s = 277;
	{8'd79,8'd94} : s = 406;
	{8'd79,8'd95} : s = 405;
	{8'd79,8'd96} : s = 485;
	{8'd79,8'd97} : s = 112;
	{8'd79,8'd98} : s = 275;
	{8'd79,8'd99} : s = 270;
	{8'd79,8'd100} : s = 403;
	{8'd79,8'd101} : s = 269;
	{8'd79,8'd102} : s = 398;
	{8'd79,8'd103} : s = 397;
	{8'd79,8'd104} : s = 483;
	{8'd79,8'd105} : s = 267;
	{8'd79,8'd106} : s = 395;
	{8'd79,8'd107} : s = 391;
	{8'd79,8'd108} : s = 476;
	{8'd79,8'd109} : s = 376;
	{8'd79,8'd110} : s = 474;
	{8'd79,8'd111} : s = 473;
	{8'd79,8'd112} : s = 506;
	{8'd79,8'd113} : s = 20;
	{8'd79,8'd114} : s = 104;
	{8'd79,8'd115} : s = 100;
	{8'd79,8'd116} : s = 263;
	{8'd79,8'd117} : s = 98;
	{8'd79,8'd118} : s = 240;
	{8'd79,8'd119} : s = 232;
	{8'd79,8'd120} : s = 372;
	{8'd79,8'd121} : s = 97;
	{8'd79,8'd122} : s = 228;
	{8'd79,8'd123} : s = 226;
	{8'd79,8'd124} : s = 370;
	{8'd79,8'd125} : s = 225;
	{8'd79,8'd126} : s = 369;
	{8'd79,8'd127} : s = 364;
	{8'd79,8'd128} : s = 470;
	{8'd79,8'd129} : s = 88;
	{8'd79,8'd130} : s = 216;
	{8'd79,8'd131} : s = 212;
	{8'd79,8'd132} : s = 362;
	{8'd79,8'd133} : s = 210;
	{8'd79,8'd134} : s = 361;
	{8'd79,8'd135} : s = 358;
	{8'd79,8'd136} : s = 469;
	{8'd79,8'd137} : s = 209;
	{8'd79,8'd138} : s = 357;
	{8'd79,8'd139} : s = 355;
	{8'd79,8'd140} : s = 467;
	{8'd79,8'd141} : s = 348;
	{8'd79,8'd142} : s = 462;
	{8'd79,8'd143} : s = 461;
	{8'd79,8'd144} : s = 505;
	{8'd79,8'd145} : s = 84;
	{8'd79,8'd146} : s = 204;
	{8'd79,8'd147} : s = 202;
	{8'd79,8'd148} : s = 346;
	{8'd79,8'd149} : s = 201;
	{8'd79,8'd150} : s = 345;
	{8'd79,8'd151} : s = 342;
	{8'd79,8'd152} : s = 459;
	{8'd79,8'd153} : s = 198;
	{8'd79,8'd154} : s = 341;
	{8'd79,8'd155} : s = 339;
	{8'd79,8'd156} : s = 455;
	{8'd79,8'd157} : s = 334;
	{8'd79,8'd158} : s = 444;
	{8'd79,8'd159} : s = 442;
	{8'd79,8'd160} : s = 502;
	{8'd79,8'd161} : s = 197;
	{8'd79,8'd162} : s = 333;
	{8'd79,8'd163} : s = 331;
	{8'd79,8'd164} : s = 441;
	{8'd79,8'd165} : s = 327;
	{8'd79,8'd166} : s = 438;
	{8'd79,8'd167} : s = 437;
	{8'd79,8'd168} : s = 501;
	{8'd79,8'd169} : s = 316;
	{8'd79,8'd170} : s = 435;
	{8'd79,8'd171} : s = 430;
	{8'd79,8'd172} : s = 499;
	{8'd79,8'd173} : s = 429;
	{8'd79,8'd174} : s = 494;
	{8'd79,8'd175} : s = 493;
	{8'd79,8'd176} : s = 510;
	{8'd79,8'd177} : s = 1;
	{8'd79,8'd178} : s = 18;
	{8'd79,8'd179} : s = 17;
	{8'd79,8'd180} : s = 82;
	{8'd79,8'd181} : s = 12;
	{8'd79,8'd182} : s = 81;
	{8'd79,8'd183} : s = 76;
	{8'd79,8'd184} : s = 195;
	{8'd79,8'd185} : s = 10;
	{8'd79,8'd186} : s = 74;
	{8'd79,8'd187} : s = 73;
	{8'd79,8'd188} : s = 184;
	{8'd79,8'd189} : s = 70;
	{8'd79,8'd190} : s = 180;
	{8'd79,8'd191} : s = 178;
	{8'd79,8'd192} : s = 314;
	{8'd79,8'd193} : s = 9;
	{8'd79,8'd194} : s = 69;
	{8'd79,8'd195} : s = 67;
	{8'd79,8'd196} : s = 177;
	{8'd79,8'd197} : s = 56;
	{8'd79,8'd198} : s = 172;
	{8'd79,8'd199} : s = 170;
	{8'd79,8'd200} : s = 313;
	{8'd79,8'd201} : s = 52;
	{8'd79,8'd202} : s = 169;
	{8'd79,8'd203} : s = 166;
	{8'd79,8'd204} : s = 310;
	{8'd79,8'd205} : s = 165;
	{8'd79,8'd206} : s = 309;
	{8'd79,8'd207} : s = 307;
	{8'd79,8'd208} : s = 427;
	{8'd79,8'd209} : s = 6;
	{8'd79,8'd210} : s = 50;
	{8'd79,8'd211} : s = 49;
	{8'd79,8'd212} : s = 163;
	{8'd79,8'd213} : s = 44;
	{8'd79,8'd214} : s = 156;
	{8'd79,8'd215} : s = 154;
	{8'd79,8'd216} : s = 302;
	{8'd79,8'd217} : s = 42;
	{8'd79,8'd218} : s = 153;
	{8'd79,8'd219} : s = 150;
	{8'd79,8'd220} : s = 301;
	{8'd79,8'd221} : s = 149;
	{8'd79,8'd222} : s = 299;
	{8'd79,8'd223} : s = 295;
	{8'd79,8'd224} : s = 423;
	{8'd79,8'd225} : s = 41;
	{8'd79,8'd226} : s = 147;
	{8'd79,8'd227} : s = 142;
	{8'd79,8'd228} : s = 286;
	{8'd79,8'd229} : s = 141;
	{8'd79,8'd230} : s = 285;
	{8'd79,8'd231} : s = 283;
	{8'd79,8'd232} : s = 414;
	{8'd79,8'd233} : s = 139;
	{8'd79,8'd234} : s = 279;
	{8'd79,8'd235} : s = 271;
	{8'd79,8'd236} : s = 413;
	{8'd79,8'd237} : s = 248;
	{8'd79,8'd238} : s = 411;
	{8'd79,8'd239} : s = 407;
	{8'd79,8'd240} : s = 491;
	{8'd79,8'd241} : s = 5;
	{8'd79,8'd242} : s = 38;
	{8'd79,8'd243} : s = 37;
	{8'd79,8'd244} : s = 135;
	{8'd79,8'd245} : s = 35;
	{8'd79,8'd246} : s = 120;
	{8'd79,8'd247} : s = 116;
	{8'd79,8'd248} : s = 244;
	{8'd79,8'd249} : s = 28;
	{8'd79,8'd250} : s = 114;
	{8'd79,8'd251} : s = 113;
	{8'd79,8'd252} : s = 242;
	{8'd79,8'd253} : s = 108;
	{8'd79,8'd254} : s = 241;
	{8'd79,8'd255} : s = 236;
	{8'd80,8'd0} : s = 66;
	{8'd80,8'd1} : s = 261;
	{8'd80,8'd2} : s = 259;
	{8'd80,8'd3} : s = 389;
	{8'd80,8'd4} : s = 224;
	{8'd80,8'd5} : s = 387;
	{8'd80,8'd6} : s = 368;
	{8'd80,8'd7} : s = 466;
	{8'd80,8'd8} : s = 208;
	{8'd80,8'd9} : s = 360;
	{8'd80,8'd10} : s = 356;
	{8'd80,8'd11} : s = 465;
	{8'd80,8'd12} : s = 354;
	{8'd80,8'd13} : s = 460;
	{8'd80,8'd14} : s = 458;
	{8'd80,8'd15} : s = 500;
	{8'd80,8'd16} : s = 65;
	{8'd80,8'd17} : s = 200;
	{8'd80,8'd18} : s = 196;
	{8'd80,8'd19} : s = 353;
	{8'd80,8'd20} : s = 194;
	{8'd80,8'd21} : s = 344;
	{8'd80,8'd22} : s = 340;
	{8'd80,8'd23} : s = 457;
	{8'd80,8'd24} : s = 193;
	{8'd80,8'd25} : s = 338;
	{8'd80,8'd26} : s = 337;
	{8'd80,8'd27} : s = 454;
	{8'd80,8'd28} : s = 332;
	{8'd80,8'd29} : s = 453;
	{8'd80,8'd30} : s = 451;
	{8'd80,8'd31} : s = 498;
	{8'd80,8'd32} : s = 176;
	{8'd80,8'd33} : s = 330;
	{8'd80,8'd34} : s = 329;
	{8'd80,8'd35} : s = 440;
	{8'd80,8'd36} : s = 326;
	{8'd80,8'd37} : s = 436;
	{8'd80,8'd38} : s = 434;
	{8'd80,8'd39} : s = 497;
	{8'd80,8'd40} : s = 325;
	{8'd80,8'd41} : s = 433;
	{8'd80,8'd42} : s = 428;
	{8'd80,8'd43} : s = 492;
	{8'd80,8'd44} : s = 426;
	{8'd80,8'd45} : s = 490;
	{8'd80,8'd46} : s = 489;
	{8'd80,8'd47} : s = 508;
	{8'd80,8'd48} : s = 2;
	{8'd80,8'd49} : s = 48;
	{8'd80,8'd50} : s = 40;
	{8'd80,8'd51} : s = 168;
	{8'd80,8'd52} : s = 36;
	{8'd80,8'd53} : s = 164;
	{8'd80,8'd54} : s = 162;
	{8'd80,8'd55} : s = 323;
	{8'd80,8'd56} : s = 34;
	{8'd80,8'd57} : s = 161;
	{8'd80,8'd58} : s = 152;
	{8'd80,8'd59} : s = 312;
	{8'd80,8'd60} : s = 148;
	{8'd80,8'd61} : s = 308;
	{8'd80,8'd62} : s = 306;
	{8'd80,8'd63} : s = 425;
	{8'd80,8'd64} : s = 33;
	{8'd80,8'd65} : s = 146;
	{8'd80,8'd66} : s = 145;
	{8'd80,8'd67} : s = 305;
	{8'd80,8'd68} : s = 140;
	{8'd80,8'd69} : s = 300;
	{8'd80,8'd70} : s = 298;
	{8'd80,8'd71} : s = 422;
	{8'd80,8'd72} : s = 138;
	{8'd80,8'd73} : s = 297;
	{8'd80,8'd74} : s = 294;
	{8'd80,8'd75} : s = 421;
	{8'd80,8'd76} : s = 293;
	{8'd80,8'd77} : s = 419;
	{8'd80,8'd78} : s = 412;
	{8'd80,8'd79} : s = 486;
	{8'd80,8'd80} : s = 24;
	{8'd80,8'd81} : s = 137;
	{8'd80,8'd82} : s = 134;
	{8'd80,8'd83} : s = 291;
	{8'd80,8'd84} : s = 133;
	{8'd80,8'd85} : s = 284;
	{8'd80,8'd86} : s = 282;
	{8'd80,8'd87} : s = 410;
	{8'd80,8'd88} : s = 131;
	{8'd80,8'd89} : s = 281;
	{8'd80,8'd90} : s = 278;
	{8'd80,8'd91} : s = 409;
	{8'd80,8'd92} : s = 277;
	{8'd80,8'd93} : s = 406;
	{8'd80,8'd94} : s = 405;
	{8'd80,8'd95} : s = 485;
	{8'd80,8'd96} : s = 112;
	{8'd80,8'd97} : s = 275;
	{8'd80,8'd98} : s = 270;
	{8'd80,8'd99} : s = 403;
	{8'd80,8'd100} : s = 269;
	{8'd80,8'd101} : s = 398;
	{8'd80,8'd102} : s = 397;
	{8'd80,8'd103} : s = 483;
	{8'd80,8'd104} : s = 267;
	{8'd80,8'd105} : s = 395;
	{8'd80,8'd106} : s = 391;
	{8'd80,8'd107} : s = 476;
	{8'd80,8'd108} : s = 376;
	{8'd80,8'd109} : s = 474;
	{8'd80,8'd110} : s = 473;
	{8'd80,8'd111} : s = 506;
	{8'd80,8'd112} : s = 20;
	{8'd80,8'd113} : s = 104;
	{8'd80,8'd114} : s = 100;
	{8'd80,8'd115} : s = 263;
	{8'd80,8'd116} : s = 98;
	{8'd80,8'd117} : s = 240;
	{8'd80,8'd118} : s = 232;
	{8'd80,8'd119} : s = 372;
	{8'd80,8'd120} : s = 97;
	{8'd80,8'd121} : s = 228;
	{8'd80,8'd122} : s = 226;
	{8'd80,8'd123} : s = 370;
	{8'd80,8'd124} : s = 225;
	{8'd80,8'd125} : s = 369;
	{8'd80,8'd126} : s = 364;
	{8'd80,8'd127} : s = 470;
	{8'd80,8'd128} : s = 88;
	{8'd80,8'd129} : s = 216;
	{8'd80,8'd130} : s = 212;
	{8'd80,8'd131} : s = 362;
	{8'd80,8'd132} : s = 210;
	{8'd80,8'd133} : s = 361;
	{8'd80,8'd134} : s = 358;
	{8'd80,8'd135} : s = 469;
	{8'd80,8'd136} : s = 209;
	{8'd80,8'd137} : s = 357;
	{8'd80,8'd138} : s = 355;
	{8'd80,8'd139} : s = 467;
	{8'd80,8'd140} : s = 348;
	{8'd80,8'd141} : s = 462;
	{8'd80,8'd142} : s = 461;
	{8'd80,8'd143} : s = 505;
	{8'd80,8'd144} : s = 84;
	{8'd80,8'd145} : s = 204;
	{8'd80,8'd146} : s = 202;
	{8'd80,8'd147} : s = 346;
	{8'd80,8'd148} : s = 201;
	{8'd80,8'd149} : s = 345;
	{8'd80,8'd150} : s = 342;
	{8'd80,8'd151} : s = 459;
	{8'd80,8'd152} : s = 198;
	{8'd80,8'd153} : s = 341;
	{8'd80,8'd154} : s = 339;
	{8'd80,8'd155} : s = 455;
	{8'd80,8'd156} : s = 334;
	{8'd80,8'd157} : s = 444;
	{8'd80,8'd158} : s = 442;
	{8'd80,8'd159} : s = 502;
	{8'd80,8'd160} : s = 197;
	{8'd80,8'd161} : s = 333;
	{8'd80,8'd162} : s = 331;
	{8'd80,8'd163} : s = 441;
	{8'd80,8'd164} : s = 327;
	{8'd80,8'd165} : s = 438;
	{8'd80,8'd166} : s = 437;
	{8'd80,8'd167} : s = 501;
	{8'd80,8'd168} : s = 316;
	{8'd80,8'd169} : s = 435;
	{8'd80,8'd170} : s = 430;
	{8'd80,8'd171} : s = 499;
	{8'd80,8'd172} : s = 429;
	{8'd80,8'd173} : s = 494;
	{8'd80,8'd174} : s = 493;
	{8'd80,8'd175} : s = 510;
	{8'd80,8'd176} : s = 1;
	{8'd80,8'd177} : s = 18;
	{8'd80,8'd178} : s = 17;
	{8'd80,8'd179} : s = 82;
	{8'd80,8'd180} : s = 12;
	{8'd80,8'd181} : s = 81;
	{8'd80,8'd182} : s = 76;
	{8'd80,8'd183} : s = 195;
	{8'd80,8'd184} : s = 10;
	{8'd80,8'd185} : s = 74;
	{8'd80,8'd186} : s = 73;
	{8'd80,8'd187} : s = 184;
	{8'd80,8'd188} : s = 70;
	{8'd80,8'd189} : s = 180;
	{8'd80,8'd190} : s = 178;
	{8'd80,8'd191} : s = 314;
	{8'd80,8'd192} : s = 9;
	{8'd80,8'd193} : s = 69;
	{8'd80,8'd194} : s = 67;
	{8'd80,8'd195} : s = 177;
	{8'd80,8'd196} : s = 56;
	{8'd80,8'd197} : s = 172;
	{8'd80,8'd198} : s = 170;
	{8'd80,8'd199} : s = 313;
	{8'd80,8'd200} : s = 52;
	{8'd80,8'd201} : s = 169;
	{8'd80,8'd202} : s = 166;
	{8'd80,8'd203} : s = 310;
	{8'd80,8'd204} : s = 165;
	{8'd80,8'd205} : s = 309;
	{8'd80,8'd206} : s = 307;
	{8'd80,8'd207} : s = 427;
	{8'd80,8'd208} : s = 6;
	{8'd80,8'd209} : s = 50;
	{8'd80,8'd210} : s = 49;
	{8'd80,8'd211} : s = 163;
	{8'd80,8'd212} : s = 44;
	{8'd80,8'd213} : s = 156;
	{8'd80,8'd214} : s = 154;
	{8'd80,8'd215} : s = 302;
	{8'd80,8'd216} : s = 42;
	{8'd80,8'd217} : s = 153;
	{8'd80,8'd218} : s = 150;
	{8'd80,8'd219} : s = 301;
	{8'd80,8'd220} : s = 149;
	{8'd80,8'd221} : s = 299;
	{8'd80,8'd222} : s = 295;
	{8'd80,8'd223} : s = 423;
	{8'd80,8'd224} : s = 41;
	{8'd80,8'd225} : s = 147;
	{8'd80,8'd226} : s = 142;
	{8'd80,8'd227} : s = 286;
	{8'd80,8'd228} : s = 141;
	{8'd80,8'd229} : s = 285;
	{8'd80,8'd230} : s = 283;
	{8'd80,8'd231} : s = 414;
	{8'd80,8'd232} : s = 139;
	{8'd80,8'd233} : s = 279;
	{8'd80,8'd234} : s = 271;
	{8'd80,8'd235} : s = 413;
	{8'd80,8'd236} : s = 248;
	{8'd80,8'd237} : s = 411;
	{8'd80,8'd238} : s = 407;
	{8'd80,8'd239} : s = 491;
	{8'd80,8'd240} : s = 5;
	{8'd80,8'd241} : s = 38;
	{8'd80,8'd242} : s = 37;
	{8'd80,8'd243} : s = 135;
	{8'd80,8'd244} : s = 35;
	{8'd80,8'd245} : s = 120;
	{8'd80,8'd246} : s = 116;
	{8'd80,8'd247} : s = 244;
	{8'd80,8'd248} : s = 28;
	{8'd80,8'd249} : s = 114;
	{8'd80,8'd250} : s = 113;
	{8'd80,8'd251} : s = 242;
	{8'd80,8'd252} : s = 108;
	{8'd80,8'd253} : s = 241;
	{8'd80,8'd254} : s = 236;
	{8'd80,8'd255} : s = 399;
	{8'd81,8'd0} : s = 261;
	{8'd81,8'd1} : s = 259;
	{8'd81,8'd2} : s = 389;
	{8'd81,8'd3} : s = 224;
	{8'd81,8'd4} : s = 387;
	{8'd81,8'd5} : s = 368;
	{8'd81,8'd6} : s = 466;
	{8'd81,8'd7} : s = 208;
	{8'd81,8'd8} : s = 360;
	{8'd81,8'd9} : s = 356;
	{8'd81,8'd10} : s = 465;
	{8'd81,8'd11} : s = 354;
	{8'd81,8'd12} : s = 460;
	{8'd81,8'd13} : s = 458;
	{8'd81,8'd14} : s = 500;
	{8'd81,8'd15} : s = 65;
	{8'd81,8'd16} : s = 200;
	{8'd81,8'd17} : s = 196;
	{8'd81,8'd18} : s = 353;
	{8'd81,8'd19} : s = 194;
	{8'd81,8'd20} : s = 344;
	{8'd81,8'd21} : s = 340;
	{8'd81,8'd22} : s = 457;
	{8'd81,8'd23} : s = 193;
	{8'd81,8'd24} : s = 338;
	{8'd81,8'd25} : s = 337;
	{8'd81,8'd26} : s = 454;
	{8'd81,8'd27} : s = 332;
	{8'd81,8'd28} : s = 453;
	{8'd81,8'd29} : s = 451;
	{8'd81,8'd30} : s = 498;
	{8'd81,8'd31} : s = 176;
	{8'd81,8'd32} : s = 330;
	{8'd81,8'd33} : s = 329;
	{8'd81,8'd34} : s = 440;
	{8'd81,8'd35} : s = 326;
	{8'd81,8'd36} : s = 436;
	{8'd81,8'd37} : s = 434;
	{8'd81,8'd38} : s = 497;
	{8'd81,8'd39} : s = 325;
	{8'd81,8'd40} : s = 433;
	{8'd81,8'd41} : s = 428;
	{8'd81,8'd42} : s = 492;
	{8'd81,8'd43} : s = 426;
	{8'd81,8'd44} : s = 490;
	{8'd81,8'd45} : s = 489;
	{8'd81,8'd46} : s = 508;
	{8'd81,8'd47} : s = 2;
	{8'd81,8'd48} : s = 48;
	{8'd81,8'd49} : s = 40;
	{8'd81,8'd50} : s = 168;
	{8'd81,8'd51} : s = 36;
	{8'd81,8'd52} : s = 164;
	{8'd81,8'd53} : s = 162;
	{8'd81,8'd54} : s = 323;
	{8'd81,8'd55} : s = 34;
	{8'd81,8'd56} : s = 161;
	{8'd81,8'd57} : s = 152;
	{8'd81,8'd58} : s = 312;
	{8'd81,8'd59} : s = 148;
	{8'd81,8'd60} : s = 308;
	{8'd81,8'd61} : s = 306;
	{8'd81,8'd62} : s = 425;
	{8'd81,8'd63} : s = 33;
	{8'd81,8'd64} : s = 146;
	{8'd81,8'd65} : s = 145;
	{8'd81,8'd66} : s = 305;
	{8'd81,8'd67} : s = 140;
	{8'd81,8'd68} : s = 300;
	{8'd81,8'd69} : s = 298;
	{8'd81,8'd70} : s = 422;
	{8'd81,8'd71} : s = 138;
	{8'd81,8'd72} : s = 297;
	{8'd81,8'd73} : s = 294;
	{8'd81,8'd74} : s = 421;
	{8'd81,8'd75} : s = 293;
	{8'd81,8'd76} : s = 419;
	{8'd81,8'd77} : s = 412;
	{8'd81,8'd78} : s = 486;
	{8'd81,8'd79} : s = 24;
	{8'd81,8'd80} : s = 137;
	{8'd81,8'd81} : s = 134;
	{8'd81,8'd82} : s = 291;
	{8'd81,8'd83} : s = 133;
	{8'd81,8'd84} : s = 284;
	{8'd81,8'd85} : s = 282;
	{8'd81,8'd86} : s = 410;
	{8'd81,8'd87} : s = 131;
	{8'd81,8'd88} : s = 281;
	{8'd81,8'd89} : s = 278;
	{8'd81,8'd90} : s = 409;
	{8'd81,8'd91} : s = 277;
	{8'd81,8'd92} : s = 406;
	{8'd81,8'd93} : s = 405;
	{8'd81,8'd94} : s = 485;
	{8'd81,8'd95} : s = 112;
	{8'd81,8'd96} : s = 275;
	{8'd81,8'd97} : s = 270;
	{8'd81,8'd98} : s = 403;
	{8'd81,8'd99} : s = 269;
	{8'd81,8'd100} : s = 398;
	{8'd81,8'd101} : s = 397;
	{8'd81,8'd102} : s = 483;
	{8'd81,8'd103} : s = 267;
	{8'd81,8'd104} : s = 395;
	{8'd81,8'd105} : s = 391;
	{8'd81,8'd106} : s = 476;
	{8'd81,8'd107} : s = 376;
	{8'd81,8'd108} : s = 474;
	{8'd81,8'd109} : s = 473;
	{8'd81,8'd110} : s = 506;
	{8'd81,8'd111} : s = 20;
	{8'd81,8'd112} : s = 104;
	{8'd81,8'd113} : s = 100;
	{8'd81,8'd114} : s = 263;
	{8'd81,8'd115} : s = 98;
	{8'd81,8'd116} : s = 240;
	{8'd81,8'd117} : s = 232;
	{8'd81,8'd118} : s = 372;
	{8'd81,8'd119} : s = 97;
	{8'd81,8'd120} : s = 228;
	{8'd81,8'd121} : s = 226;
	{8'd81,8'd122} : s = 370;
	{8'd81,8'd123} : s = 225;
	{8'd81,8'd124} : s = 369;
	{8'd81,8'd125} : s = 364;
	{8'd81,8'd126} : s = 470;
	{8'd81,8'd127} : s = 88;
	{8'd81,8'd128} : s = 216;
	{8'd81,8'd129} : s = 212;
	{8'd81,8'd130} : s = 362;
	{8'd81,8'd131} : s = 210;
	{8'd81,8'd132} : s = 361;
	{8'd81,8'd133} : s = 358;
	{8'd81,8'd134} : s = 469;
	{8'd81,8'd135} : s = 209;
	{8'd81,8'd136} : s = 357;
	{8'd81,8'd137} : s = 355;
	{8'd81,8'd138} : s = 467;
	{8'd81,8'd139} : s = 348;
	{8'd81,8'd140} : s = 462;
	{8'd81,8'd141} : s = 461;
	{8'd81,8'd142} : s = 505;
	{8'd81,8'd143} : s = 84;
	{8'd81,8'd144} : s = 204;
	{8'd81,8'd145} : s = 202;
	{8'd81,8'd146} : s = 346;
	{8'd81,8'd147} : s = 201;
	{8'd81,8'd148} : s = 345;
	{8'd81,8'd149} : s = 342;
	{8'd81,8'd150} : s = 459;
	{8'd81,8'd151} : s = 198;
	{8'd81,8'd152} : s = 341;
	{8'd81,8'd153} : s = 339;
	{8'd81,8'd154} : s = 455;
	{8'd81,8'd155} : s = 334;
	{8'd81,8'd156} : s = 444;
	{8'd81,8'd157} : s = 442;
	{8'd81,8'd158} : s = 502;
	{8'd81,8'd159} : s = 197;
	{8'd81,8'd160} : s = 333;
	{8'd81,8'd161} : s = 331;
	{8'd81,8'd162} : s = 441;
	{8'd81,8'd163} : s = 327;
	{8'd81,8'd164} : s = 438;
	{8'd81,8'd165} : s = 437;
	{8'd81,8'd166} : s = 501;
	{8'd81,8'd167} : s = 316;
	{8'd81,8'd168} : s = 435;
	{8'd81,8'd169} : s = 430;
	{8'd81,8'd170} : s = 499;
	{8'd81,8'd171} : s = 429;
	{8'd81,8'd172} : s = 494;
	{8'd81,8'd173} : s = 493;
	{8'd81,8'd174} : s = 510;
	{8'd81,8'd175} : s = 1;
	{8'd81,8'd176} : s = 18;
	{8'd81,8'd177} : s = 17;
	{8'd81,8'd178} : s = 82;
	{8'd81,8'd179} : s = 12;
	{8'd81,8'd180} : s = 81;
	{8'd81,8'd181} : s = 76;
	{8'd81,8'd182} : s = 195;
	{8'd81,8'd183} : s = 10;
	{8'd81,8'd184} : s = 74;
	{8'd81,8'd185} : s = 73;
	{8'd81,8'd186} : s = 184;
	{8'd81,8'd187} : s = 70;
	{8'd81,8'd188} : s = 180;
	{8'd81,8'd189} : s = 178;
	{8'd81,8'd190} : s = 314;
	{8'd81,8'd191} : s = 9;
	{8'd81,8'd192} : s = 69;
	{8'd81,8'd193} : s = 67;
	{8'd81,8'd194} : s = 177;
	{8'd81,8'd195} : s = 56;
	{8'd81,8'd196} : s = 172;
	{8'd81,8'd197} : s = 170;
	{8'd81,8'd198} : s = 313;
	{8'd81,8'd199} : s = 52;
	{8'd81,8'd200} : s = 169;
	{8'd81,8'd201} : s = 166;
	{8'd81,8'd202} : s = 310;
	{8'd81,8'd203} : s = 165;
	{8'd81,8'd204} : s = 309;
	{8'd81,8'd205} : s = 307;
	{8'd81,8'd206} : s = 427;
	{8'd81,8'd207} : s = 6;
	{8'd81,8'd208} : s = 50;
	{8'd81,8'd209} : s = 49;
	{8'd81,8'd210} : s = 163;
	{8'd81,8'd211} : s = 44;
	{8'd81,8'd212} : s = 156;
	{8'd81,8'd213} : s = 154;
	{8'd81,8'd214} : s = 302;
	{8'd81,8'd215} : s = 42;
	{8'd81,8'd216} : s = 153;
	{8'd81,8'd217} : s = 150;
	{8'd81,8'd218} : s = 301;
	{8'd81,8'd219} : s = 149;
	{8'd81,8'd220} : s = 299;
	{8'd81,8'd221} : s = 295;
	{8'd81,8'd222} : s = 423;
	{8'd81,8'd223} : s = 41;
	{8'd81,8'd224} : s = 147;
	{8'd81,8'd225} : s = 142;
	{8'd81,8'd226} : s = 286;
	{8'd81,8'd227} : s = 141;
	{8'd81,8'd228} : s = 285;
	{8'd81,8'd229} : s = 283;
	{8'd81,8'd230} : s = 414;
	{8'd81,8'd231} : s = 139;
	{8'd81,8'd232} : s = 279;
	{8'd81,8'd233} : s = 271;
	{8'd81,8'd234} : s = 413;
	{8'd81,8'd235} : s = 248;
	{8'd81,8'd236} : s = 411;
	{8'd81,8'd237} : s = 407;
	{8'd81,8'd238} : s = 491;
	{8'd81,8'd239} : s = 5;
	{8'd81,8'd240} : s = 38;
	{8'd81,8'd241} : s = 37;
	{8'd81,8'd242} : s = 135;
	{8'd81,8'd243} : s = 35;
	{8'd81,8'd244} : s = 120;
	{8'd81,8'd245} : s = 116;
	{8'd81,8'd246} : s = 244;
	{8'd81,8'd247} : s = 28;
	{8'd81,8'd248} : s = 114;
	{8'd81,8'd249} : s = 113;
	{8'd81,8'd250} : s = 242;
	{8'd81,8'd251} : s = 108;
	{8'd81,8'd252} : s = 241;
	{8'd81,8'd253} : s = 236;
	{8'd81,8'd254} : s = 399;
	{8'd81,8'd255} : s = 26;
	{8'd82,8'd0} : s = 259;
	{8'd82,8'd1} : s = 389;
	{8'd82,8'd2} : s = 224;
	{8'd82,8'd3} : s = 387;
	{8'd82,8'd4} : s = 368;
	{8'd82,8'd5} : s = 466;
	{8'd82,8'd6} : s = 208;
	{8'd82,8'd7} : s = 360;
	{8'd82,8'd8} : s = 356;
	{8'd82,8'd9} : s = 465;
	{8'd82,8'd10} : s = 354;
	{8'd82,8'd11} : s = 460;
	{8'd82,8'd12} : s = 458;
	{8'd82,8'd13} : s = 500;
	{8'd82,8'd14} : s = 65;
	{8'd82,8'd15} : s = 200;
	{8'd82,8'd16} : s = 196;
	{8'd82,8'd17} : s = 353;
	{8'd82,8'd18} : s = 194;
	{8'd82,8'd19} : s = 344;
	{8'd82,8'd20} : s = 340;
	{8'd82,8'd21} : s = 457;
	{8'd82,8'd22} : s = 193;
	{8'd82,8'd23} : s = 338;
	{8'd82,8'd24} : s = 337;
	{8'd82,8'd25} : s = 454;
	{8'd82,8'd26} : s = 332;
	{8'd82,8'd27} : s = 453;
	{8'd82,8'd28} : s = 451;
	{8'd82,8'd29} : s = 498;
	{8'd82,8'd30} : s = 176;
	{8'd82,8'd31} : s = 330;
	{8'd82,8'd32} : s = 329;
	{8'd82,8'd33} : s = 440;
	{8'd82,8'd34} : s = 326;
	{8'd82,8'd35} : s = 436;
	{8'd82,8'd36} : s = 434;
	{8'd82,8'd37} : s = 497;
	{8'd82,8'd38} : s = 325;
	{8'd82,8'd39} : s = 433;
	{8'd82,8'd40} : s = 428;
	{8'd82,8'd41} : s = 492;
	{8'd82,8'd42} : s = 426;
	{8'd82,8'd43} : s = 490;
	{8'd82,8'd44} : s = 489;
	{8'd82,8'd45} : s = 508;
	{8'd82,8'd46} : s = 2;
	{8'd82,8'd47} : s = 48;
	{8'd82,8'd48} : s = 40;
	{8'd82,8'd49} : s = 168;
	{8'd82,8'd50} : s = 36;
	{8'd82,8'd51} : s = 164;
	{8'd82,8'd52} : s = 162;
	{8'd82,8'd53} : s = 323;
	{8'd82,8'd54} : s = 34;
	{8'd82,8'd55} : s = 161;
	{8'd82,8'd56} : s = 152;
	{8'd82,8'd57} : s = 312;
	{8'd82,8'd58} : s = 148;
	{8'd82,8'd59} : s = 308;
	{8'd82,8'd60} : s = 306;
	{8'd82,8'd61} : s = 425;
	{8'd82,8'd62} : s = 33;
	{8'd82,8'd63} : s = 146;
	{8'd82,8'd64} : s = 145;
	{8'd82,8'd65} : s = 305;
	{8'd82,8'd66} : s = 140;
	{8'd82,8'd67} : s = 300;
	{8'd82,8'd68} : s = 298;
	{8'd82,8'd69} : s = 422;
	{8'd82,8'd70} : s = 138;
	{8'd82,8'd71} : s = 297;
	{8'd82,8'd72} : s = 294;
	{8'd82,8'd73} : s = 421;
	{8'd82,8'd74} : s = 293;
	{8'd82,8'd75} : s = 419;
	{8'd82,8'd76} : s = 412;
	{8'd82,8'd77} : s = 486;
	{8'd82,8'd78} : s = 24;
	{8'd82,8'd79} : s = 137;
	{8'd82,8'd80} : s = 134;
	{8'd82,8'd81} : s = 291;
	{8'd82,8'd82} : s = 133;
	{8'd82,8'd83} : s = 284;
	{8'd82,8'd84} : s = 282;
	{8'd82,8'd85} : s = 410;
	{8'd82,8'd86} : s = 131;
	{8'd82,8'd87} : s = 281;
	{8'd82,8'd88} : s = 278;
	{8'd82,8'd89} : s = 409;
	{8'd82,8'd90} : s = 277;
	{8'd82,8'd91} : s = 406;
	{8'd82,8'd92} : s = 405;
	{8'd82,8'd93} : s = 485;
	{8'd82,8'd94} : s = 112;
	{8'd82,8'd95} : s = 275;
	{8'd82,8'd96} : s = 270;
	{8'd82,8'd97} : s = 403;
	{8'd82,8'd98} : s = 269;
	{8'd82,8'd99} : s = 398;
	{8'd82,8'd100} : s = 397;
	{8'd82,8'd101} : s = 483;
	{8'd82,8'd102} : s = 267;
	{8'd82,8'd103} : s = 395;
	{8'd82,8'd104} : s = 391;
	{8'd82,8'd105} : s = 476;
	{8'd82,8'd106} : s = 376;
	{8'd82,8'd107} : s = 474;
	{8'd82,8'd108} : s = 473;
	{8'd82,8'd109} : s = 506;
	{8'd82,8'd110} : s = 20;
	{8'd82,8'd111} : s = 104;
	{8'd82,8'd112} : s = 100;
	{8'd82,8'd113} : s = 263;
	{8'd82,8'd114} : s = 98;
	{8'd82,8'd115} : s = 240;
	{8'd82,8'd116} : s = 232;
	{8'd82,8'd117} : s = 372;
	{8'd82,8'd118} : s = 97;
	{8'd82,8'd119} : s = 228;
	{8'd82,8'd120} : s = 226;
	{8'd82,8'd121} : s = 370;
	{8'd82,8'd122} : s = 225;
	{8'd82,8'd123} : s = 369;
	{8'd82,8'd124} : s = 364;
	{8'd82,8'd125} : s = 470;
	{8'd82,8'd126} : s = 88;
	{8'd82,8'd127} : s = 216;
	{8'd82,8'd128} : s = 212;
	{8'd82,8'd129} : s = 362;
	{8'd82,8'd130} : s = 210;
	{8'd82,8'd131} : s = 361;
	{8'd82,8'd132} : s = 358;
	{8'd82,8'd133} : s = 469;
	{8'd82,8'd134} : s = 209;
	{8'd82,8'd135} : s = 357;
	{8'd82,8'd136} : s = 355;
	{8'd82,8'd137} : s = 467;
	{8'd82,8'd138} : s = 348;
	{8'd82,8'd139} : s = 462;
	{8'd82,8'd140} : s = 461;
	{8'd82,8'd141} : s = 505;
	{8'd82,8'd142} : s = 84;
	{8'd82,8'd143} : s = 204;
	{8'd82,8'd144} : s = 202;
	{8'd82,8'd145} : s = 346;
	{8'd82,8'd146} : s = 201;
	{8'd82,8'd147} : s = 345;
	{8'd82,8'd148} : s = 342;
	{8'd82,8'd149} : s = 459;
	{8'd82,8'd150} : s = 198;
	{8'd82,8'd151} : s = 341;
	{8'd82,8'd152} : s = 339;
	{8'd82,8'd153} : s = 455;
	{8'd82,8'd154} : s = 334;
	{8'd82,8'd155} : s = 444;
	{8'd82,8'd156} : s = 442;
	{8'd82,8'd157} : s = 502;
	{8'd82,8'd158} : s = 197;
	{8'd82,8'd159} : s = 333;
	{8'd82,8'd160} : s = 331;
	{8'd82,8'd161} : s = 441;
	{8'd82,8'd162} : s = 327;
	{8'd82,8'd163} : s = 438;
	{8'd82,8'd164} : s = 437;
	{8'd82,8'd165} : s = 501;
	{8'd82,8'd166} : s = 316;
	{8'd82,8'd167} : s = 435;
	{8'd82,8'd168} : s = 430;
	{8'd82,8'd169} : s = 499;
	{8'd82,8'd170} : s = 429;
	{8'd82,8'd171} : s = 494;
	{8'd82,8'd172} : s = 493;
	{8'd82,8'd173} : s = 510;
	{8'd82,8'd174} : s = 1;
	{8'd82,8'd175} : s = 18;
	{8'd82,8'd176} : s = 17;
	{8'd82,8'd177} : s = 82;
	{8'd82,8'd178} : s = 12;
	{8'd82,8'd179} : s = 81;
	{8'd82,8'd180} : s = 76;
	{8'd82,8'd181} : s = 195;
	{8'd82,8'd182} : s = 10;
	{8'd82,8'd183} : s = 74;
	{8'd82,8'd184} : s = 73;
	{8'd82,8'd185} : s = 184;
	{8'd82,8'd186} : s = 70;
	{8'd82,8'd187} : s = 180;
	{8'd82,8'd188} : s = 178;
	{8'd82,8'd189} : s = 314;
	{8'd82,8'd190} : s = 9;
	{8'd82,8'd191} : s = 69;
	{8'd82,8'd192} : s = 67;
	{8'd82,8'd193} : s = 177;
	{8'd82,8'd194} : s = 56;
	{8'd82,8'd195} : s = 172;
	{8'd82,8'd196} : s = 170;
	{8'd82,8'd197} : s = 313;
	{8'd82,8'd198} : s = 52;
	{8'd82,8'd199} : s = 169;
	{8'd82,8'd200} : s = 166;
	{8'd82,8'd201} : s = 310;
	{8'd82,8'd202} : s = 165;
	{8'd82,8'd203} : s = 309;
	{8'd82,8'd204} : s = 307;
	{8'd82,8'd205} : s = 427;
	{8'd82,8'd206} : s = 6;
	{8'd82,8'd207} : s = 50;
	{8'd82,8'd208} : s = 49;
	{8'd82,8'd209} : s = 163;
	{8'd82,8'd210} : s = 44;
	{8'd82,8'd211} : s = 156;
	{8'd82,8'd212} : s = 154;
	{8'd82,8'd213} : s = 302;
	{8'd82,8'd214} : s = 42;
	{8'd82,8'd215} : s = 153;
	{8'd82,8'd216} : s = 150;
	{8'd82,8'd217} : s = 301;
	{8'd82,8'd218} : s = 149;
	{8'd82,8'd219} : s = 299;
	{8'd82,8'd220} : s = 295;
	{8'd82,8'd221} : s = 423;
	{8'd82,8'd222} : s = 41;
	{8'd82,8'd223} : s = 147;
	{8'd82,8'd224} : s = 142;
	{8'd82,8'd225} : s = 286;
	{8'd82,8'd226} : s = 141;
	{8'd82,8'd227} : s = 285;
	{8'd82,8'd228} : s = 283;
	{8'd82,8'd229} : s = 414;
	{8'd82,8'd230} : s = 139;
	{8'd82,8'd231} : s = 279;
	{8'd82,8'd232} : s = 271;
	{8'd82,8'd233} : s = 413;
	{8'd82,8'd234} : s = 248;
	{8'd82,8'd235} : s = 411;
	{8'd82,8'd236} : s = 407;
	{8'd82,8'd237} : s = 491;
	{8'd82,8'd238} : s = 5;
	{8'd82,8'd239} : s = 38;
	{8'd82,8'd240} : s = 37;
	{8'd82,8'd241} : s = 135;
	{8'd82,8'd242} : s = 35;
	{8'd82,8'd243} : s = 120;
	{8'd82,8'd244} : s = 116;
	{8'd82,8'd245} : s = 244;
	{8'd82,8'd246} : s = 28;
	{8'd82,8'd247} : s = 114;
	{8'd82,8'd248} : s = 113;
	{8'd82,8'd249} : s = 242;
	{8'd82,8'd250} : s = 108;
	{8'd82,8'd251} : s = 241;
	{8'd82,8'd252} : s = 236;
	{8'd82,8'd253} : s = 399;
	{8'd82,8'd254} : s = 26;
	{8'd82,8'd255} : s = 106;
	{8'd83,8'd0} : s = 389;
	{8'd83,8'd1} : s = 224;
	{8'd83,8'd2} : s = 387;
	{8'd83,8'd3} : s = 368;
	{8'd83,8'd4} : s = 466;
	{8'd83,8'd5} : s = 208;
	{8'd83,8'd6} : s = 360;
	{8'd83,8'd7} : s = 356;
	{8'd83,8'd8} : s = 465;
	{8'd83,8'd9} : s = 354;
	{8'd83,8'd10} : s = 460;
	{8'd83,8'd11} : s = 458;
	{8'd83,8'd12} : s = 500;
	{8'd83,8'd13} : s = 65;
	{8'd83,8'd14} : s = 200;
	{8'd83,8'd15} : s = 196;
	{8'd83,8'd16} : s = 353;
	{8'd83,8'd17} : s = 194;
	{8'd83,8'd18} : s = 344;
	{8'd83,8'd19} : s = 340;
	{8'd83,8'd20} : s = 457;
	{8'd83,8'd21} : s = 193;
	{8'd83,8'd22} : s = 338;
	{8'd83,8'd23} : s = 337;
	{8'd83,8'd24} : s = 454;
	{8'd83,8'd25} : s = 332;
	{8'd83,8'd26} : s = 453;
	{8'd83,8'd27} : s = 451;
	{8'd83,8'd28} : s = 498;
	{8'd83,8'd29} : s = 176;
	{8'd83,8'd30} : s = 330;
	{8'd83,8'd31} : s = 329;
	{8'd83,8'd32} : s = 440;
	{8'd83,8'd33} : s = 326;
	{8'd83,8'd34} : s = 436;
	{8'd83,8'd35} : s = 434;
	{8'd83,8'd36} : s = 497;
	{8'd83,8'd37} : s = 325;
	{8'd83,8'd38} : s = 433;
	{8'd83,8'd39} : s = 428;
	{8'd83,8'd40} : s = 492;
	{8'd83,8'd41} : s = 426;
	{8'd83,8'd42} : s = 490;
	{8'd83,8'd43} : s = 489;
	{8'd83,8'd44} : s = 508;
	{8'd83,8'd45} : s = 2;
	{8'd83,8'd46} : s = 48;
	{8'd83,8'd47} : s = 40;
	{8'd83,8'd48} : s = 168;
	{8'd83,8'd49} : s = 36;
	{8'd83,8'd50} : s = 164;
	{8'd83,8'd51} : s = 162;
	{8'd83,8'd52} : s = 323;
	{8'd83,8'd53} : s = 34;
	{8'd83,8'd54} : s = 161;
	{8'd83,8'd55} : s = 152;
	{8'd83,8'd56} : s = 312;
	{8'd83,8'd57} : s = 148;
	{8'd83,8'd58} : s = 308;
	{8'd83,8'd59} : s = 306;
	{8'd83,8'd60} : s = 425;
	{8'd83,8'd61} : s = 33;
	{8'd83,8'd62} : s = 146;
	{8'd83,8'd63} : s = 145;
	{8'd83,8'd64} : s = 305;
	{8'd83,8'd65} : s = 140;
	{8'd83,8'd66} : s = 300;
	{8'd83,8'd67} : s = 298;
	{8'd83,8'd68} : s = 422;
	{8'd83,8'd69} : s = 138;
	{8'd83,8'd70} : s = 297;
	{8'd83,8'd71} : s = 294;
	{8'd83,8'd72} : s = 421;
	{8'd83,8'd73} : s = 293;
	{8'd83,8'd74} : s = 419;
	{8'd83,8'd75} : s = 412;
	{8'd83,8'd76} : s = 486;
	{8'd83,8'd77} : s = 24;
	{8'd83,8'd78} : s = 137;
	{8'd83,8'd79} : s = 134;
	{8'd83,8'd80} : s = 291;
	{8'd83,8'd81} : s = 133;
	{8'd83,8'd82} : s = 284;
	{8'd83,8'd83} : s = 282;
	{8'd83,8'd84} : s = 410;
	{8'd83,8'd85} : s = 131;
	{8'd83,8'd86} : s = 281;
	{8'd83,8'd87} : s = 278;
	{8'd83,8'd88} : s = 409;
	{8'd83,8'd89} : s = 277;
	{8'd83,8'd90} : s = 406;
	{8'd83,8'd91} : s = 405;
	{8'd83,8'd92} : s = 485;
	{8'd83,8'd93} : s = 112;
	{8'd83,8'd94} : s = 275;
	{8'd83,8'd95} : s = 270;
	{8'd83,8'd96} : s = 403;
	{8'd83,8'd97} : s = 269;
	{8'd83,8'd98} : s = 398;
	{8'd83,8'd99} : s = 397;
	{8'd83,8'd100} : s = 483;
	{8'd83,8'd101} : s = 267;
	{8'd83,8'd102} : s = 395;
	{8'd83,8'd103} : s = 391;
	{8'd83,8'd104} : s = 476;
	{8'd83,8'd105} : s = 376;
	{8'd83,8'd106} : s = 474;
	{8'd83,8'd107} : s = 473;
	{8'd83,8'd108} : s = 506;
	{8'd83,8'd109} : s = 20;
	{8'd83,8'd110} : s = 104;
	{8'd83,8'd111} : s = 100;
	{8'd83,8'd112} : s = 263;
	{8'd83,8'd113} : s = 98;
	{8'd83,8'd114} : s = 240;
	{8'd83,8'd115} : s = 232;
	{8'd83,8'd116} : s = 372;
	{8'd83,8'd117} : s = 97;
	{8'd83,8'd118} : s = 228;
	{8'd83,8'd119} : s = 226;
	{8'd83,8'd120} : s = 370;
	{8'd83,8'd121} : s = 225;
	{8'd83,8'd122} : s = 369;
	{8'd83,8'd123} : s = 364;
	{8'd83,8'd124} : s = 470;
	{8'd83,8'd125} : s = 88;
	{8'd83,8'd126} : s = 216;
	{8'd83,8'd127} : s = 212;
	{8'd83,8'd128} : s = 362;
	{8'd83,8'd129} : s = 210;
	{8'd83,8'd130} : s = 361;
	{8'd83,8'd131} : s = 358;
	{8'd83,8'd132} : s = 469;
	{8'd83,8'd133} : s = 209;
	{8'd83,8'd134} : s = 357;
	{8'd83,8'd135} : s = 355;
	{8'd83,8'd136} : s = 467;
	{8'd83,8'd137} : s = 348;
	{8'd83,8'd138} : s = 462;
	{8'd83,8'd139} : s = 461;
	{8'd83,8'd140} : s = 505;
	{8'd83,8'd141} : s = 84;
	{8'd83,8'd142} : s = 204;
	{8'd83,8'd143} : s = 202;
	{8'd83,8'd144} : s = 346;
	{8'd83,8'd145} : s = 201;
	{8'd83,8'd146} : s = 345;
	{8'd83,8'd147} : s = 342;
	{8'd83,8'd148} : s = 459;
	{8'd83,8'd149} : s = 198;
	{8'd83,8'd150} : s = 341;
	{8'd83,8'd151} : s = 339;
	{8'd83,8'd152} : s = 455;
	{8'd83,8'd153} : s = 334;
	{8'd83,8'd154} : s = 444;
	{8'd83,8'd155} : s = 442;
	{8'd83,8'd156} : s = 502;
	{8'd83,8'd157} : s = 197;
	{8'd83,8'd158} : s = 333;
	{8'd83,8'd159} : s = 331;
	{8'd83,8'd160} : s = 441;
	{8'd83,8'd161} : s = 327;
	{8'd83,8'd162} : s = 438;
	{8'd83,8'd163} : s = 437;
	{8'd83,8'd164} : s = 501;
	{8'd83,8'd165} : s = 316;
	{8'd83,8'd166} : s = 435;
	{8'd83,8'd167} : s = 430;
	{8'd83,8'd168} : s = 499;
	{8'd83,8'd169} : s = 429;
	{8'd83,8'd170} : s = 494;
	{8'd83,8'd171} : s = 493;
	{8'd83,8'd172} : s = 510;
	{8'd83,8'd173} : s = 1;
	{8'd83,8'd174} : s = 18;
	{8'd83,8'd175} : s = 17;
	{8'd83,8'd176} : s = 82;
	{8'd83,8'd177} : s = 12;
	{8'd83,8'd178} : s = 81;
	{8'd83,8'd179} : s = 76;
	{8'd83,8'd180} : s = 195;
	{8'd83,8'd181} : s = 10;
	{8'd83,8'd182} : s = 74;
	{8'd83,8'd183} : s = 73;
	{8'd83,8'd184} : s = 184;
	{8'd83,8'd185} : s = 70;
	{8'd83,8'd186} : s = 180;
	{8'd83,8'd187} : s = 178;
	{8'd83,8'd188} : s = 314;
	{8'd83,8'd189} : s = 9;
	{8'd83,8'd190} : s = 69;
	{8'd83,8'd191} : s = 67;
	{8'd83,8'd192} : s = 177;
	{8'd83,8'd193} : s = 56;
	{8'd83,8'd194} : s = 172;
	{8'd83,8'd195} : s = 170;
	{8'd83,8'd196} : s = 313;
	{8'd83,8'd197} : s = 52;
	{8'd83,8'd198} : s = 169;
	{8'd83,8'd199} : s = 166;
	{8'd83,8'd200} : s = 310;
	{8'd83,8'd201} : s = 165;
	{8'd83,8'd202} : s = 309;
	{8'd83,8'd203} : s = 307;
	{8'd83,8'd204} : s = 427;
	{8'd83,8'd205} : s = 6;
	{8'd83,8'd206} : s = 50;
	{8'd83,8'd207} : s = 49;
	{8'd83,8'd208} : s = 163;
	{8'd83,8'd209} : s = 44;
	{8'd83,8'd210} : s = 156;
	{8'd83,8'd211} : s = 154;
	{8'd83,8'd212} : s = 302;
	{8'd83,8'd213} : s = 42;
	{8'd83,8'd214} : s = 153;
	{8'd83,8'd215} : s = 150;
	{8'd83,8'd216} : s = 301;
	{8'd83,8'd217} : s = 149;
	{8'd83,8'd218} : s = 299;
	{8'd83,8'd219} : s = 295;
	{8'd83,8'd220} : s = 423;
	{8'd83,8'd221} : s = 41;
	{8'd83,8'd222} : s = 147;
	{8'd83,8'd223} : s = 142;
	{8'd83,8'd224} : s = 286;
	{8'd83,8'd225} : s = 141;
	{8'd83,8'd226} : s = 285;
	{8'd83,8'd227} : s = 283;
	{8'd83,8'd228} : s = 414;
	{8'd83,8'd229} : s = 139;
	{8'd83,8'd230} : s = 279;
	{8'd83,8'd231} : s = 271;
	{8'd83,8'd232} : s = 413;
	{8'd83,8'd233} : s = 248;
	{8'd83,8'd234} : s = 411;
	{8'd83,8'd235} : s = 407;
	{8'd83,8'd236} : s = 491;
	{8'd83,8'd237} : s = 5;
	{8'd83,8'd238} : s = 38;
	{8'd83,8'd239} : s = 37;
	{8'd83,8'd240} : s = 135;
	{8'd83,8'd241} : s = 35;
	{8'd83,8'd242} : s = 120;
	{8'd83,8'd243} : s = 116;
	{8'd83,8'd244} : s = 244;
	{8'd83,8'd245} : s = 28;
	{8'd83,8'd246} : s = 114;
	{8'd83,8'd247} : s = 113;
	{8'd83,8'd248} : s = 242;
	{8'd83,8'd249} : s = 108;
	{8'd83,8'd250} : s = 241;
	{8'd83,8'd251} : s = 236;
	{8'd83,8'd252} : s = 399;
	{8'd83,8'd253} : s = 26;
	{8'd83,8'd254} : s = 106;
	{8'd83,8'd255} : s = 105;
	{8'd84,8'd0} : s = 224;
	{8'd84,8'd1} : s = 387;
	{8'd84,8'd2} : s = 368;
	{8'd84,8'd3} : s = 466;
	{8'd84,8'd4} : s = 208;
	{8'd84,8'd5} : s = 360;
	{8'd84,8'd6} : s = 356;
	{8'd84,8'd7} : s = 465;
	{8'd84,8'd8} : s = 354;
	{8'd84,8'd9} : s = 460;
	{8'd84,8'd10} : s = 458;
	{8'd84,8'd11} : s = 500;
	{8'd84,8'd12} : s = 65;
	{8'd84,8'd13} : s = 200;
	{8'd84,8'd14} : s = 196;
	{8'd84,8'd15} : s = 353;
	{8'd84,8'd16} : s = 194;
	{8'd84,8'd17} : s = 344;
	{8'd84,8'd18} : s = 340;
	{8'd84,8'd19} : s = 457;
	{8'd84,8'd20} : s = 193;
	{8'd84,8'd21} : s = 338;
	{8'd84,8'd22} : s = 337;
	{8'd84,8'd23} : s = 454;
	{8'd84,8'd24} : s = 332;
	{8'd84,8'd25} : s = 453;
	{8'd84,8'd26} : s = 451;
	{8'd84,8'd27} : s = 498;
	{8'd84,8'd28} : s = 176;
	{8'd84,8'd29} : s = 330;
	{8'd84,8'd30} : s = 329;
	{8'd84,8'd31} : s = 440;
	{8'd84,8'd32} : s = 326;
	{8'd84,8'd33} : s = 436;
	{8'd84,8'd34} : s = 434;
	{8'd84,8'd35} : s = 497;
	{8'd84,8'd36} : s = 325;
	{8'd84,8'd37} : s = 433;
	{8'd84,8'd38} : s = 428;
	{8'd84,8'd39} : s = 492;
	{8'd84,8'd40} : s = 426;
	{8'd84,8'd41} : s = 490;
	{8'd84,8'd42} : s = 489;
	{8'd84,8'd43} : s = 508;
	{8'd84,8'd44} : s = 2;
	{8'd84,8'd45} : s = 48;
	{8'd84,8'd46} : s = 40;
	{8'd84,8'd47} : s = 168;
	{8'd84,8'd48} : s = 36;
	{8'd84,8'd49} : s = 164;
	{8'd84,8'd50} : s = 162;
	{8'd84,8'd51} : s = 323;
	{8'd84,8'd52} : s = 34;
	{8'd84,8'd53} : s = 161;
	{8'd84,8'd54} : s = 152;
	{8'd84,8'd55} : s = 312;
	{8'd84,8'd56} : s = 148;
	{8'd84,8'd57} : s = 308;
	{8'd84,8'd58} : s = 306;
	{8'd84,8'd59} : s = 425;
	{8'd84,8'd60} : s = 33;
	{8'd84,8'd61} : s = 146;
	{8'd84,8'd62} : s = 145;
	{8'd84,8'd63} : s = 305;
	{8'd84,8'd64} : s = 140;
	{8'd84,8'd65} : s = 300;
	{8'd84,8'd66} : s = 298;
	{8'd84,8'd67} : s = 422;
	{8'd84,8'd68} : s = 138;
	{8'd84,8'd69} : s = 297;
	{8'd84,8'd70} : s = 294;
	{8'd84,8'd71} : s = 421;
	{8'd84,8'd72} : s = 293;
	{8'd84,8'd73} : s = 419;
	{8'd84,8'd74} : s = 412;
	{8'd84,8'd75} : s = 486;
	{8'd84,8'd76} : s = 24;
	{8'd84,8'd77} : s = 137;
	{8'd84,8'd78} : s = 134;
	{8'd84,8'd79} : s = 291;
	{8'd84,8'd80} : s = 133;
	{8'd84,8'd81} : s = 284;
	{8'd84,8'd82} : s = 282;
	{8'd84,8'd83} : s = 410;
	{8'd84,8'd84} : s = 131;
	{8'd84,8'd85} : s = 281;
	{8'd84,8'd86} : s = 278;
	{8'd84,8'd87} : s = 409;
	{8'd84,8'd88} : s = 277;
	{8'd84,8'd89} : s = 406;
	{8'd84,8'd90} : s = 405;
	{8'd84,8'd91} : s = 485;
	{8'd84,8'd92} : s = 112;
	{8'd84,8'd93} : s = 275;
	{8'd84,8'd94} : s = 270;
	{8'd84,8'd95} : s = 403;
	{8'd84,8'd96} : s = 269;
	{8'd84,8'd97} : s = 398;
	{8'd84,8'd98} : s = 397;
	{8'd84,8'd99} : s = 483;
	{8'd84,8'd100} : s = 267;
	{8'd84,8'd101} : s = 395;
	{8'd84,8'd102} : s = 391;
	{8'd84,8'd103} : s = 476;
	{8'd84,8'd104} : s = 376;
	{8'd84,8'd105} : s = 474;
	{8'd84,8'd106} : s = 473;
	{8'd84,8'd107} : s = 506;
	{8'd84,8'd108} : s = 20;
	{8'd84,8'd109} : s = 104;
	{8'd84,8'd110} : s = 100;
	{8'd84,8'd111} : s = 263;
	{8'd84,8'd112} : s = 98;
	{8'd84,8'd113} : s = 240;
	{8'd84,8'd114} : s = 232;
	{8'd84,8'd115} : s = 372;
	{8'd84,8'd116} : s = 97;
	{8'd84,8'd117} : s = 228;
	{8'd84,8'd118} : s = 226;
	{8'd84,8'd119} : s = 370;
	{8'd84,8'd120} : s = 225;
	{8'd84,8'd121} : s = 369;
	{8'd84,8'd122} : s = 364;
	{8'd84,8'd123} : s = 470;
	{8'd84,8'd124} : s = 88;
	{8'd84,8'd125} : s = 216;
	{8'd84,8'd126} : s = 212;
	{8'd84,8'd127} : s = 362;
	{8'd84,8'd128} : s = 210;
	{8'd84,8'd129} : s = 361;
	{8'd84,8'd130} : s = 358;
	{8'd84,8'd131} : s = 469;
	{8'd84,8'd132} : s = 209;
	{8'd84,8'd133} : s = 357;
	{8'd84,8'd134} : s = 355;
	{8'd84,8'd135} : s = 467;
	{8'd84,8'd136} : s = 348;
	{8'd84,8'd137} : s = 462;
	{8'd84,8'd138} : s = 461;
	{8'd84,8'd139} : s = 505;
	{8'd84,8'd140} : s = 84;
	{8'd84,8'd141} : s = 204;
	{8'd84,8'd142} : s = 202;
	{8'd84,8'd143} : s = 346;
	{8'd84,8'd144} : s = 201;
	{8'd84,8'd145} : s = 345;
	{8'd84,8'd146} : s = 342;
	{8'd84,8'd147} : s = 459;
	{8'd84,8'd148} : s = 198;
	{8'd84,8'd149} : s = 341;
	{8'd84,8'd150} : s = 339;
	{8'd84,8'd151} : s = 455;
	{8'd84,8'd152} : s = 334;
	{8'd84,8'd153} : s = 444;
	{8'd84,8'd154} : s = 442;
	{8'd84,8'd155} : s = 502;
	{8'd84,8'd156} : s = 197;
	{8'd84,8'd157} : s = 333;
	{8'd84,8'd158} : s = 331;
	{8'd84,8'd159} : s = 441;
	{8'd84,8'd160} : s = 327;
	{8'd84,8'd161} : s = 438;
	{8'd84,8'd162} : s = 437;
	{8'd84,8'd163} : s = 501;
	{8'd84,8'd164} : s = 316;
	{8'd84,8'd165} : s = 435;
	{8'd84,8'd166} : s = 430;
	{8'd84,8'd167} : s = 499;
	{8'd84,8'd168} : s = 429;
	{8'd84,8'd169} : s = 494;
	{8'd84,8'd170} : s = 493;
	{8'd84,8'd171} : s = 510;
	{8'd84,8'd172} : s = 1;
	{8'd84,8'd173} : s = 18;
	{8'd84,8'd174} : s = 17;
	{8'd84,8'd175} : s = 82;
	{8'd84,8'd176} : s = 12;
	{8'd84,8'd177} : s = 81;
	{8'd84,8'd178} : s = 76;
	{8'd84,8'd179} : s = 195;
	{8'd84,8'd180} : s = 10;
	{8'd84,8'd181} : s = 74;
	{8'd84,8'd182} : s = 73;
	{8'd84,8'd183} : s = 184;
	{8'd84,8'd184} : s = 70;
	{8'd84,8'd185} : s = 180;
	{8'd84,8'd186} : s = 178;
	{8'd84,8'd187} : s = 314;
	{8'd84,8'd188} : s = 9;
	{8'd84,8'd189} : s = 69;
	{8'd84,8'd190} : s = 67;
	{8'd84,8'd191} : s = 177;
	{8'd84,8'd192} : s = 56;
	{8'd84,8'd193} : s = 172;
	{8'd84,8'd194} : s = 170;
	{8'd84,8'd195} : s = 313;
	{8'd84,8'd196} : s = 52;
	{8'd84,8'd197} : s = 169;
	{8'd84,8'd198} : s = 166;
	{8'd84,8'd199} : s = 310;
	{8'd84,8'd200} : s = 165;
	{8'd84,8'd201} : s = 309;
	{8'd84,8'd202} : s = 307;
	{8'd84,8'd203} : s = 427;
	{8'd84,8'd204} : s = 6;
	{8'd84,8'd205} : s = 50;
	{8'd84,8'd206} : s = 49;
	{8'd84,8'd207} : s = 163;
	{8'd84,8'd208} : s = 44;
	{8'd84,8'd209} : s = 156;
	{8'd84,8'd210} : s = 154;
	{8'd84,8'd211} : s = 302;
	{8'd84,8'd212} : s = 42;
	{8'd84,8'd213} : s = 153;
	{8'd84,8'd214} : s = 150;
	{8'd84,8'd215} : s = 301;
	{8'd84,8'd216} : s = 149;
	{8'd84,8'd217} : s = 299;
	{8'd84,8'd218} : s = 295;
	{8'd84,8'd219} : s = 423;
	{8'd84,8'd220} : s = 41;
	{8'd84,8'd221} : s = 147;
	{8'd84,8'd222} : s = 142;
	{8'd84,8'd223} : s = 286;
	{8'd84,8'd224} : s = 141;
	{8'd84,8'd225} : s = 285;
	{8'd84,8'd226} : s = 283;
	{8'd84,8'd227} : s = 414;
	{8'd84,8'd228} : s = 139;
	{8'd84,8'd229} : s = 279;
	{8'd84,8'd230} : s = 271;
	{8'd84,8'd231} : s = 413;
	{8'd84,8'd232} : s = 248;
	{8'd84,8'd233} : s = 411;
	{8'd84,8'd234} : s = 407;
	{8'd84,8'd235} : s = 491;
	{8'd84,8'd236} : s = 5;
	{8'd84,8'd237} : s = 38;
	{8'd84,8'd238} : s = 37;
	{8'd84,8'd239} : s = 135;
	{8'd84,8'd240} : s = 35;
	{8'd84,8'd241} : s = 120;
	{8'd84,8'd242} : s = 116;
	{8'd84,8'd243} : s = 244;
	{8'd84,8'd244} : s = 28;
	{8'd84,8'd245} : s = 114;
	{8'd84,8'd246} : s = 113;
	{8'd84,8'd247} : s = 242;
	{8'd84,8'd248} : s = 108;
	{8'd84,8'd249} : s = 241;
	{8'd84,8'd250} : s = 236;
	{8'd84,8'd251} : s = 399;
	{8'd84,8'd252} : s = 26;
	{8'd84,8'd253} : s = 106;
	{8'd84,8'd254} : s = 105;
	{8'd84,8'd255} : s = 234;
	{8'd85,8'd0} : s = 387;
	{8'd85,8'd1} : s = 368;
	{8'd85,8'd2} : s = 466;
	{8'd85,8'd3} : s = 208;
	{8'd85,8'd4} : s = 360;
	{8'd85,8'd5} : s = 356;
	{8'd85,8'd6} : s = 465;
	{8'd85,8'd7} : s = 354;
	{8'd85,8'd8} : s = 460;
	{8'd85,8'd9} : s = 458;
	{8'd85,8'd10} : s = 500;
	{8'd85,8'd11} : s = 65;
	{8'd85,8'd12} : s = 200;
	{8'd85,8'd13} : s = 196;
	{8'd85,8'd14} : s = 353;
	{8'd85,8'd15} : s = 194;
	{8'd85,8'd16} : s = 344;
	{8'd85,8'd17} : s = 340;
	{8'd85,8'd18} : s = 457;
	{8'd85,8'd19} : s = 193;
	{8'd85,8'd20} : s = 338;
	{8'd85,8'd21} : s = 337;
	{8'd85,8'd22} : s = 454;
	{8'd85,8'd23} : s = 332;
	{8'd85,8'd24} : s = 453;
	{8'd85,8'd25} : s = 451;
	{8'd85,8'd26} : s = 498;
	{8'd85,8'd27} : s = 176;
	{8'd85,8'd28} : s = 330;
	{8'd85,8'd29} : s = 329;
	{8'd85,8'd30} : s = 440;
	{8'd85,8'd31} : s = 326;
	{8'd85,8'd32} : s = 436;
	{8'd85,8'd33} : s = 434;
	{8'd85,8'd34} : s = 497;
	{8'd85,8'd35} : s = 325;
	{8'd85,8'd36} : s = 433;
	{8'd85,8'd37} : s = 428;
	{8'd85,8'd38} : s = 492;
	{8'd85,8'd39} : s = 426;
	{8'd85,8'd40} : s = 490;
	{8'd85,8'd41} : s = 489;
	{8'd85,8'd42} : s = 508;
	{8'd85,8'd43} : s = 2;
	{8'd85,8'd44} : s = 48;
	{8'd85,8'd45} : s = 40;
	{8'd85,8'd46} : s = 168;
	{8'd85,8'd47} : s = 36;
	{8'd85,8'd48} : s = 164;
	{8'd85,8'd49} : s = 162;
	{8'd85,8'd50} : s = 323;
	{8'd85,8'd51} : s = 34;
	{8'd85,8'd52} : s = 161;
	{8'd85,8'd53} : s = 152;
	{8'd85,8'd54} : s = 312;
	{8'd85,8'd55} : s = 148;
	{8'd85,8'd56} : s = 308;
	{8'd85,8'd57} : s = 306;
	{8'd85,8'd58} : s = 425;
	{8'd85,8'd59} : s = 33;
	{8'd85,8'd60} : s = 146;
	{8'd85,8'd61} : s = 145;
	{8'd85,8'd62} : s = 305;
	{8'd85,8'd63} : s = 140;
	{8'd85,8'd64} : s = 300;
	{8'd85,8'd65} : s = 298;
	{8'd85,8'd66} : s = 422;
	{8'd85,8'd67} : s = 138;
	{8'd85,8'd68} : s = 297;
	{8'd85,8'd69} : s = 294;
	{8'd85,8'd70} : s = 421;
	{8'd85,8'd71} : s = 293;
	{8'd85,8'd72} : s = 419;
	{8'd85,8'd73} : s = 412;
	{8'd85,8'd74} : s = 486;
	{8'd85,8'd75} : s = 24;
	{8'd85,8'd76} : s = 137;
	{8'd85,8'd77} : s = 134;
	{8'd85,8'd78} : s = 291;
	{8'd85,8'd79} : s = 133;
	{8'd85,8'd80} : s = 284;
	{8'd85,8'd81} : s = 282;
	{8'd85,8'd82} : s = 410;
	{8'd85,8'd83} : s = 131;
	{8'd85,8'd84} : s = 281;
	{8'd85,8'd85} : s = 278;
	{8'd85,8'd86} : s = 409;
	{8'd85,8'd87} : s = 277;
	{8'd85,8'd88} : s = 406;
	{8'd85,8'd89} : s = 405;
	{8'd85,8'd90} : s = 485;
	{8'd85,8'd91} : s = 112;
	{8'd85,8'd92} : s = 275;
	{8'd85,8'd93} : s = 270;
	{8'd85,8'd94} : s = 403;
	{8'd85,8'd95} : s = 269;
	{8'd85,8'd96} : s = 398;
	{8'd85,8'd97} : s = 397;
	{8'd85,8'd98} : s = 483;
	{8'd85,8'd99} : s = 267;
	{8'd85,8'd100} : s = 395;
	{8'd85,8'd101} : s = 391;
	{8'd85,8'd102} : s = 476;
	{8'd85,8'd103} : s = 376;
	{8'd85,8'd104} : s = 474;
	{8'd85,8'd105} : s = 473;
	{8'd85,8'd106} : s = 506;
	{8'd85,8'd107} : s = 20;
	{8'd85,8'd108} : s = 104;
	{8'd85,8'd109} : s = 100;
	{8'd85,8'd110} : s = 263;
	{8'd85,8'd111} : s = 98;
	{8'd85,8'd112} : s = 240;
	{8'd85,8'd113} : s = 232;
	{8'd85,8'd114} : s = 372;
	{8'd85,8'd115} : s = 97;
	{8'd85,8'd116} : s = 228;
	{8'd85,8'd117} : s = 226;
	{8'd85,8'd118} : s = 370;
	{8'd85,8'd119} : s = 225;
	{8'd85,8'd120} : s = 369;
	{8'd85,8'd121} : s = 364;
	{8'd85,8'd122} : s = 470;
	{8'd85,8'd123} : s = 88;
	{8'd85,8'd124} : s = 216;
	{8'd85,8'd125} : s = 212;
	{8'd85,8'd126} : s = 362;
	{8'd85,8'd127} : s = 210;
	{8'd85,8'd128} : s = 361;
	{8'd85,8'd129} : s = 358;
	{8'd85,8'd130} : s = 469;
	{8'd85,8'd131} : s = 209;
	{8'd85,8'd132} : s = 357;
	{8'd85,8'd133} : s = 355;
	{8'd85,8'd134} : s = 467;
	{8'd85,8'd135} : s = 348;
	{8'd85,8'd136} : s = 462;
	{8'd85,8'd137} : s = 461;
	{8'd85,8'd138} : s = 505;
	{8'd85,8'd139} : s = 84;
	{8'd85,8'd140} : s = 204;
	{8'd85,8'd141} : s = 202;
	{8'd85,8'd142} : s = 346;
	{8'd85,8'd143} : s = 201;
	{8'd85,8'd144} : s = 345;
	{8'd85,8'd145} : s = 342;
	{8'd85,8'd146} : s = 459;
	{8'd85,8'd147} : s = 198;
	{8'd85,8'd148} : s = 341;
	{8'd85,8'd149} : s = 339;
	{8'd85,8'd150} : s = 455;
	{8'd85,8'd151} : s = 334;
	{8'd85,8'd152} : s = 444;
	{8'd85,8'd153} : s = 442;
	{8'd85,8'd154} : s = 502;
	{8'd85,8'd155} : s = 197;
	{8'd85,8'd156} : s = 333;
	{8'd85,8'd157} : s = 331;
	{8'd85,8'd158} : s = 441;
	{8'd85,8'd159} : s = 327;
	{8'd85,8'd160} : s = 438;
	{8'd85,8'd161} : s = 437;
	{8'd85,8'd162} : s = 501;
	{8'd85,8'd163} : s = 316;
	{8'd85,8'd164} : s = 435;
	{8'd85,8'd165} : s = 430;
	{8'd85,8'd166} : s = 499;
	{8'd85,8'd167} : s = 429;
	{8'd85,8'd168} : s = 494;
	{8'd85,8'd169} : s = 493;
	{8'd85,8'd170} : s = 510;
	{8'd85,8'd171} : s = 1;
	{8'd85,8'd172} : s = 18;
	{8'd85,8'd173} : s = 17;
	{8'd85,8'd174} : s = 82;
	{8'd85,8'd175} : s = 12;
	{8'd85,8'd176} : s = 81;
	{8'd85,8'd177} : s = 76;
	{8'd85,8'd178} : s = 195;
	{8'd85,8'd179} : s = 10;
	{8'd85,8'd180} : s = 74;
	{8'd85,8'd181} : s = 73;
	{8'd85,8'd182} : s = 184;
	{8'd85,8'd183} : s = 70;
	{8'd85,8'd184} : s = 180;
	{8'd85,8'd185} : s = 178;
	{8'd85,8'd186} : s = 314;
	{8'd85,8'd187} : s = 9;
	{8'd85,8'd188} : s = 69;
	{8'd85,8'd189} : s = 67;
	{8'd85,8'd190} : s = 177;
	{8'd85,8'd191} : s = 56;
	{8'd85,8'd192} : s = 172;
	{8'd85,8'd193} : s = 170;
	{8'd85,8'd194} : s = 313;
	{8'd85,8'd195} : s = 52;
	{8'd85,8'd196} : s = 169;
	{8'd85,8'd197} : s = 166;
	{8'd85,8'd198} : s = 310;
	{8'd85,8'd199} : s = 165;
	{8'd85,8'd200} : s = 309;
	{8'd85,8'd201} : s = 307;
	{8'd85,8'd202} : s = 427;
	{8'd85,8'd203} : s = 6;
	{8'd85,8'd204} : s = 50;
	{8'd85,8'd205} : s = 49;
	{8'd85,8'd206} : s = 163;
	{8'd85,8'd207} : s = 44;
	{8'd85,8'd208} : s = 156;
	{8'd85,8'd209} : s = 154;
	{8'd85,8'd210} : s = 302;
	{8'd85,8'd211} : s = 42;
	{8'd85,8'd212} : s = 153;
	{8'd85,8'd213} : s = 150;
	{8'd85,8'd214} : s = 301;
	{8'd85,8'd215} : s = 149;
	{8'd85,8'd216} : s = 299;
	{8'd85,8'd217} : s = 295;
	{8'd85,8'd218} : s = 423;
	{8'd85,8'd219} : s = 41;
	{8'd85,8'd220} : s = 147;
	{8'd85,8'd221} : s = 142;
	{8'd85,8'd222} : s = 286;
	{8'd85,8'd223} : s = 141;
	{8'd85,8'd224} : s = 285;
	{8'd85,8'd225} : s = 283;
	{8'd85,8'd226} : s = 414;
	{8'd85,8'd227} : s = 139;
	{8'd85,8'd228} : s = 279;
	{8'd85,8'd229} : s = 271;
	{8'd85,8'd230} : s = 413;
	{8'd85,8'd231} : s = 248;
	{8'd85,8'd232} : s = 411;
	{8'd85,8'd233} : s = 407;
	{8'd85,8'd234} : s = 491;
	{8'd85,8'd235} : s = 5;
	{8'd85,8'd236} : s = 38;
	{8'd85,8'd237} : s = 37;
	{8'd85,8'd238} : s = 135;
	{8'd85,8'd239} : s = 35;
	{8'd85,8'd240} : s = 120;
	{8'd85,8'd241} : s = 116;
	{8'd85,8'd242} : s = 244;
	{8'd85,8'd243} : s = 28;
	{8'd85,8'd244} : s = 114;
	{8'd85,8'd245} : s = 113;
	{8'd85,8'd246} : s = 242;
	{8'd85,8'd247} : s = 108;
	{8'd85,8'd248} : s = 241;
	{8'd85,8'd249} : s = 236;
	{8'd85,8'd250} : s = 399;
	{8'd85,8'd251} : s = 26;
	{8'd85,8'd252} : s = 106;
	{8'd85,8'd253} : s = 105;
	{8'd85,8'd254} : s = 234;
	{8'd85,8'd255} : s = 102;
	{8'd86,8'd0} : s = 368;
	{8'd86,8'd1} : s = 466;
	{8'd86,8'd2} : s = 208;
	{8'd86,8'd3} : s = 360;
	{8'd86,8'd4} : s = 356;
	{8'd86,8'd5} : s = 465;
	{8'd86,8'd6} : s = 354;
	{8'd86,8'd7} : s = 460;
	{8'd86,8'd8} : s = 458;
	{8'd86,8'd9} : s = 500;
	{8'd86,8'd10} : s = 65;
	{8'd86,8'd11} : s = 200;
	{8'd86,8'd12} : s = 196;
	{8'd86,8'd13} : s = 353;
	{8'd86,8'd14} : s = 194;
	{8'd86,8'd15} : s = 344;
	{8'd86,8'd16} : s = 340;
	{8'd86,8'd17} : s = 457;
	{8'd86,8'd18} : s = 193;
	{8'd86,8'd19} : s = 338;
	{8'd86,8'd20} : s = 337;
	{8'd86,8'd21} : s = 454;
	{8'd86,8'd22} : s = 332;
	{8'd86,8'd23} : s = 453;
	{8'd86,8'd24} : s = 451;
	{8'd86,8'd25} : s = 498;
	{8'd86,8'd26} : s = 176;
	{8'd86,8'd27} : s = 330;
	{8'd86,8'd28} : s = 329;
	{8'd86,8'd29} : s = 440;
	{8'd86,8'd30} : s = 326;
	{8'd86,8'd31} : s = 436;
	{8'd86,8'd32} : s = 434;
	{8'd86,8'd33} : s = 497;
	{8'd86,8'd34} : s = 325;
	{8'd86,8'd35} : s = 433;
	{8'd86,8'd36} : s = 428;
	{8'd86,8'd37} : s = 492;
	{8'd86,8'd38} : s = 426;
	{8'd86,8'd39} : s = 490;
	{8'd86,8'd40} : s = 489;
	{8'd86,8'd41} : s = 508;
	{8'd86,8'd42} : s = 2;
	{8'd86,8'd43} : s = 48;
	{8'd86,8'd44} : s = 40;
	{8'd86,8'd45} : s = 168;
	{8'd86,8'd46} : s = 36;
	{8'd86,8'd47} : s = 164;
	{8'd86,8'd48} : s = 162;
	{8'd86,8'd49} : s = 323;
	{8'd86,8'd50} : s = 34;
	{8'd86,8'd51} : s = 161;
	{8'd86,8'd52} : s = 152;
	{8'd86,8'd53} : s = 312;
	{8'd86,8'd54} : s = 148;
	{8'd86,8'd55} : s = 308;
	{8'd86,8'd56} : s = 306;
	{8'd86,8'd57} : s = 425;
	{8'd86,8'd58} : s = 33;
	{8'd86,8'd59} : s = 146;
	{8'd86,8'd60} : s = 145;
	{8'd86,8'd61} : s = 305;
	{8'd86,8'd62} : s = 140;
	{8'd86,8'd63} : s = 300;
	{8'd86,8'd64} : s = 298;
	{8'd86,8'd65} : s = 422;
	{8'd86,8'd66} : s = 138;
	{8'd86,8'd67} : s = 297;
	{8'd86,8'd68} : s = 294;
	{8'd86,8'd69} : s = 421;
	{8'd86,8'd70} : s = 293;
	{8'd86,8'd71} : s = 419;
	{8'd86,8'd72} : s = 412;
	{8'd86,8'd73} : s = 486;
	{8'd86,8'd74} : s = 24;
	{8'd86,8'd75} : s = 137;
	{8'd86,8'd76} : s = 134;
	{8'd86,8'd77} : s = 291;
	{8'd86,8'd78} : s = 133;
	{8'd86,8'd79} : s = 284;
	{8'd86,8'd80} : s = 282;
	{8'd86,8'd81} : s = 410;
	{8'd86,8'd82} : s = 131;
	{8'd86,8'd83} : s = 281;
	{8'd86,8'd84} : s = 278;
	{8'd86,8'd85} : s = 409;
	{8'd86,8'd86} : s = 277;
	{8'd86,8'd87} : s = 406;
	{8'd86,8'd88} : s = 405;
	{8'd86,8'd89} : s = 485;
	{8'd86,8'd90} : s = 112;
	{8'd86,8'd91} : s = 275;
	{8'd86,8'd92} : s = 270;
	{8'd86,8'd93} : s = 403;
	{8'd86,8'd94} : s = 269;
	{8'd86,8'd95} : s = 398;
	{8'd86,8'd96} : s = 397;
	{8'd86,8'd97} : s = 483;
	{8'd86,8'd98} : s = 267;
	{8'd86,8'd99} : s = 395;
	{8'd86,8'd100} : s = 391;
	{8'd86,8'd101} : s = 476;
	{8'd86,8'd102} : s = 376;
	{8'd86,8'd103} : s = 474;
	{8'd86,8'd104} : s = 473;
	{8'd86,8'd105} : s = 506;
	{8'd86,8'd106} : s = 20;
	{8'd86,8'd107} : s = 104;
	{8'd86,8'd108} : s = 100;
	{8'd86,8'd109} : s = 263;
	{8'd86,8'd110} : s = 98;
	{8'd86,8'd111} : s = 240;
	{8'd86,8'd112} : s = 232;
	{8'd86,8'd113} : s = 372;
	{8'd86,8'd114} : s = 97;
	{8'd86,8'd115} : s = 228;
	{8'd86,8'd116} : s = 226;
	{8'd86,8'd117} : s = 370;
	{8'd86,8'd118} : s = 225;
	{8'd86,8'd119} : s = 369;
	{8'd86,8'd120} : s = 364;
	{8'd86,8'd121} : s = 470;
	{8'd86,8'd122} : s = 88;
	{8'd86,8'd123} : s = 216;
	{8'd86,8'd124} : s = 212;
	{8'd86,8'd125} : s = 362;
	{8'd86,8'd126} : s = 210;
	{8'd86,8'd127} : s = 361;
	{8'd86,8'd128} : s = 358;
	{8'd86,8'd129} : s = 469;
	{8'd86,8'd130} : s = 209;
	{8'd86,8'd131} : s = 357;
	{8'd86,8'd132} : s = 355;
	{8'd86,8'd133} : s = 467;
	{8'd86,8'd134} : s = 348;
	{8'd86,8'd135} : s = 462;
	{8'd86,8'd136} : s = 461;
	{8'd86,8'd137} : s = 505;
	{8'd86,8'd138} : s = 84;
	{8'd86,8'd139} : s = 204;
	{8'd86,8'd140} : s = 202;
	{8'd86,8'd141} : s = 346;
	{8'd86,8'd142} : s = 201;
	{8'd86,8'd143} : s = 345;
	{8'd86,8'd144} : s = 342;
	{8'd86,8'd145} : s = 459;
	{8'd86,8'd146} : s = 198;
	{8'd86,8'd147} : s = 341;
	{8'd86,8'd148} : s = 339;
	{8'd86,8'd149} : s = 455;
	{8'd86,8'd150} : s = 334;
	{8'd86,8'd151} : s = 444;
	{8'd86,8'd152} : s = 442;
	{8'd86,8'd153} : s = 502;
	{8'd86,8'd154} : s = 197;
	{8'd86,8'd155} : s = 333;
	{8'd86,8'd156} : s = 331;
	{8'd86,8'd157} : s = 441;
	{8'd86,8'd158} : s = 327;
	{8'd86,8'd159} : s = 438;
	{8'd86,8'd160} : s = 437;
	{8'd86,8'd161} : s = 501;
	{8'd86,8'd162} : s = 316;
	{8'd86,8'd163} : s = 435;
	{8'd86,8'd164} : s = 430;
	{8'd86,8'd165} : s = 499;
	{8'd86,8'd166} : s = 429;
	{8'd86,8'd167} : s = 494;
	{8'd86,8'd168} : s = 493;
	{8'd86,8'd169} : s = 510;
	{8'd86,8'd170} : s = 1;
	{8'd86,8'd171} : s = 18;
	{8'd86,8'd172} : s = 17;
	{8'd86,8'd173} : s = 82;
	{8'd86,8'd174} : s = 12;
	{8'd86,8'd175} : s = 81;
	{8'd86,8'd176} : s = 76;
	{8'd86,8'd177} : s = 195;
	{8'd86,8'd178} : s = 10;
	{8'd86,8'd179} : s = 74;
	{8'd86,8'd180} : s = 73;
	{8'd86,8'd181} : s = 184;
	{8'd86,8'd182} : s = 70;
	{8'd86,8'd183} : s = 180;
	{8'd86,8'd184} : s = 178;
	{8'd86,8'd185} : s = 314;
	{8'd86,8'd186} : s = 9;
	{8'd86,8'd187} : s = 69;
	{8'd86,8'd188} : s = 67;
	{8'd86,8'd189} : s = 177;
	{8'd86,8'd190} : s = 56;
	{8'd86,8'd191} : s = 172;
	{8'd86,8'd192} : s = 170;
	{8'd86,8'd193} : s = 313;
	{8'd86,8'd194} : s = 52;
	{8'd86,8'd195} : s = 169;
	{8'd86,8'd196} : s = 166;
	{8'd86,8'd197} : s = 310;
	{8'd86,8'd198} : s = 165;
	{8'd86,8'd199} : s = 309;
	{8'd86,8'd200} : s = 307;
	{8'd86,8'd201} : s = 427;
	{8'd86,8'd202} : s = 6;
	{8'd86,8'd203} : s = 50;
	{8'd86,8'd204} : s = 49;
	{8'd86,8'd205} : s = 163;
	{8'd86,8'd206} : s = 44;
	{8'd86,8'd207} : s = 156;
	{8'd86,8'd208} : s = 154;
	{8'd86,8'd209} : s = 302;
	{8'd86,8'd210} : s = 42;
	{8'd86,8'd211} : s = 153;
	{8'd86,8'd212} : s = 150;
	{8'd86,8'd213} : s = 301;
	{8'd86,8'd214} : s = 149;
	{8'd86,8'd215} : s = 299;
	{8'd86,8'd216} : s = 295;
	{8'd86,8'd217} : s = 423;
	{8'd86,8'd218} : s = 41;
	{8'd86,8'd219} : s = 147;
	{8'd86,8'd220} : s = 142;
	{8'd86,8'd221} : s = 286;
	{8'd86,8'd222} : s = 141;
	{8'd86,8'd223} : s = 285;
	{8'd86,8'd224} : s = 283;
	{8'd86,8'd225} : s = 414;
	{8'd86,8'd226} : s = 139;
	{8'd86,8'd227} : s = 279;
	{8'd86,8'd228} : s = 271;
	{8'd86,8'd229} : s = 413;
	{8'd86,8'd230} : s = 248;
	{8'd86,8'd231} : s = 411;
	{8'd86,8'd232} : s = 407;
	{8'd86,8'd233} : s = 491;
	{8'd86,8'd234} : s = 5;
	{8'd86,8'd235} : s = 38;
	{8'd86,8'd236} : s = 37;
	{8'd86,8'd237} : s = 135;
	{8'd86,8'd238} : s = 35;
	{8'd86,8'd239} : s = 120;
	{8'd86,8'd240} : s = 116;
	{8'd86,8'd241} : s = 244;
	{8'd86,8'd242} : s = 28;
	{8'd86,8'd243} : s = 114;
	{8'd86,8'd244} : s = 113;
	{8'd86,8'd245} : s = 242;
	{8'd86,8'd246} : s = 108;
	{8'd86,8'd247} : s = 241;
	{8'd86,8'd248} : s = 236;
	{8'd86,8'd249} : s = 399;
	{8'd86,8'd250} : s = 26;
	{8'd86,8'd251} : s = 106;
	{8'd86,8'd252} : s = 105;
	{8'd86,8'd253} : s = 234;
	{8'd86,8'd254} : s = 102;
	{8'd86,8'd255} : s = 233;
	{8'd87,8'd0} : s = 466;
	{8'd87,8'd1} : s = 208;
	{8'd87,8'd2} : s = 360;
	{8'd87,8'd3} : s = 356;
	{8'd87,8'd4} : s = 465;
	{8'd87,8'd5} : s = 354;
	{8'd87,8'd6} : s = 460;
	{8'd87,8'd7} : s = 458;
	{8'd87,8'd8} : s = 500;
	{8'd87,8'd9} : s = 65;
	{8'd87,8'd10} : s = 200;
	{8'd87,8'd11} : s = 196;
	{8'd87,8'd12} : s = 353;
	{8'd87,8'd13} : s = 194;
	{8'd87,8'd14} : s = 344;
	{8'd87,8'd15} : s = 340;
	{8'd87,8'd16} : s = 457;
	{8'd87,8'd17} : s = 193;
	{8'd87,8'd18} : s = 338;
	{8'd87,8'd19} : s = 337;
	{8'd87,8'd20} : s = 454;
	{8'd87,8'd21} : s = 332;
	{8'd87,8'd22} : s = 453;
	{8'd87,8'd23} : s = 451;
	{8'd87,8'd24} : s = 498;
	{8'd87,8'd25} : s = 176;
	{8'd87,8'd26} : s = 330;
	{8'd87,8'd27} : s = 329;
	{8'd87,8'd28} : s = 440;
	{8'd87,8'd29} : s = 326;
	{8'd87,8'd30} : s = 436;
	{8'd87,8'd31} : s = 434;
	{8'd87,8'd32} : s = 497;
	{8'd87,8'd33} : s = 325;
	{8'd87,8'd34} : s = 433;
	{8'd87,8'd35} : s = 428;
	{8'd87,8'd36} : s = 492;
	{8'd87,8'd37} : s = 426;
	{8'd87,8'd38} : s = 490;
	{8'd87,8'd39} : s = 489;
	{8'd87,8'd40} : s = 508;
	{8'd87,8'd41} : s = 2;
	{8'd87,8'd42} : s = 48;
	{8'd87,8'd43} : s = 40;
	{8'd87,8'd44} : s = 168;
	{8'd87,8'd45} : s = 36;
	{8'd87,8'd46} : s = 164;
	{8'd87,8'd47} : s = 162;
	{8'd87,8'd48} : s = 323;
	{8'd87,8'd49} : s = 34;
	{8'd87,8'd50} : s = 161;
	{8'd87,8'd51} : s = 152;
	{8'd87,8'd52} : s = 312;
	{8'd87,8'd53} : s = 148;
	{8'd87,8'd54} : s = 308;
	{8'd87,8'd55} : s = 306;
	{8'd87,8'd56} : s = 425;
	{8'd87,8'd57} : s = 33;
	{8'd87,8'd58} : s = 146;
	{8'd87,8'd59} : s = 145;
	{8'd87,8'd60} : s = 305;
	{8'd87,8'd61} : s = 140;
	{8'd87,8'd62} : s = 300;
	{8'd87,8'd63} : s = 298;
	{8'd87,8'd64} : s = 422;
	{8'd87,8'd65} : s = 138;
	{8'd87,8'd66} : s = 297;
	{8'd87,8'd67} : s = 294;
	{8'd87,8'd68} : s = 421;
	{8'd87,8'd69} : s = 293;
	{8'd87,8'd70} : s = 419;
	{8'd87,8'd71} : s = 412;
	{8'd87,8'd72} : s = 486;
	{8'd87,8'd73} : s = 24;
	{8'd87,8'd74} : s = 137;
	{8'd87,8'd75} : s = 134;
	{8'd87,8'd76} : s = 291;
	{8'd87,8'd77} : s = 133;
	{8'd87,8'd78} : s = 284;
	{8'd87,8'd79} : s = 282;
	{8'd87,8'd80} : s = 410;
	{8'd87,8'd81} : s = 131;
	{8'd87,8'd82} : s = 281;
	{8'd87,8'd83} : s = 278;
	{8'd87,8'd84} : s = 409;
	{8'd87,8'd85} : s = 277;
	{8'd87,8'd86} : s = 406;
	{8'd87,8'd87} : s = 405;
	{8'd87,8'd88} : s = 485;
	{8'd87,8'd89} : s = 112;
	{8'd87,8'd90} : s = 275;
	{8'd87,8'd91} : s = 270;
	{8'd87,8'd92} : s = 403;
	{8'd87,8'd93} : s = 269;
	{8'd87,8'd94} : s = 398;
	{8'd87,8'd95} : s = 397;
	{8'd87,8'd96} : s = 483;
	{8'd87,8'd97} : s = 267;
	{8'd87,8'd98} : s = 395;
	{8'd87,8'd99} : s = 391;
	{8'd87,8'd100} : s = 476;
	{8'd87,8'd101} : s = 376;
	{8'd87,8'd102} : s = 474;
	{8'd87,8'd103} : s = 473;
	{8'd87,8'd104} : s = 506;
	{8'd87,8'd105} : s = 20;
	{8'd87,8'd106} : s = 104;
	{8'd87,8'd107} : s = 100;
	{8'd87,8'd108} : s = 263;
	{8'd87,8'd109} : s = 98;
	{8'd87,8'd110} : s = 240;
	{8'd87,8'd111} : s = 232;
	{8'd87,8'd112} : s = 372;
	{8'd87,8'd113} : s = 97;
	{8'd87,8'd114} : s = 228;
	{8'd87,8'd115} : s = 226;
	{8'd87,8'd116} : s = 370;
	{8'd87,8'd117} : s = 225;
	{8'd87,8'd118} : s = 369;
	{8'd87,8'd119} : s = 364;
	{8'd87,8'd120} : s = 470;
	{8'd87,8'd121} : s = 88;
	{8'd87,8'd122} : s = 216;
	{8'd87,8'd123} : s = 212;
	{8'd87,8'd124} : s = 362;
	{8'd87,8'd125} : s = 210;
	{8'd87,8'd126} : s = 361;
	{8'd87,8'd127} : s = 358;
	{8'd87,8'd128} : s = 469;
	{8'd87,8'd129} : s = 209;
	{8'd87,8'd130} : s = 357;
	{8'd87,8'd131} : s = 355;
	{8'd87,8'd132} : s = 467;
	{8'd87,8'd133} : s = 348;
	{8'd87,8'd134} : s = 462;
	{8'd87,8'd135} : s = 461;
	{8'd87,8'd136} : s = 505;
	{8'd87,8'd137} : s = 84;
	{8'd87,8'd138} : s = 204;
	{8'd87,8'd139} : s = 202;
	{8'd87,8'd140} : s = 346;
	{8'd87,8'd141} : s = 201;
	{8'd87,8'd142} : s = 345;
	{8'd87,8'd143} : s = 342;
	{8'd87,8'd144} : s = 459;
	{8'd87,8'd145} : s = 198;
	{8'd87,8'd146} : s = 341;
	{8'd87,8'd147} : s = 339;
	{8'd87,8'd148} : s = 455;
	{8'd87,8'd149} : s = 334;
	{8'd87,8'd150} : s = 444;
	{8'd87,8'd151} : s = 442;
	{8'd87,8'd152} : s = 502;
	{8'd87,8'd153} : s = 197;
	{8'd87,8'd154} : s = 333;
	{8'd87,8'd155} : s = 331;
	{8'd87,8'd156} : s = 441;
	{8'd87,8'd157} : s = 327;
	{8'd87,8'd158} : s = 438;
	{8'd87,8'd159} : s = 437;
	{8'd87,8'd160} : s = 501;
	{8'd87,8'd161} : s = 316;
	{8'd87,8'd162} : s = 435;
	{8'd87,8'd163} : s = 430;
	{8'd87,8'd164} : s = 499;
	{8'd87,8'd165} : s = 429;
	{8'd87,8'd166} : s = 494;
	{8'd87,8'd167} : s = 493;
	{8'd87,8'd168} : s = 510;
	{8'd87,8'd169} : s = 1;
	{8'd87,8'd170} : s = 18;
	{8'd87,8'd171} : s = 17;
	{8'd87,8'd172} : s = 82;
	{8'd87,8'd173} : s = 12;
	{8'd87,8'd174} : s = 81;
	{8'd87,8'd175} : s = 76;
	{8'd87,8'd176} : s = 195;
	{8'd87,8'd177} : s = 10;
	{8'd87,8'd178} : s = 74;
	{8'd87,8'd179} : s = 73;
	{8'd87,8'd180} : s = 184;
	{8'd87,8'd181} : s = 70;
	{8'd87,8'd182} : s = 180;
	{8'd87,8'd183} : s = 178;
	{8'd87,8'd184} : s = 314;
	{8'd87,8'd185} : s = 9;
	{8'd87,8'd186} : s = 69;
	{8'd87,8'd187} : s = 67;
	{8'd87,8'd188} : s = 177;
	{8'd87,8'd189} : s = 56;
	{8'd87,8'd190} : s = 172;
	{8'd87,8'd191} : s = 170;
	{8'd87,8'd192} : s = 313;
	{8'd87,8'd193} : s = 52;
	{8'd87,8'd194} : s = 169;
	{8'd87,8'd195} : s = 166;
	{8'd87,8'd196} : s = 310;
	{8'd87,8'd197} : s = 165;
	{8'd87,8'd198} : s = 309;
	{8'd87,8'd199} : s = 307;
	{8'd87,8'd200} : s = 427;
	{8'd87,8'd201} : s = 6;
	{8'd87,8'd202} : s = 50;
	{8'd87,8'd203} : s = 49;
	{8'd87,8'd204} : s = 163;
	{8'd87,8'd205} : s = 44;
	{8'd87,8'd206} : s = 156;
	{8'd87,8'd207} : s = 154;
	{8'd87,8'd208} : s = 302;
	{8'd87,8'd209} : s = 42;
	{8'd87,8'd210} : s = 153;
	{8'd87,8'd211} : s = 150;
	{8'd87,8'd212} : s = 301;
	{8'd87,8'd213} : s = 149;
	{8'd87,8'd214} : s = 299;
	{8'd87,8'd215} : s = 295;
	{8'd87,8'd216} : s = 423;
	{8'd87,8'd217} : s = 41;
	{8'd87,8'd218} : s = 147;
	{8'd87,8'd219} : s = 142;
	{8'd87,8'd220} : s = 286;
	{8'd87,8'd221} : s = 141;
	{8'd87,8'd222} : s = 285;
	{8'd87,8'd223} : s = 283;
	{8'd87,8'd224} : s = 414;
	{8'd87,8'd225} : s = 139;
	{8'd87,8'd226} : s = 279;
	{8'd87,8'd227} : s = 271;
	{8'd87,8'd228} : s = 413;
	{8'd87,8'd229} : s = 248;
	{8'd87,8'd230} : s = 411;
	{8'd87,8'd231} : s = 407;
	{8'd87,8'd232} : s = 491;
	{8'd87,8'd233} : s = 5;
	{8'd87,8'd234} : s = 38;
	{8'd87,8'd235} : s = 37;
	{8'd87,8'd236} : s = 135;
	{8'd87,8'd237} : s = 35;
	{8'd87,8'd238} : s = 120;
	{8'd87,8'd239} : s = 116;
	{8'd87,8'd240} : s = 244;
	{8'd87,8'd241} : s = 28;
	{8'd87,8'd242} : s = 114;
	{8'd87,8'd243} : s = 113;
	{8'd87,8'd244} : s = 242;
	{8'd87,8'd245} : s = 108;
	{8'd87,8'd246} : s = 241;
	{8'd87,8'd247} : s = 236;
	{8'd87,8'd248} : s = 399;
	{8'd87,8'd249} : s = 26;
	{8'd87,8'd250} : s = 106;
	{8'd87,8'd251} : s = 105;
	{8'd87,8'd252} : s = 234;
	{8'd87,8'd253} : s = 102;
	{8'd87,8'd254} : s = 233;
	{8'd87,8'd255} : s = 230;
	{8'd88,8'd0} : s = 208;
	{8'd88,8'd1} : s = 360;
	{8'd88,8'd2} : s = 356;
	{8'd88,8'd3} : s = 465;
	{8'd88,8'd4} : s = 354;
	{8'd88,8'd5} : s = 460;
	{8'd88,8'd6} : s = 458;
	{8'd88,8'd7} : s = 500;
	{8'd88,8'd8} : s = 65;
	{8'd88,8'd9} : s = 200;
	{8'd88,8'd10} : s = 196;
	{8'd88,8'd11} : s = 353;
	{8'd88,8'd12} : s = 194;
	{8'd88,8'd13} : s = 344;
	{8'd88,8'd14} : s = 340;
	{8'd88,8'd15} : s = 457;
	{8'd88,8'd16} : s = 193;
	{8'd88,8'd17} : s = 338;
	{8'd88,8'd18} : s = 337;
	{8'd88,8'd19} : s = 454;
	{8'd88,8'd20} : s = 332;
	{8'd88,8'd21} : s = 453;
	{8'd88,8'd22} : s = 451;
	{8'd88,8'd23} : s = 498;
	{8'd88,8'd24} : s = 176;
	{8'd88,8'd25} : s = 330;
	{8'd88,8'd26} : s = 329;
	{8'd88,8'd27} : s = 440;
	{8'd88,8'd28} : s = 326;
	{8'd88,8'd29} : s = 436;
	{8'd88,8'd30} : s = 434;
	{8'd88,8'd31} : s = 497;
	{8'd88,8'd32} : s = 325;
	{8'd88,8'd33} : s = 433;
	{8'd88,8'd34} : s = 428;
	{8'd88,8'd35} : s = 492;
	{8'd88,8'd36} : s = 426;
	{8'd88,8'd37} : s = 490;
	{8'd88,8'd38} : s = 489;
	{8'd88,8'd39} : s = 508;
	{8'd88,8'd40} : s = 2;
	{8'd88,8'd41} : s = 48;
	{8'd88,8'd42} : s = 40;
	{8'd88,8'd43} : s = 168;
	{8'd88,8'd44} : s = 36;
	{8'd88,8'd45} : s = 164;
	{8'd88,8'd46} : s = 162;
	{8'd88,8'd47} : s = 323;
	{8'd88,8'd48} : s = 34;
	{8'd88,8'd49} : s = 161;
	{8'd88,8'd50} : s = 152;
	{8'd88,8'd51} : s = 312;
	{8'd88,8'd52} : s = 148;
	{8'd88,8'd53} : s = 308;
	{8'd88,8'd54} : s = 306;
	{8'd88,8'd55} : s = 425;
	{8'd88,8'd56} : s = 33;
	{8'd88,8'd57} : s = 146;
	{8'd88,8'd58} : s = 145;
	{8'd88,8'd59} : s = 305;
	{8'd88,8'd60} : s = 140;
	{8'd88,8'd61} : s = 300;
	{8'd88,8'd62} : s = 298;
	{8'd88,8'd63} : s = 422;
	{8'd88,8'd64} : s = 138;
	{8'd88,8'd65} : s = 297;
	{8'd88,8'd66} : s = 294;
	{8'd88,8'd67} : s = 421;
	{8'd88,8'd68} : s = 293;
	{8'd88,8'd69} : s = 419;
	{8'd88,8'd70} : s = 412;
	{8'd88,8'd71} : s = 486;
	{8'd88,8'd72} : s = 24;
	{8'd88,8'd73} : s = 137;
	{8'd88,8'd74} : s = 134;
	{8'd88,8'd75} : s = 291;
	{8'd88,8'd76} : s = 133;
	{8'd88,8'd77} : s = 284;
	{8'd88,8'd78} : s = 282;
	{8'd88,8'd79} : s = 410;
	{8'd88,8'd80} : s = 131;
	{8'd88,8'd81} : s = 281;
	{8'd88,8'd82} : s = 278;
	{8'd88,8'd83} : s = 409;
	{8'd88,8'd84} : s = 277;
	{8'd88,8'd85} : s = 406;
	{8'd88,8'd86} : s = 405;
	{8'd88,8'd87} : s = 485;
	{8'd88,8'd88} : s = 112;
	{8'd88,8'd89} : s = 275;
	{8'd88,8'd90} : s = 270;
	{8'd88,8'd91} : s = 403;
	{8'd88,8'd92} : s = 269;
	{8'd88,8'd93} : s = 398;
	{8'd88,8'd94} : s = 397;
	{8'd88,8'd95} : s = 483;
	{8'd88,8'd96} : s = 267;
	{8'd88,8'd97} : s = 395;
	{8'd88,8'd98} : s = 391;
	{8'd88,8'd99} : s = 476;
	{8'd88,8'd100} : s = 376;
	{8'd88,8'd101} : s = 474;
	{8'd88,8'd102} : s = 473;
	{8'd88,8'd103} : s = 506;
	{8'd88,8'd104} : s = 20;
	{8'd88,8'd105} : s = 104;
	{8'd88,8'd106} : s = 100;
	{8'd88,8'd107} : s = 263;
	{8'd88,8'd108} : s = 98;
	{8'd88,8'd109} : s = 240;
	{8'd88,8'd110} : s = 232;
	{8'd88,8'd111} : s = 372;
	{8'd88,8'd112} : s = 97;
	{8'd88,8'd113} : s = 228;
	{8'd88,8'd114} : s = 226;
	{8'd88,8'd115} : s = 370;
	{8'd88,8'd116} : s = 225;
	{8'd88,8'd117} : s = 369;
	{8'd88,8'd118} : s = 364;
	{8'd88,8'd119} : s = 470;
	{8'd88,8'd120} : s = 88;
	{8'd88,8'd121} : s = 216;
	{8'd88,8'd122} : s = 212;
	{8'd88,8'd123} : s = 362;
	{8'd88,8'd124} : s = 210;
	{8'd88,8'd125} : s = 361;
	{8'd88,8'd126} : s = 358;
	{8'd88,8'd127} : s = 469;
	{8'd88,8'd128} : s = 209;
	{8'd88,8'd129} : s = 357;
	{8'd88,8'd130} : s = 355;
	{8'd88,8'd131} : s = 467;
	{8'd88,8'd132} : s = 348;
	{8'd88,8'd133} : s = 462;
	{8'd88,8'd134} : s = 461;
	{8'd88,8'd135} : s = 505;
	{8'd88,8'd136} : s = 84;
	{8'd88,8'd137} : s = 204;
	{8'd88,8'd138} : s = 202;
	{8'd88,8'd139} : s = 346;
	{8'd88,8'd140} : s = 201;
	{8'd88,8'd141} : s = 345;
	{8'd88,8'd142} : s = 342;
	{8'd88,8'd143} : s = 459;
	{8'd88,8'd144} : s = 198;
	{8'd88,8'd145} : s = 341;
	{8'd88,8'd146} : s = 339;
	{8'd88,8'd147} : s = 455;
	{8'd88,8'd148} : s = 334;
	{8'd88,8'd149} : s = 444;
	{8'd88,8'd150} : s = 442;
	{8'd88,8'd151} : s = 502;
	{8'd88,8'd152} : s = 197;
	{8'd88,8'd153} : s = 333;
	{8'd88,8'd154} : s = 331;
	{8'd88,8'd155} : s = 441;
	{8'd88,8'd156} : s = 327;
	{8'd88,8'd157} : s = 438;
	{8'd88,8'd158} : s = 437;
	{8'd88,8'd159} : s = 501;
	{8'd88,8'd160} : s = 316;
	{8'd88,8'd161} : s = 435;
	{8'd88,8'd162} : s = 430;
	{8'd88,8'd163} : s = 499;
	{8'd88,8'd164} : s = 429;
	{8'd88,8'd165} : s = 494;
	{8'd88,8'd166} : s = 493;
	{8'd88,8'd167} : s = 510;
	{8'd88,8'd168} : s = 1;
	{8'd88,8'd169} : s = 18;
	{8'd88,8'd170} : s = 17;
	{8'd88,8'd171} : s = 82;
	{8'd88,8'd172} : s = 12;
	{8'd88,8'd173} : s = 81;
	{8'd88,8'd174} : s = 76;
	{8'd88,8'd175} : s = 195;
	{8'd88,8'd176} : s = 10;
	{8'd88,8'd177} : s = 74;
	{8'd88,8'd178} : s = 73;
	{8'd88,8'd179} : s = 184;
	{8'd88,8'd180} : s = 70;
	{8'd88,8'd181} : s = 180;
	{8'd88,8'd182} : s = 178;
	{8'd88,8'd183} : s = 314;
	{8'd88,8'd184} : s = 9;
	{8'd88,8'd185} : s = 69;
	{8'd88,8'd186} : s = 67;
	{8'd88,8'd187} : s = 177;
	{8'd88,8'd188} : s = 56;
	{8'd88,8'd189} : s = 172;
	{8'd88,8'd190} : s = 170;
	{8'd88,8'd191} : s = 313;
	{8'd88,8'd192} : s = 52;
	{8'd88,8'd193} : s = 169;
	{8'd88,8'd194} : s = 166;
	{8'd88,8'd195} : s = 310;
	{8'd88,8'd196} : s = 165;
	{8'd88,8'd197} : s = 309;
	{8'd88,8'd198} : s = 307;
	{8'd88,8'd199} : s = 427;
	{8'd88,8'd200} : s = 6;
	{8'd88,8'd201} : s = 50;
	{8'd88,8'd202} : s = 49;
	{8'd88,8'd203} : s = 163;
	{8'd88,8'd204} : s = 44;
	{8'd88,8'd205} : s = 156;
	{8'd88,8'd206} : s = 154;
	{8'd88,8'd207} : s = 302;
	{8'd88,8'd208} : s = 42;
	{8'd88,8'd209} : s = 153;
	{8'd88,8'd210} : s = 150;
	{8'd88,8'd211} : s = 301;
	{8'd88,8'd212} : s = 149;
	{8'd88,8'd213} : s = 299;
	{8'd88,8'd214} : s = 295;
	{8'd88,8'd215} : s = 423;
	{8'd88,8'd216} : s = 41;
	{8'd88,8'd217} : s = 147;
	{8'd88,8'd218} : s = 142;
	{8'd88,8'd219} : s = 286;
	{8'd88,8'd220} : s = 141;
	{8'd88,8'd221} : s = 285;
	{8'd88,8'd222} : s = 283;
	{8'd88,8'd223} : s = 414;
	{8'd88,8'd224} : s = 139;
	{8'd88,8'd225} : s = 279;
	{8'd88,8'd226} : s = 271;
	{8'd88,8'd227} : s = 413;
	{8'd88,8'd228} : s = 248;
	{8'd88,8'd229} : s = 411;
	{8'd88,8'd230} : s = 407;
	{8'd88,8'd231} : s = 491;
	{8'd88,8'd232} : s = 5;
	{8'd88,8'd233} : s = 38;
	{8'd88,8'd234} : s = 37;
	{8'd88,8'd235} : s = 135;
	{8'd88,8'd236} : s = 35;
	{8'd88,8'd237} : s = 120;
	{8'd88,8'd238} : s = 116;
	{8'd88,8'd239} : s = 244;
	{8'd88,8'd240} : s = 28;
	{8'd88,8'd241} : s = 114;
	{8'd88,8'd242} : s = 113;
	{8'd88,8'd243} : s = 242;
	{8'd88,8'd244} : s = 108;
	{8'd88,8'd245} : s = 241;
	{8'd88,8'd246} : s = 236;
	{8'd88,8'd247} : s = 399;
	{8'd88,8'd248} : s = 26;
	{8'd88,8'd249} : s = 106;
	{8'd88,8'd250} : s = 105;
	{8'd88,8'd251} : s = 234;
	{8'd88,8'd252} : s = 102;
	{8'd88,8'd253} : s = 233;
	{8'd88,8'd254} : s = 230;
	{8'd88,8'd255} : s = 380;
	{8'd89,8'd0} : s = 360;
	{8'd89,8'd1} : s = 356;
	{8'd89,8'd2} : s = 465;
	{8'd89,8'd3} : s = 354;
	{8'd89,8'd4} : s = 460;
	{8'd89,8'd5} : s = 458;
	{8'd89,8'd6} : s = 500;
	{8'd89,8'd7} : s = 65;
	{8'd89,8'd8} : s = 200;
	{8'd89,8'd9} : s = 196;
	{8'd89,8'd10} : s = 353;
	{8'd89,8'd11} : s = 194;
	{8'd89,8'd12} : s = 344;
	{8'd89,8'd13} : s = 340;
	{8'd89,8'd14} : s = 457;
	{8'd89,8'd15} : s = 193;
	{8'd89,8'd16} : s = 338;
	{8'd89,8'd17} : s = 337;
	{8'd89,8'd18} : s = 454;
	{8'd89,8'd19} : s = 332;
	{8'd89,8'd20} : s = 453;
	{8'd89,8'd21} : s = 451;
	{8'd89,8'd22} : s = 498;
	{8'd89,8'd23} : s = 176;
	{8'd89,8'd24} : s = 330;
	{8'd89,8'd25} : s = 329;
	{8'd89,8'd26} : s = 440;
	{8'd89,8'd27} : s = 326;
	{8'd89,8'd28} : s = 436;
	{8'd89,8'd29} : s = 434;
	{8'd89,8'd30} : s = 497;
	{8'd89,8'd31} : s = 325;
	{8'd89,8'd32} : s = 433;
	{8'd89,8'd33} : s = 428;
	{8'd89,8'd34} : s = 492;
	{8'd89,8'd35} : s = 426;
	{8'd89,8'd36} : s = 490;
	{8'd89,8'd37} : s = 489;
	{8'd89,8'd38} : s = 508;
	{8'd89,8'd39} : s = 2;
	{8'd89,8'd40} : s = 48;
	{8'd89,8'd41} : s = 40;
	{8'd89,8'd42} : s = 168;
	{8'd89,8'd43} : s = 36;
	{8'd89,8'd44} : s = 164;
	{8'd89,8'd45} : s = 162;
	{8'd89,8'd46} : s = 323;
	{8'd89,8'd47} : s = 34;
	{8'd89,8'd48} : s = 161;
	{8'd89,8'd49} : s = 152;
	{8'd89,8'd50} : s = 312;
	{8'd89,8'd51} : s = 148;
	{8'd89,8'd52} : s = 308;
	{8'd89,8'd53} : s = 306;
	{8'd89,8'd54} : s = 425;
	{8'd89,8'd55} : s = 33;
	{8'd89,8'd56} : s = 146;
	{8'd89,8'd57} : s = 145;
	{8'd89,8'd58} : s = 305;
	{8'd89,8'd59} : s = 140;
	{8'd89,8'd60} : s = 300;
	{8'd89,8'd61} : s = 298;
	{8'd89,8'd62} : s = 422;
	{8'd89,8'd63} : s = 138;
	{8'd89,8'd64} : s = 297;
	{8'd89,8'd65} : s = 294;
	{8'd89,8'd66} : s = 421;
	{8'd89,8'd67} : s = 293;
	{8'd89,8'd68} : s = 419;
	{8'd89,8'd69} : s = 412;
	{8'd89,8'd70} : s = 486;
	{8'd89,8'd71} : s = 24;
	{8'd89,8'd72} : s = 137;
	{8'd89,8'd73} : s = 134;
	{8'd89,8'd74} : s = 291;
	{8'd89,8'd75} : s = 133;
	{8'd89,8'd76} : s = 284;
	{8'd89,8'd77} : s = 282;
	{8'd89,8'd78} : s = 410;
	{8'd89,8'd79} : s = 131;
	{8'd89,8'd80} : s = 281;
	{8'd89,8'd81} : s = 278;
	{8'd89,8'd82} : s = 409;
	{8'd89,8'd83} : s = 277;
	{8'd89,8'd84} : s = 406;
	{8'd89,8'd85} : s = 405;
	{8'd89,8'd86} : s = 485;
	{8'd89,8'd87} : s = 112;
	{8'd89,8'd88} : s = 275;
	{8'd89,8'd89} : s = 270;
	{8'd89,8'd90} : s = 403;
	{8'd89,8'd91} : s = 269;
	{8'd89,8'd92} : s = 398;
	{8'd89,8'd93} : s = 397;
	{8'd89,8'd94} : s = 483;
	{8'd89,8'd95} : s = 267;
	{8'd89,8'd96} : s = 395;
	{8'd89,8'd97} : s = 391;
	{8'd89,8'd98} : s = 476;
	{8'd89,8'd99} : s = 376;
	{8'd89,8'd100} : s = 474;
	{8'd89,8'd101} : s = 473;
	{8'd89,8'd102} : s = 506;
	{8'd89,8'd103} : s = 20;
	{8'd89,8'd104} : s = 104;
	{8'd89,8'd105} : s = 100;
	{8'd89,8'd106} : s = 263;
	{8'd89,8'd107} : s = 98;
	{8'd89,8'd108} : s = 240;
	{8'd89,8'd109} : s = 232;
	{8'd89,8'd110} : s = 372;
	{8'd89,8'd111} : s = 97;
	{8'd89,8'd112} : s = 228;
	{8'd89,8'd113} : s = 226;
	{8'd89,8'd114} : s = 370;
	{8'd89,8'd115} : s = 225;
	{8'd89,8'd116} : s = 369;
	{8'd89,8'd117} : s = 364;
	{8'd89,8'd118} : s = 470;
	{8'd89,8'd119} : s = 88;
	{8'd89,8'd120} : s = 216;
	{8'd89,8'd121} : s = 212;
	{8'd89,8'd122} : s = 362;
	{8'd89,8'd123} : s = 210;
	{8'd89,8'd124} : s = 361;
	{8'd89,8'd125} : s = 358;
	{8'd89,8'd126} : s = 469;
	{8'd89,8'd127} : s = 209;
	{8'd89,8'd128} : s = 357;
	{8'd89,8'd129} : s = 355;
	{8'd89,8'd130} : s = 467;
	{8'd89,8'd131} : s = 348;
	{8'd89,8'd132} : s = 462;
	{8'd89,8'd133} : s = 461;
	{8'd89,8'd134} : s = 505;
	{8'd89,8'd135} : s = 84;
	{8'd89,8'd136} : s = 204;
	{8'd89,8'd137} : s = 202;
	{8'd89,8'd138} : s = 346;
	{8'd89,8'd139} : s = 201;
	{8'd89,8'd140} : s = 345;
	{8'd89,8'd141} : s = 342;
	{8'd89,8'd142} : s = 459;
	{8'd89,8'd143} : s = 198;
	{8'd89,8'd144} : s = 341;
	{8'd89,8'd145} : s = 339;
	{8'd89,8'd146} : s = 455;
	{8'd89,8'd147} : s = 334;
	{8'd89,8'd148} : s = 444;
	{8'd89,8'd149} : s = 442;
	{8'd89,8'd150} : s = 502;
	{8'd89,8'd151} : s = 197;
	{8'd89,8'd152} : s = 333;
	{8'd89,8'd153} : s = 331;
	{8'd89,8'd154} : s = 441;
	{8'd89,8'd155} : s = 327;
	{8'd89,8'd156} : s = 438;
	{8'd89,8'd157} : s = 437;
	{8'd89,8'd158} : s = 501;
	{8'd89,8'd159} : s = 316;
	{8'd89,8'd160} : s = 435;
	{8'd89,8'd161} : s = 430;
	{8'd89,8'd162} : s = 499;
	{8'd89,8'd163} : s = 429;
	{8'd89,8'd164} : s = 494;
	{8'd89,8'd165} : s = 493;
	{8'd89,8'd166} : s = 510;
	{8'd89,8'd167} : s = 1;
	{8'd89,8'd168} : s = 18;
	{8'd89,8'd169} : s = 17;
	{8'd89,8'd170} : s = 82;
	{8'd89,8'd171} : s = 12;
	{8'd89,8'd172} : s = 81;
	{8'd89,8'd173} : s = 76;
	{8'd89,8'd174} : s = 195;
	{8'd89,8'd175} : s = 10;
	{8'd89,8'd176} : s = 74;
	{8'd89,8'd177} : s = 73;
	{8'd89,8'd178} : s = 184;
	{8'd89,8'd179} : s = 70;
	{8'd89,8'd180} : s = 180;
	{8'd89,8'd181} : s = 178;
	{8'd89,8'd182} : s = 314;
	{8'd89,8'd183} : s = 9;
	{8'd89,8'd184} : s = 69;
	{8'd89,8'd185} : s = 67;
	{8'd89,8'd186} : s = 177;
	{8'd89,8'd187} : s = 56;
	{8'd89,8'd188} : s = 172;
	{8'd89,8'd189} : s = 170;
	{8'd89,8'd190} : s = 313;
	{8'd89,8'd191} : s = 52;
	{8'd89,8'd192} : s = 169;
	{8'd89,8'd193} : s = 166;
	{8'd89,8'd194} : s = 310;
	{8'd89,8'd195} : s = 165;
	{8'd89,8'd196} : s = 309;
	{8'd89,8'd197} : s = 307;
	{8'd89,8'd198} : s = 427;
	{8'd89,8'd199} : s = 6;
	{8'd89,8'd200} : s = 50;
	{8'd89,8'd201} : s = 49;
	{8'd89,8'd202} : s = 163;
	{8'd89,8'd203} : s = 44;
	{8'd89,8'd204} : s = 156;
	{8'd89,8'd205} : s = 154;
	{8'd89,8'd206} : s = 302;
	{8'd89,8'd207} : s = 42;
	{8'd89,8'd208} : s = 153;
	{8'd89,8'd209} : s = 150;
	{8'd89,8'd210} : s = 301;
	{8'd89,8'd211} : s = 149;
	{8'd89,8'd212} : s = 299;
	{8'd89,8'd213} : s = 295;
	{8'd89,8'd214} : s = 423;
	{8'd89,8'd215} : s = 41;
	{8'd89,8'd216} : s = 147;
	{8'd89,8'd217} : s = 142;
	{8'd89,8'd218} : s = 286;
	{8'd89,8'd219} : s = 141;
	{8'd89,8'd220} : s = 285;
	{8'd89,8'd221} : s = 283;
	{8'd89,8'd222} : s = 414;
	{8'd89,8'd223} : s = 139;
	{8'd89,8'd224} : s = 279;
	{8'd89,8'd225} : s = 271;
	{8'd89,8'd226} : s = 413;
	{8'd89,8'd227} : s = 248;
	{8'd89,8'd228} : s = 411;
	{8'd89,8'd229} : s = 407;
	{8'd89,8'd230} : s = 491;
	{8'd89,8'd231} : s = 5;
	{8'd89,8'd232} : s = 38;
	{8'd89,8'd233} : s = 37;
	{8'd89,8'd234} : s = 135;
	{8'd89,8'd235} : s = 35;
	{8'd89,8'd236} : s = 120;
	{8'd89,8'd237} : s = 116;
	{8'd89,8'd238} : s = 244;
	{8'd89,8'd239} : s = 28;
	{8'd89,8'd240} : s = 114;
	{8'd89,8'd241} : s = 113;
	{8'd89,8'd242} : s = 242;
	{8'd89,8'd243} : s = 108;
	{8'd89,8'd244} : s = 241;
	{8'd89,8'd245} : s = 236;
	{8'd89,8'd246} : s = 399;
	{8'd89,8'd247} : s = 26;
	{8'd89,8'd248} : s = 106;
	{8'd89,8'd249} : s = 105;
	{8'd89,8'd250} : s = 234;
	{8'd89,8'd251} : s = 102;
	{8'd89,8'd252} : s = 233;
	{8'd89,8'd253} : s = 230;
	{8'd89,8'd254} : s = 380;
	{8'd89,8'd255} : s = 101;
	{8'd90,8'd0} : s = 356;
	{8'd90,8'd1} : s = 465;
	{8'd90,8'd2} : s = 354;
	{8'd90,8'd3} : s = 460;
	{8'd90,8'd4} : s = 458;
	{8'd90,8'd5} : s = 500;
	{8'd90,8'd6} : s = 65;
	{8'd90,8'd7} : s = 200;
	{8'd90,8'd8} : s = 196;
	{8'd90,8'd9} : s = 353;
	{8'd90,8'd10} : s = 194;
	{8'd90,8'd11} : s = 344;
	{8'd90,8'd12} : s = 340;
	{8'd90,8'd13} : s = 457;
	{8'd90,8'd14} : s = 193;
	{8'd90,8'd15} : s = 338;
	{8'd90,8'd16} : s = 337;
	{8'd90,8'd17} : s = 454;
	{8'd90,8'd18} : s = 332;
	{8'd90,8'd19} : s = 453;
	{8'd90,8'd20} : s = 451;
	{8'd90,8'd21} : s = 498;
	{8'd90,8'd22} : s = 176;
	{8'd90,8'd23} : s = 330;
	{8'd90,8'd24} : s = 329;
	{8'd90,8'd25} : s = 440;
	{8'd90,8'd26} : s = 326;
	{8'd90,8'd27} : s = 436;
	{8'd90,8'd28} : s = 434;
	{8'd90,8'd29} : s = 497;
	{8'd90,8'd30} : s = 325;
	{8'd90,8'd31} : s = 433;
	{8'd90,8'd32} : s = 428;
	{8'd90,8'd33} : s = 492;
	{8'd90,8'd34} : s = 426;
	{8'd90,8'd35} : s = 490;
	{8'd90,8'd36} : s = 489;
	{8'd90,8'd37} : s = 508;
	{8'd90,8'd38} : s = 2;
	{8'd90,8'd39} : s = 48;
	{8'd90,8'd40} : s = 40;
	{8'd90,8'd41} : s = 168;
	{8'd90,8'd42} : s = 36;
	{8'd90,8'd43} : s = 164;
	{8'd90,8'd44} : s = 162;
	{8'd90,8'd45} : s = 323;
	{8'd90,8'd46} : s = 34;
	{8'd90,8'd47} : s = 161;
	{8'd90,8'd48} : s = 152;
	{8'd90,8'd49} : s = 312;
	{8'd90,8'd50} : s = 148;
	{8'd90,8'd51} : s = 308;
	{8'd90,8'd52} : s = 306;
	{8'd90,8'd53} : s = 425;
	{8'd90,8'd54} : s = 33;
	{8'd90,8'd55} : s = 146;
	{8'd90,8'd56} : s = 145;
	{8'd90,8'd57} : s = 305;
	{8'd90,8'd58} : s = 140;
	{8'd90,8'd59} : s = 300;
	{8'd90,8'd60} : s = 298;
	{8'd90,8'd61} : s = 422;
	{8'd90,8'd62} : s = 138;
	{8'd90,8'd63} : s = 297;
	{8'd90,8'd64} : s = 294;
	{8'd90,8'd65} : s = 421;
	{8'd90,8'd66} : s = 293;
	{8'd90,8'd67} : s = 419;
	{8'd90,8'd68} : s = 412;
	{8'd90,8'd69} : s = 486;
	{8'd90,8'd70} : s = 24;
	{8'd90,8'd71} : s = 137;
	{8'd90,8'd72} : s = 134;
	{8'd90,8'd73} : s = 291;
	{8'd90,8'd74} : s = 133;
	{8'd90,8'd75} : s = 284;
	{8'd90,8'd76} : s = 282;
	{8'd90,8'd77} : s = 410;
	{8'd90,8'd78} : s = 131;
	{8'd90,8'd79} : s = 281;
	{8'd90,8'd80} : s = 278;
	{8'd90,8'd81} : s = 409;
	{8'd90,8'd82} : s = 277;
	{8'd90,8'd83} : s = 406;
	{8'd90,8'd84} : s = 405;
	{8'd90,8'd85} : s = 485;
	{8'd90,8'd86} : s = 112;
	{8'd90,8'd87} : s = 275;
	{8'd90,8'd88} : s = 270;
	{8'd90,8'd89} : s = 403;
	{8'd90,8'd90} : s = 269;
	{8'd90,8'd91} : s = 398;
	{8'd90,8'd92} : s = 397;
	{8'd90,8'd93} : s = 483;
	{8'd90,8'd94} : s = 267;
	{8'd90,8'd95} : s = 395;
	{8'd90,8'd96} : s = 391;
	{8'd90,8'd97} : s = 476;
	{8'd90,8'd98} : s = 376;
	{8'd90,8'd99} : s = 474;
	{8'd90,8'd100} : s = 473;
	{8'd90,8'd101} : s = 506;
	{8'd90,8'd102} : s = 20;
	{8'd90,8'd103} : s = 104;
	{8'd90,8'd104} : s = 100;
	{8'd90,8'd105} : s = 263;
	{8'd90,8'd106} : s = 98;
	{8'd90,8'd107} : s = 240;
	{8'd90,8'd108} : s = 232;
	{8'd90,8'd109} : s = 372;
	{8'd90,8'd110} : s = 97;
	{8'd90,8'd111} : s = 228;
	{8'd90,8'd112} : s = 226;
	{8'd90,8'd113} : s = 370;
	{8'd90,8'd114} : s = 225;
	{8'd90,8'd115} : s = 369;
	{8'd90,8'd116} : s = 364;
	{8'd90,8'd117} : s = 470;
	{8'd90,8'd118} : s = 88;
	{8'd90,8'd119} : s = 216;
	{8'd90,8'd120} : s = 212;
	{8'd90,8'd121} : s = 362;
	{8'd90,8'd122} : s = 210;
	{8'd90,8'd123} : s = 361;
	{8'd90,8'd124} : s = 358;
	{8'd90,8'd125} : s = 469;
	{8'd90,8'd126} : s = 209;
	{8'd90,8'd127} : s = 357;
	{8'd90,8'd128} : s = 355;
	{8'd90,8'd129} : s = 467;
	{8'd90,8'd130} : s = 348;
	{8'd90,8'd131} : s = 462;
	{8'd90,8'd132} : s = 461;
	{8'd90,8'd133} : s = 505;
	{8'd90,8'd134} : s = 84;
	{8'd90,8'd135} : s = 204;
	{8'd90,8'd136} : s = 202;
	{8'd90,8'd137} : s = 346;
	{8'd90,8'd138} : s = 201;
	{8'd90,8'd139} : s = 345;
	{8'd90,8'd140} : s = 342;
	{8'd90,8'd141} : s = 459;
	{8'd90,8'd142} : s = 198;
	{8'd90,8'd143} : s = 341;
	{8'd90,8'd144} : s = 339;
	{8'd90,8'd145} : s = 455;
	{8'd90,8'd146} : s = 334;
	{8'd90,8'd147} : s = 444;
	{8'd90,8'd148} : s = 442;
	{8'd90,8'd149} : s = 502;
	{8'd90,8'd150} : s = 197;
	{8'd90,8'd151} : s = 333;
	{8'd90,8'd152} : s = 331;
	{8'd90,8'd153} : s = 441;
	{8'd90,8'd154} : s = 327;
	{8'd90,8'd155} : s = 438;
	{8'd90,8'd156} : s = 437;
	{8'd90,8'd157} : s = 501;
	{8'd90,8'd158} : s = 316;
	{8'd90,8'd159} : s = 435;
	{8'd90,8'd160} : s = 430;
	{8'd90,8'd161} : s = 499;
	{8'd90,8'd162} : s = 429;
	{8'd90,8'd163} : s = 494;
	{8'd90,8'd164} : s = 493;
	{8'd90,8'd165} : s = 510;
	{8'd90,8'd166} : s = 1;
	{8'd90,8'd167} : s = 18;
	{8'd90,8'd168} : s = 17;
	{8'd90,8'd169} : s = 82;
	{8'd90,8'd170} : s = 12;
	{8'd90,8'd171} : s = 81;
	{8'd90,8'd172} : s = 76;
	{8'd90,8'd173} : s = 195;
	{8'd90,8'd174} : s = 10;
	{8'd90,8'd175} : s = 74;
	{8'd90,8'd176} : s = 73;
	{8'd90,8'd177} : s = 184;
	{8'd90,8'd178} : s = 70;
	{8'd90,8'd179} : s = 180;
	{8'd90,8'd180} : s = 178;
	{8'd90,8'd181} : s = 314;
	{8'd90,8'd182} : s = 9;
	{8'd90,8'd183} : s = 69;
	{8'd90,8'd184} : s = 67;
	{8'd90,8'd185} : s = 177;
	{8'd90,8'd186} : s = 56;
	{8'd90,8'd187} : s = 172;
	{8'd90,8'd188} : s = 170;
	{8'd90,8'd189} : s = 313;
	{8'd90,8'd190} : s = 52;
	{8'd90,8'd191} : s = 169;
	{8'd90,8'd192} : s = 166;
	{8'd90,8'd193} : s = 310;
	{8'd90,8'd194} : s = 165;
	{8'd90,8'd195} : s = 309;
	{8'd90,8'd196} : s = 307;
	{8'd90,8'd197} : s = 427;
	{8'd90,8'd198} : s = 6;
	{8'd90,8'd199} : s = 50;
	{8'd90,8'd200} : s = 49;
	{8'd90,8'd201} : s = 163;
	{8'd90,8'd202} : s = 44;
	{8'd90,8'd203} : s = 156;
	{8'd90,8'd204} : s = 154;
	{8'd90,8'd205} : s = 302;
	{8'd90,8'd206} : s = 42;
	{8'd90,8'd207} : s = 153;
	{8'd90,8'd208} : s = 150;
	{8'd90,8'd209} : s = 301;
	{8'd90,8'd210} : s = 149;
	{8'd90,8'd211} : s = 299;
	{8'd90,8'd212} : s = 295;
	{8'd90,8'd213} : s = 423;
	{8'd90,8'd214} : s = 41;
	{8'd90,8'd215} : s = 147;
	{8'd90,8'd216} : s = 142;
	{8'd90,8'd217} : s = 286;
	{8'd90,8'd218} : s = 141;
	{8'd90,8'd219} : s = 285;
	{8'd90,8'd220} : s = 283;
	{8'd90,8'd221} : s = 414;
	{8'd90,8'd222} : s = 139;
	{8'd90,8'd223} : s = 279;
	{8'd90,8'd224} : s = 271;
	{8'd90,8'd225} : s = 413;
	{8'd90,8'd226} : s = 248;
	{8'd90,8'd227} : s = 411;
	{8'd90,8'd228} : s = 407;
	{8'd90,8'd229} : s = 491;
	{8'd90,8'd230} : s = 5;
	{8'd90,8'd231} : s = 38;
	{8'd90,8'd232} : s = 37;
	{8'd90,8'd233} : s = 135;
	{8'd90,8'd234} : s = 35;
	{8'd90,8'd235} : s = 120;
	{8'd90,8'd236} : s = 116;
	{8'd90,8'd237} : s = 244;
	{8'd90,8'd238} : s = 28;
	{8'd90,8'd239} : s = 114;
	{8'd90,8'd240} : s = 113;
	{8'd90,8'd241} : s = 242;
	{8'd90,8'd242} : s = 108;
	{8'd90,8'd243} : s = 241;
	{8'd90,8'd244} : s = 236;
	{8'd90,8'd245} : s = 399;
	{8'd90,8'd246} : s = 26;
	{8'd90,8'd247} : s = 106;
	{8'd90,8'd248} : s = 105;
	{8'd90,8'd249} : s = 234;
	{8'd90,8'd250} : s = 102;
	{8'd90,8'd251} : s = 233;
	{8'd90,8'd252} : s = 230;
	{8'd90,8'd253} : s = 380;
	{8'd90,8'd254} : s = 101;
	{8'd90,8'd255} : s = 229;
	{8'd91,8'd0} : s = 465;
	{8'd91,8'd1} : s = 354;
	{8'd91,8'd2} : s = 460;
	{8'd91,8'd3} : s = 458;
	{8'd91,8'd4} : s = 500;
	{8'd91,8'd5} : s = 65;
	{8'd91,8'd6} : s = 200;
	{8'd91,8'd7} : s = 196;
	{8'd91,8'd8} : s = 353;
	{8'd91,8'd9} : s = 194;
	{8'd91,8'd10} : s = 344;
	{8'd91,8'd11} : s = 340;
	{8'd91,8'd12} : s = 457;
	{8'd91,8'd13} : s = 193;
	{8'd91,8'd14} : s = 338;
	{8'd91,8'd15} : s = 337;
	{8'd91,8'd16} : s = 454;
	{8'd91,8'd17} : s = 332;
	{8'd91,8'd18} : s = 453;
	{8'd91,8'd19} : s = 451;
	{8'd91,8'd20} : s = 498;
	{8'd91,8'd21} : s = 176;
	{8'd91,8'd22} : s = 330;
	{8'd91,8'd23} : s = 329;
	{8'd91,8'd24} : s = 440;
	{8'd91,8'd25} : s = 326;
	{8'd91,8'd26} : s = 436;
	{8'd91,8'd27} : s = 434;
	{8'd91,8'd28} : s = 497;
	{8'd91,8'd29} : s = 325;
	{8'd91,8'd30} : s = 433;
	{8'd91,8'd31} : s = 428;
	{8'd91,8'd32} : s = 492;
	{8'd91,8'd33} : s = 426;
	{8'd91,8'd34} : s = 490;
	{8'd91,8'd35} : s = 489;
	{8'd91,8'd36} : s = 508;
	{8'd91,8'd37} : s = 2;
	{8'd91,8'd38} : s = 48;
	{8'd91,8'd39} : s = 40;
	{8'd91,8'd40} : s = 168;
	{8'd91,8'd41} : s = 36;
	{8'd91,8'd42} : s = 164;
	{8'd91,8'd43} : s = 162;
	{8'd91,8'd44} : s = 323;
	{8'd91,8'd45} : s = 34;
	{8'd91,8'd46} : s = 161;
	{8'd91,8'd47} : s = 152;
	{8'd91,8'd48} : s = 312;
	{8'd91,8'd49} : s = 148;
	{8'd91,8'd50} : s = 308;
	{8'd91,8'd51} : s = 306;
	{8'd91,8'd52} : s = 425;
	{8'd91,8'd53} : s = 33;
	{8'd91,8'd54} : s = 146;
	{8'd91,8'd55} : s = 145;
	{8'd91,8'd56} : s = 305;
	{8'd91,8'd57} : s = 140;
	{8'd91,8'd58} : s = 300;
	{8'd91,8'd59} : s = 298;
	{8'd91,8'd60} : s = 422;
	{8'd91,8'd61} : s = 138;
	{8'd91,8'd62} : s = 297;
	{8'd91,8'd63} : s = 294;
	{8'd91,8'd64} : s = 421;
	{8'd91,8'd65} : s = 293;
	{8'd91,8'd66} : s = 419;
	{8'd91,8'd67} : s = 412;
	{8'd91,8'd68} : s = 486;
	{8'd91,8'd69} : s = 24;
	{8'd91,8'd70} : s = 137;
	{8'd91,8'd71} : s = 134;
	{8'd91,8'd72} : s = 291;
	{8'd91,8'd73} : s = 133;
	{8'd91,8'd74} : s = 284;
	{8'd91,8'd75} : s = 282;
	{8'd91,8'd76} : s = 410;
	{8'd91,8'd77} : s = 131;
	{8'd91,8'd78} : s = 281;
	{8'd91,8'd79} : s = 278;
	{8'd91,8'd80} : s = 409;
	{8'd91,8'd81} : s = 277;
	{8'd91,8'd82} : s = 406;
	{8'd91,8'd83} : s = 405;
	{8'd91,8'd84} : s = 485;
	{8'd91,8'd85} : s = 112;
	{8'd91,8'd86} : s = 275;
	{8'd91,8'd87} : s = 270;
	{8'd91,8'd88} : s = 403;
	{8'd91,8'd89} : s = 269;
	{8'd91,8'd90} : s = 398;
	{8'd91,8'd91} : s = 397;
	{8'd91,8'd92} : s = 483;
	{8'd91,8'd93} : s = 267;
	{8'd91,8'd94} : s = 395;
	{8'd91,8'd95} : s = 391;
	{8'd91,8'd96} : s = 476;
	{8'd91,8'd97} : s = 376;
	{8'd91,8'd98} : s = 474;
	{8'd91,8'd99} : s = 473;
	{8'd91,8'd100} : s = 506;
	{8'd91,8'd101} : s = 20;
	{8'd91,8'd102} : s = 104;
	{8'd91,8'd103} : s = 100;
	{8'd91,8'd104} : s = 263;
	{8'd91,8'd105} : s = 98;
	{8'd91,8'd106} : s = 240;
	{8'd91,8'd107} : s = 232;
	{8'd91,8'd108} : s = 372;
	{8'd91,8'd109} : s = 97;
	{8'd91,8'd110} : s = 228;
	{8'd91,8'd111} : s = 226;
	{8'd91,8'd112} : s = 370;
	{8'd91,8'd113} : s = 225;
	{8'd91,8'd114} : s = 369;
	{8'd91,8'd115} : s = 364;
	{8'd91,8'd116} : s = 470;
	{8'd91,8'd117} : s = 88;
	{8'd91,8'd118} : s = 216;
	{8'd91,8'd119} : s = 212;
	{8'd91,8'd120} : s = 362;
	{8'd91,8'd121} : s = 210;
	{8'd91,8'd122} : s = 361;
	{8'd91,8'd123} : s = 358;
	{8'd91,8'd124} : s = 469;
	{8'd91,8'd125} : s = 209;
	{8'd91,8'd126} : s = 357;
	{8'd91,8'd127} : s = 355;
	{8'd91,8'd128} : s = 467;
	{8'd91,8'd129} : s = 348;
	{8'd91,8'd130} : s = 462;
	{8'd91,8'd131} : s = 461;
	{8'd91,8'd132} : s = 505;
	{8'd91,8'd133} : s = 84;
	{8'd91,8'd134} : s = 204;
	{8'd91,8'd135} : s = 202;
	{8'd91,8'd136} : s = 346;
	{8'd91,8'd137} : s = 201;
	{8'd91,8'd138} : s = 345;
	{8'd91,8'd139} : s = 342;
	{8'd91,8'd140} : s = 459;
	{8'd91,8'd141} : s = 198;
	{8'd91,8'd142} : s = 341;
	{8'd91,8'd143} : s = 339;
	{8'd91,8'd144} : s = 455;
	{8'd91,8'd145} : s = 334;
	{8'd91,8'd146} : s = 444;
	{8'd91,8'd147} : s = 442;
	{8'd91,8'd148} : s = 502;
	{8'd91,8'd149} : s = 197;
	{8'd91,8'd150} : s = 333;
	{8'd91,8'd151} : s = 331;
	{8'd91,8'd152} : s = 441;
	{8'd91,8'd153} : s = 327;
	{8'd91,8'd154} : s = 438;
	{8'd91,8'd155} : s = 437;
	{8'd91,8'd156} : s = 501;
	{8'd91,8'd157} : s = 316;
	{8'd91,8'd158} : s = 435;
	{8'd91,8'd159} : s = 430;
	{8'd91,8'd160} : s = 499;
	{8'd91,8'd161} : s = 429;
	{8'd91,8'd162} : s = 494;
	{8'd91,8'd163} : s = 493;
	{8'd91,8'd164} : s = 510;
	{8'd91,8'd165} : s = 1;
	{8'd91,8'd166} : s = 18;
	{8'd91,8'd167} : s = 17;
	{8'd91,8'd168} : s = 82;
	{8'd91,8'd169} : s = 12;
	{8'd91,8'd170} : s = 81;
	{8'd91,8'd171} : s = 76;
	{8'd91,8'd172} : s = 195;
	{8'd91,8'd173} : s = 10;
	{8'd91,8'd174} : s = 74;
	{8'd91,8'd175} : s = 73;
	{8'd91,8'd176} : s = 184;
	{8'd91,8'd177} : s = 70;
	{8'd91,8'd178} : s = 180;
	{8'd91,8'd179} : s = 178;
	{8'd91,8'd180} : s = 314;
	{8'd91,8'd181} : s = 9;
	{8'd91,8'd182} : s = 69;
	{8'd91,8'd183} : s = 67;
	{8'd91,8'd184} : s = 177;
	{8'd91,8'd185} : s = 56;
	{8'd91,8'd186} : s = 172;
	{8'd91,8'd187} : s = 170;
	{8'd91,8'd188} : s = 313;
	{8'd91,8'd189} : s = 52;
	{8'd91,8'd190} : s = 169;
	{8'd91,8'd191} : s = 166;
	{8'd91,8'd192} : s = 310;
	{8'd91,8'd193} : s = 165;
	{8'd91,8'd194} : s = 309;
	{8'd91,8'd195} : s = 307;
	{8'd91,8'd196} : s = 427;
	{8'd91,8'd197} : s = 6;
	{8'd91,8'd198} : s = 50;
	{8'd91,8'd199} : s = 49;
	{8'd91,8'd200} : s = 163;
	{8'd91,8'd201} : s = 44;
	{8'd91,8'd202} : s = 156;
	{8'd91,8'd203} : s = 154;
	{8'd91,8'd204} : s = 302;
	{8'd91,8'd205} : s = 42;
	{8'd91,8'd206} : s = 153;
	{8'd91,8'd207} : s = 150;
	{8'd91,8'd208} : s = 301;
	{8'd91,8'd209} : s = 149;
	{8'd91,8'd210} : s = 299;
	{8'd91,8'd211} : s = 295;
	{8'd91,8'd212} : s = 423;
	{8'd91,8'd213} : s = 41;
	{8'd91,8'd214} : s = 147;
	{8'd91,8'd215} : s = 142;
	{8'd91,8'd216} : s = 286;
	{8'd91,8'd217} : s = 141;
	{8'd91,8'd218} : s = 285;
	{8'd91,8'd219} : s = 283;
	{8'd91,8'd220} : s = 414;
	{8'd91,8'd221} : s = 139;
	{8'd91,8'd222} : s = 279;
	{8'd91,8'd223} : s = 271;
	{8'd91,8'd224} : s = 413;
	{8'd91,8'd225} : s = 248;
	{8'd91,8'd226} : s = 411;
	{8'd91,8'd227} : s = 407;
	{8'd91,8'd228} : s = 491;
	{8'd91,8'd229} : s = 5;
	{8'd91,8'd230} : s = 38;
	{8'd91,8'd231} : s = 37;
	{8'd91,8'd232} : s = 135;
	{8'd91,8'd233} : s = 35;
	{8'd91,8'd234} : s = 120;
	{8'd91,8'd235} : s = 116;
	{8'd91,8'd236} : s = 244;
	{8'd91,8'd237} : s = 28;
	{8'd91,8'd238} : s = 114;
	{8'd91,8'd239} : s = 113;
	{8'd91,8'd240} : s = 242;
	{8'd91,8'd241} : s = 108;
	{8'd91,8'd242} : s = 241;
	{8'd91,8'd243} : s = 236;
	{8'd91,8'd244} : s = 399;
	{8'd91,8'd245} : s = 26;
	{8'd91,8'd246} : s = 106;
	{8'd91,8'd247} : s = 105;
	{8'd91,8'd248} : s = 234;
	{8'd91,8'd249} : s = 102;
	{8'd91,8'd250} : s = 233;
	{8'd91,8'd251} : s = 230;
	{8'd91,8'd252} : s = 380;
	{8'd91,8'd253} : s = 101;
	{8'd91,8'd254} : s = 229;
	{8'd91,8'd255} : s = 227;
	{8'd92,8'd0} : s = 354;
	{8'd92,8'd1} : s = 460;
	{8'd92,8'd2} : s = 458;
	{8'd92,8'd3} : s = 500;
	{8'd92,8'd4} : s = 65;
	{8'd92,8'd5} : s = 200;
	{8'd92,8'd6} : s = 196;
	{8'd92,8'd7} : s = 353;
	{8'd92,8'd8} : s = 194;
	{8'd92,8'd9} : s = 344;
	{8'd92,8'd10} : s = 340;
	{8'd92,8'd11} : s = 457;
	{8'd92,8'd12} : s = 193;
	{8'd92,8'd13} : s = 338;
	{8'd92,8'd14} : s = 337;
	{8'd92,8'd15} : s = 454;
	{8'd92,8'd16} : s = 332;
	{8'd92,8'd17} : s = 453;
	{8'd92,8'd18} : s = 451;
	{8'd92,8'd19} : s = 498;
	{8'd92,8'd20} : s = 176;
	{8'd92,8'd21} : s = 330;
	{8'd92,8'd22} : s = 329;
	{8'd92,8'd23} : s = 440;
	{8'd92,8'd24} : s = 326;
	{8'd92,8'd25} : s = 436;
	{8'd92,8'd26} : s = 434;
	{8'd92,8'd27} : s = 497;
	{8'd92,8'd28} : s = 325;
	{8'd92,8'd29} : s = 433;
	{8'd92,8'd30} : s = 428;
	{8'd92,8'd31} : s = 492;
	{8'd92,8'd32} : s = 426;
	{8'd92,8'd33} : s = 490;
	{8'd92,8'd34} : s = 489;
	{8'd92,8'd35} : s = 508;
	{8'd92,8'd36} : s = 2;
	{8'd92,8'd37} : s = 48;
	{8'd92,8'd38} : s = 40;
	{8'd92,8'd39} : s = 168;
	{8'd92,8'd40} : s = 36;
	{8'd92,8'd41} : s = 164;
	{8'd92,8'd42} : s = 162;
	{8'd92,8'd43} : s = 323;
	{8'd92,8'd44} : s = 34;
	{8'd92,8'd45} : s = 161;
	{8'd92,8'd46} : s = 152;
	{8'd92,8'd47} : s = 312;
	{8'd92,8'd48} : s = 148;
	{8'd92,8'd49} : s = 308;
	{8'd92,8'd50} : s = 306;
	{8'd92,8'd51} : s = 425;
	{8'd92,8'd52} : s = 33;
	{8'd92,8'd53} : s = 146;
	{8'd92,8'd54} : s = 145;
	{8'd92,8'd55} : s = 305;
	{8'd92,8'd56} : s = 140;
	{8'd92,8'd57} : s = 300;
	{8'd92,8'd58} : s = 298;
	{8'd92,8'd59} : s = 422;
	{8'd92,8'd60} : s = 138;
	{8'd92,8'd61} : s = 297;
	{8'd92,8'd62} : s = 294;
	{8'd92,8'd63} : s = 421;
	{8'd92,8'd64} : s = 293;
	{8'd92,8'd65} : s = 419;
	{8'd92,8'd66} : s = 412;
	{8'd92,8'd67} : s = 486;
	{8'd92,8'd68} : s = 24;
	{8'd92,8'd69} : s = 137;
	{8'd92,8'd70} : s = 134;
	{8'd92,8'd71} : s = 291;
	{8'd92,8'd72} : s = 133;
	{8'd92,8'd73} : s = 284;
	{8'd92,8'd74} : s = 282;
	{8'd92,8'd75} : s = 410;
	{8'd92,8'd76} : s = 131;
	{8'd92,8'd77} : s = 281;
	{8'd92,8'd78} : s = 278;
	{8'd92,8'd79} : s = 409;
	{8'd92,8'd80} : s = 277;
	{8'd92,8'd81} : s = 406;
	{8'd92,8'd82} : s = 405;
	{8'd92,8'd83} : s = 485;
	{8'd92,8'd84} : s = 112;
	{8'd92,8'd85} : s = 275;
	{8'd92,8'd86} : s = 270;
	{8'd92,8'd87} : s = 403;
	{8'd92,8'd88} : s = 269;
	{8'd92,8'd89} : s = 398;
	{8'd92,8'd90} : s = 397;
	{8'd92,8'd91} : s = 483;
	{8'd92,8'd92} : s = 267;
	{8'd92,8'd93} : s = 395;
	{8'd92,8'd94} : s = 391;
	{8'd92,8'd95} : s = 476;
	{8'd92,8'd96} : s = 376;
	{8'd92,8'd97} : s = 474;
	{8'd92,8'd98} : s = 473;
	{8'd92,8'd99} : s = 506;
	{8'd92,8'd100} : s = 20;
	{8'd92,8'd101} : s = 104;
	{8'd92,8'd102} : s = 100;
	{8'd92,8'd103} : s = 263;
	{8'd92,8'd104} : s = 98;
	{8'd92,8'd105} : s = 240;
	{8'd92,8'd106} : s = 232;
	{8'd92,8'd107} : s = 372;
	{8'd92,8'd108} : s = 97;
	{8'd92,8'd109} : s = 228;
	{8'd92,8'd110} : s = 226;
	{8'd92,8'd111} : s = 370;
	{8'd92,8'd112} : s = 225;
	{8'd92,8'd113} : s = 369;
	{8'd92,8'd114} : s = 364;
	{8'd92,8'd115} : s = 470;
	{8'd92,8'd116} : s = 88;
	{8'd92,8'd117} : s = 216;
	{8'd92,8'd118} : s = 212;
	{8'd92,8'd119} : s = 362;
	{8'd92,8'd120} : s = 210;
	{8'd92,8'd121} : s = 361;
	{8'd92,8'd122} : s = 358;
	{8'd92,8'd123} : s = 469;
	{8'd92,8'd124} : s = 209;
	{8'd92,8'd125} : s = 357;
	{8'd92,8'd126} : s = 355;
	{8'd92,8'd127} : s = 467;
	{8'd92,8'd128} : s = 348;
	{8'd92,8'd129} : s = 462;
	{8'd92,8'd130} : s = 461;
	{8'd92,8'd131} : s = 505;
	{8'd92,8'd132} : s = 84;
	{8'd92,8'd133} : s = 204;
	{8'd92,8'd134} : s = 202;
	{8'd92,8'd135} : s = 346;
	{8'd92,8'd136} : s = 201;
	{8'd92,8'd137} : s = 345;
	{8'd92,8'd138} : s = 342;
	{8'd92,8'd139} : s = 459;
	{8'd92,8'd140} : s = 198;
	{8'd92,8'd141} : s = 341;
	{8'd92,8'd142} : s = 339;
	{8'd92,8'd143} : s = 455;
	{8'd92,8'd144} : s = 334;
	{8'd92,8'd145} : s = 444;
	{8'd92,8'd146} : s = 442;
	{8'd92,8'd147} : s = 502;
	{8'd92,8'd148} : s = 197;
	{8'd92,8'd149} : s = 333;
	{8'd92,8'd150} : s = 331;
	{8'd92,8'd151} : s = 441;
	{8'd92,8'd152} : s = 327;
	{8'd92,8'd153} : s = 438;
	{8'd92,8'd154} : s = 437;
	{8'd92,8'd155} : s = 501;
	{8'd92,8'd156} : s = 316;
	{8'd92,8'd157} : s = 435;
	{8'd92,8'd158} : s = 430;
	{8'd92,8'd159} : s = 499;
	{8'd92,8'd160} : s = 429;
	{8'd92,8'd161} : s = 494;
	{8'd92,8'd162} : s = 493;
	{8'd92,8'd163} : s = 510;
	{8'd92,8'd164} : s = 1;
	{8'd92,8'd165} : s = 18;
	{8'd92,8'd166} : s = 17;
	{8'd92,8'd167} : s = 82;
	{8'd92,8'd168} : s = 12;
	{8'd92,8'd169} : s = 81;
	{8'd92,8'd170} : s = 76;
	{8'd92,8'd171} : s = 195;
	{8'd92,8'd172} : s = 10;
	{8'd92,8'd173} : s = 74;
	{8'd92,8'd174} : s = 73;
	{8'd92,8'd175} : s = 184;
	{8'd92,8'd176} : s = 70;
	{8'd92,8'd177} : s = 180;
	{8'd92,8'd178} : s = 178;
	{8'd92,8'd179} : s = 314;
	{8'd92,8'd180} : s = 9;
	{8'd92,8'd181} : s = 69;
	{8'd92,8'd182} : s = 67;
	{8'd92,8'd183} : s = 177;
	{8'd92,8'd184} : s = 56;
	{8'd92,8'd185} : s = 172;
	{8'd92,8'd186} : s = 170;
	{8'd92,8'd187} : s = 313;
	{8'd92,8'd188} : s = 52;
	{8'd92,8'd189} : s = 169;
	{8'd92,8'd190} : s = 166;
	{8'd92,8'd191} : s = 310;
	{8'd92,8'd192} : s = 165;
	{8'd92,8'd193} : s = 309;
	{8'd92,8'd194} : s = 307;
	{8'd92,8'd195} : s = 427;
	{8'd92,8'd196} : s = 6;
	{8'd92,8'd197} : s = 50;
	{8'd92,8'd198} : s = 49;
	{8'd92,8'd199} : s = 163;
	{8'd92,8'd200} : s = 44;
	{8'd92,8'd201} : s = 156;
	{8'd92,8'd202} : s = 154;
	{8'd92,8'd203} : s = 302;
	{8'd92,8'd204} : s = 42;
	{8'd92,8'd205} : s = 153;
	{8'd92,8'd206} : s = 150;
	{8'd92,8'd207} : s = 301;
	{8'd92,8'd208} : s = 149;
	{8'd92,8'd209} : s = 299;
	{8'd92,8'd210} : s = 295;
	{8'd92,8'd211} : s = 423;
	{8'd92,8'd212} : s = 41;
	{8'd92,8'd213} : s = 147;
	{8'd92,8'd214} : s = 142;
	{8'd92,8'd215} : s = 286;
	{8'd92,8'd216} : s = 141;
	{8'd92,8'd217} : s = 285;
	{8'd92,8'd218} : s = 283;
	{8'd92,8'd219} : s = 414;
	{8'd92,8'd220} : s = 139;
	{8'd92,8'd221} : s = 279;
	{8'd92,8'd222} : s = 271;
	{8'd92,8'd223} : s = 413;
	{8'd92,8'd224} : s = 248;
	{8'd92,8'd225} : s = 411;
	{8'd92,8'd226} : s = 407;
	{8'd92,8'd227} : s = 491;
	{8'd92,8'd228} : s = 5;
	{8'd92,8'd229} : s = 38;
	{8'd92,8'd230} : s = 37;
	{8'd92,8'd231} : s = 135;
	{8'd92,8'd232} : s = 35;
	{8'd92,8'd233} : s = 120;
	{8'd92,8'd234} : s = 116;
	{8'd92,8'd235} : s = 244;
	{8'd92,8'd236} : s = 28;
	{8'd92,8'd237} : s = 114;
	{8'd92,8'd238} : s = 113;
	{8'd92,8'd239} : s = 242;
	{8'd92,8'd240} : s = 108;
	{8'd92,8'd241} : s = 241;
	{8'd92,8'd242} : s = 236;
	{8'd92,8'd243} : s = 399;
	{8'd92,8'd244} : s = 26;
	{8'd92,8'd245} : s = 106;
	{8'd92,8'd246} : s = 105;
	{8'd92,8'd247} : s = 234;
	{8'd92,8'd248} : s = 102;
	{8'd92,8'd249} : s = 233;
	{8'd92,8'd250} : s = 230;
	{8'd92,8'd251} : s = 380;
	{8'd92,8'd252} : s = 101;
	{8'd92,8'd253} : s = 229;
	{8'd92,8'd254} : s = 227;
	{8'd92,8'd255} : s = 378;
	{8'd93,8'd0} : s = 460;
	{8'd93,8'd1} : s = 458;
	{8'd93,8'd2} : s = 500;
	{8'd93,8'd3} : s = 65;
	{8'd93,8'd4} : s = 200;
	{8'd93,8'd5} : s = 196;
	{8'd93,8'd6} : s = 353;
	{8'd93,8'd7} : s = 194;
	{8'd93,8'd8} : s = 344;
	{8'd93,8'd9} : s = 340;
	{8'd93,8'd10} : s = 457;
	{8'd93,8'd11} : s = 193;
	{8'd93,8'd12} : s = 338;
	{8'd93,8'd13} : s = 337;
	{8'd93,8'd14} : s = 454;
	{8'd93,8'd15} : s = 332;
	{8'd93,8'd16} : s = 453;
	{8'd93,8'd17} : s = 451;
	{8'd93,8'd18} : s = 498;
	{8'd93,8'd19} : s = 176;
	{8'd93,8'd20} : s = 330;
	{8'd93,8'd21} : s = 329;
	{8'd93,8'd22} : s = 440;
	{8'd93,8'd23} : s = 326;
	{8'd93,8'd24} : s = 436;
	{8'd93,8'd25} : s = 434;
	{8'd93,8'd26} : s = 497;
	{8'd93,8'd27} : s = 325;
	{8'd93,8'd28} : s = 433;
	{8'd93,8'd29} : s = 428;
	{8'd93,8'd30} : s = 492;
	{8'd93,8'd31} : s = 426;
	{8'd93,8'd32} : s = 490;
	{8'd93,8'd33} : s = 489;
	{8'd93,8'd34} : s = 508;
	{8'd93,8'd35} : s = 2;
	{8'd93,8'd36} : s = 48;
	{8'd93,8'd37} : s = 40;
	{8'd93,8'd38} : s = 168;
	{8'd93,8'd39} : s = 36;
	{8'd93,8'd40} : s = 164;
	{8'd93,8'd41} : s = 162;
	{8'd93,8'd42} : s = 323;
	{8'd93,8'd43} : s = 34;
	{8'd93,8'd44} : s = 161;
	{8'd93,8'd45} : s = 152;
	{8'd93,8'd46} : s = 312;
	{8'd93,8'd47} : s = 148;
	{8'd93,8'd48} : s = 308;
	{8'd93,8'd49} : s = 306;
	{8'd93,8'd50} : s = 425;
	{8'd93,8'd51} : s = 33;
	{8'd93,8'd52} : s = 146;
	{8'd93,8'd53} : s = 145;
	{8'd93,8'd54} : s = 305;
	{8'd93,8'd55} : s = 140;
	{8'd93,8'd56} : s = 300;
	{8'd93,8'd57} : s = 298;
	{8'd93,8'd58} : s = 422;
	{8'd93,8'd59} : s = 138;
	{8'd93,8'd60} : s = 297;
	{8'd93,8'd61} : s = 294;
	{8'd93,8'd62} : s = 421;
	{8'd93,8'd63} : s = 293;
	{8'd93,8'd64} : s = 419;
	{8'd93,8'd65} : s = 412;
	{8'd93,8'd66} : s = 486;
	{8'd93,8'd67} : s = 24;
	{8'd93,8'd68} : s = 137;
	{8'd93,8'd69} : s = 134;
	{8'd93,8'd70} : s = 291;
	{8'd93,8'd71} : s = 133;
	{8'd93,8'd72} : s = 284;
	{8'd93,8'd73} : s = 282;
	{8'd93,8'd74} : s = 410;
	{8'd93,8'd75} : s = 131;
	{8'd93,8'd76} : s = 281;
	{8'd93,8'd77} : s = 278;
	{8'd93,8'd78} : s = 409;
	{8'd93,8'd79} : s = 277;
	{8'd93,8'd80} : s = 406;
	{8'd93,8'd81} : s = 405;
	{8'd93,8'd82} : s = 485;
	{8'd93,8'd83} : s = 112;
	{8'd93,8'd84} : s = 275;
	{8'd93,8'd85} : s = 270;
	{8'd93,8'd86} : s = 403;
	{8'd93,8'd87} : s = 269;
	{8'd93,8'd88} : s = 398;
	{8'd93,8'd89} : s = 397;
	{8'd93,8'd90} : s = 483;
	{8'd93,8'd91} : s = 267;
	{8'd93,8'd92} : s = 395;
	{8'd93,8'd93} : s = 391;
	{8'd93,8'd94} : s = 476;
	{8'd93,8'd95} : s = 376;
	{8'd93,8'd96} : s = 474;
	{8'd93,8'd97} : s = 473;
	{8'd93,8'd98} : s = 506;
	{8'd93,8'd99} : s = 20;
	{8'd93,8'd100} : s = 104;
	{8'd93,8'd101} : s = 100;
	{8'd93,8'd102} : s = 263;
	{8'd93,8'd103} : s = 98;
	{8'd93,8'd104} : s = 240;
	{8'd93,8'd105} : s = 232;
	{8'd93,8'd106} : s = 372;
	{8'd93,8'd107} : s = 97;
	{8'd93,8'd108} : s = 228;
	{8'd93,8'd109} : s = 226;
	{8'd93,8'd110} : s = 370;
	{8'd93,8'd111} : s = 225;
	{8'd93,8'd112} : s = 369;
	{8'd93,8'd113} : s = 364;
	{8'd93,8'd114} : s = 470;
	{8'd93,8'd115} : s = 88;
	{8'd93,8'd116} : s = 216;
	{8'd93,8'd117} : s = 212;
	{8'd93,8'd118} : s = 362;
	{8'd93,8'd119} : s = 210;
	{8'd93,8'd120} : s = 361;
	{8'd93,8'd121} : s = 358;
	{8'd93,8'd122} : s = 469;
	{8'd93,8'd123} : s = 209;
	{8'd93,8'd124} : s = 357;
	{8'd93,8'd125} : s = 355;
	{8'd93,8'd126} : s = 467;
	{8'd93,8'd127} : s = 348;
	{8'd93,8'd128} : s = 462;
	{8'd93,8'd129} : s = 461;
	{8'd93,8'd130} : s = 505;
	{8'd93,8'd131} : s = 84;
	{8'd93,8'd132} : s = 204;
	{8'd93,8'd133} : s = 202;
	{8'd93,8'd134} : s = 346;
	{8'd93,8'd135} : s = 201;
	{8'd93,8'd136} : s = 345;
	{8'd93,8'd137} : s = 342;
	{8'd93,8'd138} : s = 459;
	{8'd93,8'd139} : s = 198;
	{8'd93,8'd140} : s = 341;
	{8'd93,8'd141} : s = 339;
	{8'd93,8'd142} : s = 455;
	{8'd93,8'd143} : s = 334;
	{8'd93,8'd144} : s = 444;
	{8'd93,8'd145} : s = 442;
	{8'd93,8'd146} : s = 502;
	{8'd93,8'd147} : s = 197;
	{8'd93,8'd148} : s = 333;
	{8'd93,8'd149} : s = 331;
	{8'd93,8'd150} : s = 441;
	{8'd93,8'd151} : s = 327;
	{8'd93,8'd152} : s = 438;
	{8'd93,8'd153} : s = 437;
	{8'd93,8'd154} : s = 501;
	{8'd93,8'd155} : s = 316;
	{8'd93,8'd156} : s = 435;
	{8'd93,8'd157} : s = 430;
	{8'd93,8'd158} : s = 499;
	{8'd93,8'd159} : s = 429;
	{8'd93,8'd160} : s = 494;
	{8'd93,8'd161} : s = 493;
	{8'd93,8'd162} : s = 510;
	{8'd93,8'd163} : s = 1;
	{8'd93,8'd164} : s = 18;
	{8'd93,8'd165} : s = 17;
	{8'd93,8'd166} : s = 82;
	{8'd93,8'd167} : s = 12;
	{8'd93,8'd168} : s = 81;
	{8'd93,8'd169} : s = 76;
	{8'd93,8'd170} : s = 195;
	{8'd93,8'd171} : s = 10;
	{8'd93,8'd172} : s = 74;
	{8'd93,8'd173} : s = 73;
	{8'd93,8'd174} : s = 184;
	{8'd93,8'd175} : s = 70;
	{8'd93,8'd176} : s = 180;
	{8'd93,8'd177} : s = 178;
	{8'd93,8'd178} : s = 314;
	{8'd93,8'd179} : s = 9;
	{8'd93,8'd180} : s = 69;
	{8'd93,8'd181} : s = 67;
	{8'd93,8'd182} : s = 177;
	{8'd93,8'd183} : s = 56;
	{8'd93,8'd184} : s = 172;
	{8'd93,8'd185} : s = 170;
	{8'd93,8'd186} : s = 313;
	{8'd93,8'd187} : s = 52;
	{8'd93,8'd188} : s = 169;
	{8'd93,8'd189} : s = 166;
	{8'd93,8'd190} : s = 310;
	{8'd93,8'd191} : s = 165;
	{8'd93,8'd192} : s = 309;
	{8'd93,8'd193} : s = 307;
	{8'd93,8'd194} : s = 427;
	{8'd93,8'd195} : s = 6;
	{8'd93,8'd196} : s = 50;
	{8'd93,8'd197} : s = 49;
	{8'd93,8'd198} : s = 163;
	{8'd93,8'd199} : s = 44;
	{8'd93,8'd200} : s = 156;
	{8'd93,8'd201} : s = 154;
	{8'd93,8'd202} : s = 302;
	{8'd93,8'd203} : s = 42;
	{8'd93,8'd204} : s = 153;
	{8'd93,8'd205} : s = 150;
	{8'd93,8'd206} : s = 301;
	{8'd93,8'd207} : s = 149;
	{8'd93,8'd208} : s = 299;
	{8'd93,8'd209} : s = 295;
	{8'd93,8'd210} : s = 423;
	{8'd93,8'd211} : s = 41;
	{8'd93,8'd212} : s = 147;
	{8'd93,8'd213} : s = 142;
	{8'd93,8'd214} : s = 286;
	{8'd93,8'd215} : s = 141;
	{8'd93,8'd216} : s = 285;
	{8'd93,8'd217} : s = 283;
	{8'd93,8'd218} : s = 414;
	{8'd93,8'd219} : s = 139;
	{8'd93,8'd220} : s = 279;
	{8'd93,8'd221} : s = 271;
	{8'd93,8'd222} : s = 413;
	{8'd93,8'd223} : s = 248;
	{8'd93,8'd224} : s = 411;
	{8'd93,8'd225} : s = 407;
	{8'd93,8'd226} : s = 491;
	{8'd93,8'd227} : s = 5;
	{8'd93,8'd228} : s = 38;
	{8'd93,8'd229} : s = 37;
	{8'd93,8'd230} : s = 135;
	{8'd93,8'd231} : s = 35;
	{8'd93,8'd232} : s = 120;
	{8'd93,8'd233} : s = 116;
	{8'd93,8'd234} : s = 244;
	{8'd93,8'd235} : s = 28;
	{8'd93,8'd236} : s = 114;
	{8'd93,8'd237} : s = 113;
	{8'd93,8'd238} : s = 242;
	{8'd93,8'd239} : s = 108;
	{8'd93,8'd240} : s = 241;
	{8'd93,8'd241} : s = 236;
	{8'd93,8'd242} : s = 399;
	{8'd93,8'd243} : s = 26;
	{8'd93,8'd244} : s = 106;
	{8'd93,8'd245} : s = 105;
	{8'd93,8'd246} : s = 234;
	{8'd93,8'd247} : s = 102;
	{8'd93,8'd248} : s = 233;
	{8'd93,8'd249} : s = 230;
	{8'd93,8'd250} : s = 380;
	{8'd93,8'd251} : s = 101;
	{8'd93,8'd252} : s = 229;
	{8'd93,8'd253} : s = 227;
	{8'd93,8'd254} : s = 378;
	{8'd93,8'd255} : s = 220;
	{8'd94,8'd0} : s = 458;
	{8'd94,8'd1} : s = 500;
	{8'd94,8'd2} : s = 65;
	{8'd94,8'd3} : s = 200;
	{8'd94,8'd4} : s = 196;
	{8'd94,8'd5} : s = 353;
	{8'd94,8'd6} : s = 194;
	{8'd94,8'd7} : s = 344;
	{8'd94,8'd8} : s = 340;
	{8'd94,8'd9} : s = 457;
	{8'd94,8'd10} : s = 193;
	{8'd94,8'd11} : s = 338;
	{8'd94,8'd12} : s = 337;
	{8'd94,8'd13} : s = 454;
	{8'd94,8'd14} : s = 332;
	{8'd94,8'd15} : s = 453;
	{8'd94,8'd16} : s = 451;
	{8'd94,8'd17} : s = 498;
	{8'd94,8'd18} : s = 176;
	{8'd94,8'd19} : s = 330;
	{8'd94,8'd20} : s = 329;
	{8'd94,8'd21} : s = 440;
	{8'd94,8'd22} : s = 326;
	{8'd94,8'd23} : s = 436;
	{8'd94,8'd24} : s = 434;
	{8'd94,8'd25} : s = 497;
	{8'd94,8'd26} : s = 325;
	{8'd94,8'd27} : s = 433;
	{8'd94,8'd28} : s = 428;
	{8'd94,8'd29} : s = 492;
	{8'd94,8'd30} : s = 426;
	{8'd94,8'd31} : s = 490;
	{8'd94,8'd32} : s = 489;
	{8'd94,8'd33} : s = 508;
	{8'd94,8'd34} : s = 2;
	{8'd94,8'd35} : s = 48;
	{8'd94,8'd36} : s = 40;
	{8'd94,8'd37} : s = 168;
	{8'd94,8'd38} : s = 36;
	{8'd94,8'd39} : s = 164;
	{8'd94,8'd40} : s = 162;
	{8'd94,8'd41} : s = 323;
	{8'd94,8'd42} : s = 34;
	{8'd94,8'd43} : s = 161;
	{8'd94,8'd44} : s = 152;
	{8'd94,8'd45} : s = 312;
	{8'd94,8'd46} : s = 148;
	{8'd94,8'd47} : s = 308;
	{8'd94,8'd48} : s = 306;
	{8'd94,8'd49} : s = 425;
	{8'd94,8'd50} : s = 33;
	{8'd94,8'd51} : s = 146;
	{8'd94,8'd52} : s = 145;
	{8'd94,8'd53} : s = 305;
	{8'd94,8'd54} : s = 140;
	{8'd94,8'd55} : s = 300;
	{8'd94,8'd56} : s = 298;
	{8'd94,8'd57} : s = 422;
	{8'd94,8'd58} : s = 138;
	{8'd94,8'd59} : s = 297;
	{8'd94,8'd60} : s = 294;
	{8'd94,8'd61} : s = 421;
	{8'd94,8'd62} : s = 293;
	{8'd94,8'd63} : s = 419;
	{8'd94,8'd64} : s = 412;
	{8'd94,8'd65} : s = 486;
	{8'd94,8'd66} : s = 24;
	{8'd94,8'd67} : s = 137;
	{8'd94,8'd68} : s = 134;
	{8'd94,8'd69} : s = 291;
	{8'd94,8'd70} : s = 133;
	{8'd94,8'd71} : s = 284;
	{8'd94,8'd72} : s = 282;
	{8'd94,8'd73} : s = 410;
	{8'd94,8'd74} : s = 131;
	{8'd94,8'd75} : s = 281;
	{8'd94,8'd76} : s = 278;
	{8'd94,8'd77} : s = 409;
	{8'd94,8'd78} : s = 277;
	{8'd94,8'd79} : s = 406;
	{8'd94,8'd80} : s = 405;
	{8'd94,8'd81} : s = 485;
	{8'd94,8'd82} : s = 112;
	{8'd94,8'd83} : s = 275;
	{8'd94,8'd84} : s = 270;
	{8'd94,8'd85} : s = 403;
	{8'd94,8'd86} : s = 269;
	{8'd94,8'd87} : s = 398;
	{8'd94,8'd88} : s = 397;
	{8'd94,8'd89} : s = 483;
	{8'd94,8'd90} : s = 267;
	{8'd94,8'd91} : s = 395;
	{8'd94,8'd92} : s = 391;
	{8'd94,8'd93} : s = 476;
	{8'd94,8'd94} : s = 376;
	{8'd94,8'd95} : s = 474;
	{8'd94,8'd96} : s = 473;
	{8'd94,8'd97} : s = 506;
	{8'd94,8'd98} : s = 20;
	{8'd94,8'd99} : s = 104;
	{8'd94,8'd100} : s = 100;
	{8'd94,8'd101} : s = 263;
	{8'd94,8'd102} : s = 98;
	{8'd94,8'd103} : s = 240;
	{8'd94,8'd104} : s = 232;
	{8'd94,8'd105} : s = 372;
	{8'd94,8'd106} : s = 97;
	{8'd94,8'd107} : s = 228;
	{8'd94,8'd108} : s = 226;
	{8'd94,8'd109} : s = 370;
	{8'd94,8'd110} : s = 225;
	{8'd94,8'd111} : s = 369;
	{8'd94,8'd112} : s = 364;
	{8'd94,8'd113} : s = 470;
	{8'd94,8'd114} : s = 88;
	{8'd94,8'd115} : s = 216;
	{8'd94,8'd116} : s = 212;
	{8'd94,8'd117} : s = 362;
	{8'd94,8'd118} : s = 210;
	{8'd94,8'd119} : s = 361;
	{8'd94,8'd120} : s = 358;
	{8'd94,8'd121} : s = 469;
	{8'd94,8'd122} : s = 209;
	{8'd94,8'd123} : s = 357;
	{8'd94,8'd124} : s = 355;
	{8'd94,8'd125} : s = 467;
	{8'd94,8'd126} : s = 348;
	{8'd94,8'd127} : s = 462;
	{8'd94,8'd128} : s = 461;
	{8'd94,8'd129} : s = 505;
	{8'd94,8'd130} : s = 84;
	{8'd94,8'd131} : s = 204;
	{8'd94,8'd132} : s = 202;
	{8'd94,8'd133} : s = 346;
	{8'd94,8'd134} : s = 201;
	{8'd94,8'd135} : s = 345;
	{8'd94,8'd136} : s = 342;
	{8'd94,8'd137} : s = 459;
	{8'd94,8'd138} : s = 198;
	{8'd94,8'd139} : s = 341;
	{8'd94,8'd140} : s = 339;
	{8'd94,8'd141} : s = 455;
	{8'd94,8'd142} : s = 334;
	{8'd94,8'd143} : s = 444;
	{8'd94,8'd144} : s = 442;
	{8'd94,8'd145} : s = 502;
	{8'd94,8'd146} : s = 197;
	{8'd94,8'd147} : s = 333;
	{8'd94,8'd148} : s = 331;
	{8'd94,8'd149} : s = 441;
	{8'd94,8'd150} : s = 327;
	{8'd94,8'd151} : s = 438;
	{8'd94,8'd152} : s = 437;
	{8'd94,8'd153} : s = 501;
	{8'd94,8'd154} : s = 316;
	{8'd94,8'd155} : s = 435;
	{8'd94,8'd156} : s = 430;
	{8'd94,8'd157} : s = 499;
	{8'd94,8'd158} : s = 429;
	{8'd94,8'd159} : s = 494;
	{8'd94,8'd160} : s = 493;
	{8'd94,8'd161} : s = 510;
	{8'd94,8'd162} : s = 1;
	{8'd94,8'd163} : s = 18;
	{8'd94,8'd164} : s = 17;
	{8'd94,8'd165} : s = 82;
	{8'd94,8'd166} : s = 12;
	{8'd94,8'd167} : s = 81;
	{8'd94,8'd168} : s = 76;
	{8'd94,8'd169} : s = 195;
	{8'd94,8'd170} : s = 10;
	{8'd94,8'd171} : s = 74;
	{8'd94,8'd172} : s = 73;
	{8'd94,8'd173} : s = 184;
	{8'd94,8'd174} : s = 70;
	{8'd94,8'd175} : s = 180;
	{8'd94,8'd176} : s = 178;
	{8'd94,8'd177} : s = 314;
	{8'd94,8'd178} : s = 9;
	{8'd94,8'd179} : s = 69;
	{8'd94,8'd180} : s = 67;
	{8'd94,8'd181} : s = 177;
	{8'd94,8'd182} : s = 56;
	{8'd94,8'd183} : s = 172;
	{8'd94,8'd184} : s = 170;
	{8'd94,8'd185} : s = 313;
	{8'd94,8'd186} : s = 52;
	{8'd94,8'd187} : s = 169;
	{8'd94,8'd188} : s = 166;
	{8'd94,8'd189} : s = 310;
	{8'd94,8'd190} : s = 165;
	{8'd94,8'd191} : s = 309;
	{8'd94,8'd192} : s = 307;
	{8'd94,8'd193} : s = 427;
	{8'd94,8'd194} : s = 6;
	{8'd94,8'd195} : s = 50;
	{8'd94,8'd196} : s = 49;
	{8'd94,8'd197} : s = 163;
	{8'd94,8'd198} : s = 44;
	{8'd94,8'd199} : s = 156;
	{8'd94,8'd200} : s = 154;
	{8'd94,8'd201} : s = 302;
	{8'd94,8'd202} : s = 42;
	{8'd94,8'd203} : s = 153;
	{8'd94,8'd204} : s = 150;
	{8'd94,8'd205} : s = 301;
	{8'd94,8'd206} : s = 149;
	{8'd94,8'd207} : s = 299;
	{8'd94,8'd208} : s = 295;
	{8'd94,8'd209} : s = 423;
	{8'd94,8'd210} : s = 41;
	{8'd94,8'd211} : s = 147;
	{8'd94,8'd212} : s = 142;
	{8'd94,8'd213} : s = 286;
	{8'd94,8'd214} : s = 141;
	{8'd94,8'd215} : s = 285;
	{8'd94,8'd216} : s = 283;
	{8'd94,8'd217} : s = 414;
	{8'd94,8'd218} : s = 139;
	{8'd94,8'd219} : s = 279;
	{8'd94,8'd220} : s = 271;
	{8'd94,8'd221} : s = 413;
	{8'd94,8'd222} : s = 248;
	{8'd94,8'd223} : s = 411;
	{8'd94,8'd224} : s = 407;
	{8'd94,8'd225} : s = 491;
	{8'd94,8'd226} : s = 5;
	{8'd94,8'd227} : s = 38;
	{8'd94,8'd228} : s = 37;
	{8'd94,8'd229} : s = 135;
	{8'd94,8'd230} : s = 35;
	{8'd94,8'd231} : s = 120;
	{8'd94,8'd232} : s = 116;
	{8'd94,8'd233} : s = 244;
	{8'd94,8'd234} : s = 28;
	{8'd94,8'd235} : s = 114;
	{8'd94,8'd236} : s = 113;
	{8'd94,8'd237} : s = 242;
	{8'd94,8'd238} : s = 108;
	{8'd94,8'd239} : s = 241;
	{8'd94,8'd240} : s = 236;
	{8'd94,8'd241} : s = 399;
	{8'd94,8'd242} : s = 26;
	{8'd94,8'd243} : s = 106;
	{8'd94,8'd244} : s = 105;
	{8'd94,8'd245} : s = 234;
	{8'd94,8'd246} : s = 102;
	{8'd94,8'd247} : s = 233;
	{8'd94,8'd248} : s = 230;
	{8'd94,8'd249} : s = 380;
	{8'd94,8'd250} : s = 101;
	{8'd94,8'd251} : s = 229;
	{8'd94,8'd252} : s = 227;
	{8'd94,8'd253} : s = 378;
	{8'd94,8'd254} : s = 220;
	{8'd94,8'd255} : s = 377;
	{8'd95,8'd0} : s = 500;
	{8'd95,8'd1} : s = 65;
	{8'd95,8'd2} : s = 200;
	{8'd95,8'd3} : s = 196;
	{8'd95,8'd4} : s = 353;
	{8'd95,8'd5} : s = 194;
	{8'd95,8'd6} : s = 344;
	{8'd95,8'd7} : s = 340;
	{8'd95,8'd8} : s = 457;
	{8'd95,8'd9} : s = 193;
	{8'd95,8'd10} : s = 338;
	{8'd95,8'd11} : s = 337;
	{8'd95,8'd12} : s = 454;
	{8'd95,8'd13} : s = 332;
	{8'd95,8'd14} : s = 453;
	{8'd95,8'd15} : s = 451;
	{8'd95,8'd16} : s = 498;
	{8'd95,8'd17} : s = 176;
	{8'd95,8'd18} : s = 330;
	{8'd95,8'd19} : s = 329;
	{8'd95,8'd20} : s = 440;
	{8'd95,8'd21} : s = 326;
	{8'd95,8'd22} : s = 436;
	{8'd95,8'd23} : s = 434;
	{8'd95,8'd24} : s = 497;
	{8'd95,8'd25} : s = 325;
	{8'd95,8'd26} : s = 433;
	{8'd95,8'd27} : s = 428;
	{8'd95,8'd28} : s = 492;
	{8'd95,8'd29} : s = 426;
	{8'd95,8'd30} : s = 490;
	{8'd95,8'd31} : s = 489;
	{8'd95,8'd32} : s = 508;
	{8'd95,8'd33} : s = 2;
	{8'd95,8'd34} : s = 48;
	{8'd95,8'd35} : s = 40;
	{8'd95,8'd36} : s = 168;
	{8'd95,8'd37} : s = 36;
	{8'd95,8'd38} : s = 164;
	{8'd95,8'd39} : s = 162;
	{8'd95,8'd40} : s = 323;
	{8'd95,8'd41} : s = 34;
	{8'd95,8'd42} : s = 161;
	{8'd95,8'd43} : s = 152;
	{8'd95,8'd44} : s = 312;
	{8'd95,8'd45} : s = 148;
	{8'd95,8'd46} : s = 308;
	{8'd95,8'd47} : s = 306;
	{8'd95,8'd48} : s = 425;
	{8'd95,8'd49} : s = 33;
	{8'd95,8'd50} : s = 146;
	{8'd95,8'd51} : s = 145;
	{8'd95,8'd52} : s = 305;
	{8'd95,8'd53} : s = 140;
	{8'd95,8'd54} : s = 300;
	{8'd95,8'd55} : s = 298;
	{8'd95,8'd56} : s = 422;
	{8'd95,8'd57} : s = 138;
	{8'd95,8'd58} : s = 297;
	{8'd95,8'd59} : s = 294;
	{8'd95,8'd60} : s = 421;
	{8'd95,8'd61} : s = 293;
	{8'd95,8'd62} : s = 419;
	{8'd95,8'd63} : s = 412;
	{8'd95,8'd64} : s = 486;
	{8'd95,8'd65} : s = 24;
	{8'd95,8'd66} : s = 137;
	{8'd95,8'd67} : s = 134;
	{8'd95,8'd68} : s = 291;
	{8'd95,8'd69} : s = 133;
	{8'd95,8'd70} : s = 284;
	{8'd95,8'd71} : s = 282;
	{8'd95,8'd72} : s = 410;
	{8'd95,8'd73} : s = 131;
	{8'd95,8'd74} : s = 281;
	{8'd95,8'd75} : s = 278;
	{8'd95,8'd76} : s = 409;
	{8'd95,8'd77} : s = 277;
	{8'd95,8'd78} : s = 406;
	{8'd95,8'd79} : s = 405;
	{8'd95,8'd80} : s = 485;
	{8'd95,8'd81} : s = 112;
	{8'd95,8'd82} : s = 275;
	{8'd95,8'd83} : s = 270;
	{8'd95,8'd84} : s = 403;
	{8'd95,8'd85} : s = 269;
	{8'd95,8'd86} : s = 398;
	{8'd95,8'd87} : s = 397;
	{8'd95,8'd88} : s = 483;
	{8'd95,8'd89} : s = 267;
	{8'd95,8'd90} : s = 395;
	{8'd95,8'd91} : s = 391;
	{8'd95,8'd92} : s = 476;
	{8'd95,8'd93} : s = 376;
	{8'd95,8'd94} : s = 474;
	{8'd95,8'd95} : s = 473;
	{8'd95,8'd96} : s = 506;
	{8'd95,8'd97} : s = 20;
	{8'd95,8'd98} : s = 104;
	{8'd95,8'd99} : s = 100;
	{8'd95,8'd100} : s = 263;
	{8'd95,8'd101} : s = 98;
	{8'd95,8'd102} : s = 240;
	{8'd95,8'd103} : s = 232;
	{8'd95,8'd104} : s = 372;
	{8'd95,8'd105} : s = 97;
	{8'd95,8'd106} : s = 228;
	{8'd95,8'd107} : s = 226;
	{8'd95,8'd108} : s = 370;
	{8'd95,8'd109} : s = 225;
	{8'd95,8'd110} : s = 369;
	{8'd95,8'd111} : s = 364;
	{8'd95,8'd112} : s = 470;
	{8'd95,8'd113} : s = 88;
	{8'd95,8'd114} : s = 216;
	{8'd95,8'd115} : s = 212;
	{8'd95,8'd116} : s = 362;
	{8'd95,8'd117} : s = 210;
	{8'd95,8'd118} : s = 361;
	{8'd95,8'd119} : s = 358;
	{8'd95,8'd120} : s = 469;
	{8'd95,8'd121} : s = 209;
	{8'd95,8'd122} : s = 357;
	{8'd95,8'd123} : s = 355;
	{8'd95,8'd124} : s = 467;
	{8'd95,8'd125} : s = 348;
	{8'd95,8'd126} : s = 462;
	{8'd95,8'd127} : s = 461;
	{8'd95,8'd128} : s = 505;
	{8'd95,8'd129} : s = 84;
	{8'd95,8'd130} : s = 204;
	{8'd95,8'd131} : s = 202;
	{8'd95,8'd132} : s = 346;
	{8'd95,8'd133} : s = 201;
	{8'd95,8'd134} : s = 345;
	{8'd95,8'd135} : s = 342;
	{8'd95,8'd136} : s = 459;
	{8'd95,8'd137} : s = 198;
	{8'd95,8'd138} : s = 341;
	{8'd95,8'd139} : s = 339;
	{8'd95,8'd140} : s = 455;
	{8'd95,8'd141} : s = 334;
	{8'd95,8'd142} : s = 444;
	{8'd95,8'd143} : s = 442;
	{8'd95,8'd144} : s = 502;
	{8'd95,8'd145} : s = 197;
	{8'd95,8'd146} : s = 333;
	{8'd95,8'd147} : s = 331;
	{8'd95,8'd148} : s = 441;
	{8'd95,8'd149} : s = 327;
	{8'd95,8'd150} : s = 438;
	{8'd95,8'd151} : s = 437;
	{8'd95,8'd152} : s = 501;
	{8'd95,8'd153} : s = 316;
	{8'd95,8'd154} : s = 435;
	{8'd95,8'd155} : s = 430;
	{8'd95,8'd156} : s = 499;
	{8'd95,8'd157} : s = 429;
	{8'd95,8'd158} : s = 494;
	{8'd95,8'd159} : s = 493;
	{8'd95,8'd160} : s = 510;
	{8'd95,8'd161} : s = 1;
	{8'd95,8'd162} : s = 18;
	{8'd95,8'd163} : s = 17;
	{8'd95,8'd164} : s = 82;
	{8'd95,8'd165} : s = 12;
	{8'd95,8'd166} : s = 81;
	{8'd95,8'd167} : s = 76;
	{8'd95,8'd168} : s = 195;
	{8'd95,8'd169} : s = 10;
	{8'd95,8'd170} : s = 74;
	{8'd95,8'd171} : s = 73;
	{8'd95,8'd172} : s = 184;
	{8'd95,8'd173} : s = 70;
	{8'd95,8'd174} : s = 180;
	{8'd95,8'd175} : s = 178;
	{8'd95,8'd176} : s = 314;
	{8'd95,8'd177} : s = 9;
	{8'd95,8'd178} : s = 69;
	{8'd95,8'd179} : s = 67;
	{8'd95,8'd180} : s = 177;
	{8'd95,8'd181} : s = 56;
	{8'd95,8'd182} : s = 172;
	{8'd95,8'd183} : s = 170;
	{8'd95,8'd184} : s = 313;
	{8'd95,8'd185} : s = 52;
	{8'd95,8'd186} : s = 169;
	{8'd95,8'd187} : s = 166;
	{8'd95,8'd188} : s = 310;
	{8'd95,8'd189} : s = 165;
	{8'd95,8'd190} : s = 309;
	{8'd95,8'd191} : s = 307;
	{8'd95,8'd192} : s = 427;
	{8'd95,8'd193} : s = 6;
	{8'd95,8'd194} : s = 50;
	{8'd95,8'd195} : s = 49;
	{8'd95,8'd196} : s = 163;
	{8'd95,8'd197} : s = 44;
	{8'd95,8'd198} : s = 156;
	{8'd95,8'd199} : s = 154;
	{8'd95,8'd200} : s = 302;
	{8'd95,8'd201} : s = 42;
	{8'd95,8'd202} : s = 153;
	{8'd95,8'd203} : s = 150;
	{8'd95,8'd204} : s = 301;
	{8'd95,8'd205} : s = 149;
	{8'd95,8'd206} : s = 299;
	{8'd95,8'd207} : s = 295;
	{8'd95,8'd208} : s = 423;
	{8'd95,8'd209} : s = 41;
	{8'd95,8'd210} : s = 147;
	{8'd95,8'd211} : s = 142;
	{8'd95,8'd212} : s = 286;
	{8'd95,8'd213} : s = 141;
	{8'd95,8'd214} : s = 285;
	{8'd95,8'd215} : s = 283;
	{8'd95,8'd216} : s = 414;
	{8'd95,8'd217} : s = 139;
	{8'd95,8'd218} : s = 279;
	{8'd95,8'd219} : s = 271;
	{8'd95,8'd220} : s = 413;
	{8'd95,8'd221} : s = 248;
	{8'd95,8'd222} : s = 411;
	{8'd95,8'd223} : s = 407;
	{8'd95,8'd224} : s = 491;
	{8'd95,8'd225} : s = 5;
	{8'd95,8'd226} : s = 38;
	{8'd95,8'd227} : s = 37;
	{8'd95,8'd228} : s = 135;
	{8'd95,8'd229} : s = 35;
	{8'd95,8'd230} : s = 120;
	{8'd95,8'd231} : s = 116;
	{8'd95,8'd232} : s = 244;
	{8'd95,8'd233} : s = 28;
	{8'd95,8'd234} : s = 114;
	{8'd95,8'd235} : s = 113;
	{8'd95,8'd236} : s = 242;
	{8'd95,8'd237} : s = 108;
	{8'd95,8'd238} : s = 241;
	{8'd95,8'd239} : s = 236;
	{8'd95,8'd240} : s = 399;
	{8'd95,8'd241} : s = 26;
	{8'd95,8'd242} : s = 106;
	{8'd95,8'd243} : s = 105;
	{8'd95,8'd244} : s = 234;
	{8'd95,8'd245} : s = 102;
	{8'd95,8'd246} : s = 233;
	{8'd95,8'd247} : s = 230;
	{8'd95,8'd248} : s = 380;
	{8'd95,8'd249} : s = 101;
	{8'd95,8'd250} : s = 229;
	{8'd95,8'd251} : s = 227;
	{8'd95,8'd252} : s = 378;
	{8'd95,8'd253} : s = 220;
	{8'd95,8'd254} : s = 377;
	{8'd95,8'd255} : s = 374;
	{8'd96,8'd0} : s = 65;
	{8'd96,8'd1} : s = 200;
	{8'd96,8'd2} : s = 196;
	{8'd96,8'd3} : s = 353;
	{8'd96,8'd4} : s = 194;
	{8'd96,8'd5} : s = 344;
	{8'd96,8'd6} : s = 340;
	{8'd96,8'd7} : s = 457;
	{8'd96,8'd8} : s = 193;
	{8'd96,8'd9} : s = 338;
	{8'd96,8'd10} : s = 337;
	{8'd96,8'd11} : s = 454;
	{8'd96,8'd12} : s = 332;
	{8'd96,8'd13} : s = 453;
	{8'd96,8'd14} : s = 451;
	{8'd96,8'd15} : s = 498;
	{8'd96,8'd16} : s = 176;
	{8'd96,8'd17} : s = 330;
	{8'd96,8'd18} : s = 329;
	{8'd96,8'd19} : s = 440;
	{8'd96,8'd20} : s = 326;
	{8'd96,8'd21} : s = 436;
	{8'd96,8'd22} : s = 434;
	{8'd96,8'd23} : s = 497;
	{8'd96,8'd24} : s = 325;
	{8'd96,8'd25} : s = 433;
	{8'd96,8'd26} : s = 428;
	{8'd96,8'd27} : s = 492;
	{8'd96,8'd28} : s = 426;
	{8'd96,8'd29} : s = 490;
	{8'd96,8'd30} : s = 489;
	{8'd96,8'd31} : s = 508;
	{8'd96,8'd32} : s = 2;
	{8'd96,8'd33} : s = 48;
	{8'd96,8'd34} : s = 40;
	{8'd96,8'd35} : s = 168;
	{8'd96,8'd36} : s = 36;
	{8'd96,8'd37} : s = 164;
	{8'd96,8'd38} : s = 162;
	{8'd96,8'd39} : s = 323;
	{8'd96,8'd40} : s = 34;
	{8'd96,8'd41} : s = 161;
	{8'd96,8'd42} : s = 152;
	{8'd96,8'd43} : s = 312;
	{8'd96,8'd44} : s = 148;
	{8'd96,8'd45} : s = 308;
	{8'd96,8'd46} : s = 306;
	{8'd96,8'd47} : s = 425;
	{8'd96,8'd48} : s = 33;
	{8'd96,8'd49} : s = 146;
	{8'd96,8'd50} : s = 145;
	{8'd96,8'd51} : s = 305;
	{8'd96,8'd52} : s = 140;
	{8'd96,8'd53} : s = 300;
	{8'd96,8'd54} : s = 298;
	{8'd96,8'd55} : s = 422;
	{8'd96,8'd56} : s = 138;
	{8'd96,8'd57} : s = 297;
	{8'd96,8'd58} : s = 294;
	{8'd96,8'd59} : s = 421;
	{8'd96,8'd60} : s = 293;
	{8'd96,8'd61} : s = 419;
	{8'd96,8'd62} : s = 412;
	{8'd96,8'd63} : s = 486;
	{8'd96,8'd64} : s = 24;
	{8'd96,8'd65} : s = 137;
	{8'd96,8'd66} : s = 134;
	{8'd96,8'd67} : s = 291;
	{8'd96,8'd68} : s = 133;
	{8'd96,8'd69} : s = 284;
	{8'd96,8'd70} : s = 282;
	{8'd96,8'd71} : s = 410;
	{8'd96,8'd72} : s = 131;
	{8'd96,8'd73} : s = 281;
	{8'd96,8'd74} : s = 278;
	{8'd96,8'd75} : s = 409;
	{8'd96,8'd76} : s = 277;
	{8'd96,8'd77} : s = 406;
	{8'd96,8'd78} : s = 405;
	{8'd96,8'd79} : s = 485;
	{8'd96,8'd80} : s = 112;
	{8'd96,8'd81} : s = 275;
	{8'd96,8'd82} : s = 270;
	{8'd96,8'd83} : s = 403;
	{8'd96,8'd84} : s = 269;
	{8'd96,8'd85} : s = 398;
	{8'd96,8'd86} : s = 397;
	{8'd96,8'd87} : s = 483;
	{8'd96,8'd88} : s = 267;
	{8'd96,8'd89} : s = 395;
	{8'd96,8'd90} : s = 391;
	{8'd96,8'd91} : s = 476;
	{8'd96,8'd92} : s = 376;
	{8'd96,8'd93} : s = 474;
	{8'd96,8'd94} : s = 473;
	{8'd96,8'd95} : s = 506;
	{8'd96,8'd96} : s = 20;
	{8'd96,8'd97} : s = 104;
	{8'd96,8'd98} : s = 100;
	{8'd96,8'd99} : s = 263;
	{8'd96,8'd100} : s = 98;
	{8'd96,8'd101} : s = 240;
	{8'd96,8'd102} : s = 232;
	{8'd96,8'd103} : s = 372;
	{8'd96,8'd104} : s = 97;
	{8'd96,8'd105} : s = 228;
	{8'd96,8'd106} : s = 226;
	{8'd96,8'd107} : s = 370;
	{8'd96,8'd108} : s = 225;
	{8'd96,8'd109} : s = 369;
	{8'd96,8'd110} : s = 364;
	{8'd96,8'd111} : s = 470;
	{8'd96,8'd112} : s = 88;
	{8'd96,8'd113} : s = 216;
	{8'd96,8'd114} : s = 212;
	{8'd96,8'd115} : s = 362;
	{8'd96,8'd116} : s = 210;
	{8'd96,8'd117} : s = 361;
	{8'd96,8'd118} : s = 358;
	{8'd96,8'd119} : s = 469;
	{8'd96,8'd120} : s = 209;
	{8'd96,8'd121} : s = 357;
	{8'd96,8'd122} : s = 355;
	{8'd96,8'd123} : s = 467;
	{8'd96,8'd124} : s = 348;
	{8'd96,8'd125} : s = 462;
	{8'd96,8'd126} : s = 461;
	{8'd96,8'd127} : s = 505;
	{8'd96,8'd128} : s = 84;
	{8'd96,8'd129} : s = 204;
	{8'd96,8'd130} : s = 202;
	{8'd96,8'd131} : s = 346;
	{8'd96,8'd132} : s = 201;
	{8'd96,8'd133} : s = 345;
	{8'd96,8'd134} : s = 342;
	{8'd96,8'd135} : s = 459;
	{8'd96,8'd136} : s = 198;
	{8'd96,8'd137} : s = 341;
	{8'd96,8'd138} : s = 339;
	{8'd96,8'd139} : s = 455;
	{8'd96,8'd140} : s = 334;
	{8'd96,8'd141} : s = 444;
	{8'd96,8'd142} : s = 442;
	{8'd96,8'd143} : s = 502;
	{8'd96,8'd144} : s = 197;
	{8'd96,8'd145} : s = 333;
	{8'd96,8'd146} : s = 331;
	{8'd96,8'd147} : s = 441;
	{8'd96,8'd148} : s = 327;
	{8'd96,8'd149} : s = 438;
	{8'd96,8'd150} : s = 437;
	{8'd96,8'd151} : s = 501;
	{8'd96,8'd152} : s = 316;
	{8'd96,8'd153} : s = 435;
	{8'd96,8'd154} : s = 430;
	{8'd96,8'd155} : s = 499;
	{8'd96,8'd156} : s = 429;
	{8'd96,8'd157} : s = 494;
	{8'd96,8'd158} : s = 493;
	{8'd96,8'd159} : s = 510;
	{8'd96,8'd160} : s = 1;
	{8'd96,8'd161} : s = 18;
	{8'd96,8'd162} : s = 17;
	{8'd96,8'd163} : s = 82;
	{8'd96,8'd164} : s = 12;
	{8'd96,8'd165} : s = 81;
	{8'd96,8'd166} : s = 76;
	{8'd96,8'd167} : s = 195;
	{8'd96,8'd168} : s = 10;
	{8'd96,8'd169} : s = 74;
	{8'd96,8'd170} : s = 73;
	{8'd96,8'd171} : s = 184;
	{8'd96,8'd172} : s = 70;
	{8'd96,8'd173} : s = 180;
	{8'd96,8'd174} : s = 178;
	{8'd96,8'd175} : s = 314;
	{8'd96,8'd176} : s = 9;
	{8'd96,8'd177} : s = 69;
	{8'd96,8'd178} : s = 67;
	{8'd96,8'd179} : s = 177;
	{8'd96,8'd180} : s = 56;
	{8'd96,8'd181} : s = 172;
	{8'd96,8'd182} : s = 170;
	{8'd96,8'd183} : s = 313;
	{8'd96,8'd184} : s = 52;
	{8'd96,8'd185} : s = 169;
	{8'd96,8'd186} : s = 166;
	{8'd96,8'd187} : s = 310;
	{8'd96,8'd188} : s = 165;
	{8'd96,8'd189} : s = 309;
	{8'd96,8'd190} : s = 307;
	{8'd96,8'd191} : s = 427;
	{8'd96,8'd192} : s = 6;
	{8'd96,8'd193} : s = 50;
	{8'd96,8'd194} : s = 49;
	{8'd96,8'd195} : s = 163;
	{8'd96,8'd196} : s = 44;
	{8'd96,8'd197} : s = 156;
	{8'd96,8'd198} : s = 154;
	{8'd96,8'd199} : s = 302;
	{8'd96,8'd200} : s = 42;
	{8'd96,8'd201} : s = 153;
	{8'd96,8'd202} : s = 150;
	{8'd96,8'd203} : s = 301;
	{8'd96,8'd204} : s = 149;
	{8'd96,8'd205} : s = 299;
	{8'd96,8'd206} : s = 295;
	{8'd96,8'd207} : s = 423;
	{8'd96,8'd208} : s = 41;
	{8'd96,8'd209} : s = 147;
	{8'd96,8'd210} : s = 142;
	{8'd96,8'd211} : s = 286;
	{8'd96,8'd212} : s = 141;
	{8'd96,8'd213} : s = 285;
	{8'd96,8'd214} : s = 283;
	{8'd96,8'd215} : s = 414;
	{8'd96,8'd216} : s = 139;
	{8'd96,8'd217} : s = 279;
	{8'd96,8'd218} : s = 271;
	{8'd96,8'd219} : s = 413;
	{8'd96,8'd220} : s = 248;
	{8'd96,8'd221} : s = 411;
	{8'd96,8'd222} : s = 407;
	{8'd96,8'd223} : s = 491;
	{8'd96,8'd224} : s = 5;
	{8'd96,8'd225} : s = 38;
	{8'd96,8'd226} : s = 37;
	{8'd96,8'd227} : s = 135;
	{8'd96,8'd228} : s = 35;
	{8'd96,8'd229} : s = 120;
	{8'd96,8'd230} : s = 116;
	{8'd96,8'd231} : s = 244;
	{8'd96,8'd232} : s = 28;
	{8'd96,8'd233} : s = 114;
	{8'd96,8'd234} : s = 113;
	{8'd96,8'd235} : s = 242;
	{8'd96,8'd236} : s = 108;
	{8'd96,8'd237} : s = 241;
	{8'd96,8'd238} : s = 236;
	{8'd96,8'd239} : s = 399;
	{8'd96,8'd240} : s = 26;
	{8'd96,8'd241} : s = 106;
	{8'd96,8'd242} : s = 105;
	{8'd96,8'd243} : s = 234;
	{8'd96,8'd244} : s = 102;
	{8'd96,8'd245} : s = 233;
	{8'd96,8'd246} : s = 230;
	{8'd96,8'd247} : s = 380;
	{8'd96,8'd248} : s = 101;
	{8'd96,8'd249} : s = 229;
	{8'd96,8'd250} : s = 227;
	{8'd96,8'd251} : s = 378;
	{8'd96,8'd252} : s = 220;
	{8'd96,8'd253} : s = 377;
	{8'd96,8'd254} : s = 374;
	{8'd96,8'd255} : s = 487;
	{8'd97,8'd0} : s = 200;
	{8'd97,8'd1} : s = 196;
	{8'd97,8'd2} : s = 353;
	{8'd97,8'd3} : s = 194;
	{8'd97,8'd4} : s = 344;
	{8'd97,8'd5} : s = 340;
	{8'd97,8'd6} : s = 457;
	{8'd97,8'd7} : s = 193;
	{8'd97,8'd8} : s = 338;
	{8'd97,8'd9} : s = 337;
	{8'd97,8'd10} : s = 454;
	{8'd97,8'd11} : s = 332;
	{8'd97,8'd12} : s = 453;
	{8'd97,8'd13} : s = 451;
	{8'd97,8'd14} : s = 498;
	{8'd97,8'd15} : s = 176;
	{8'd97,8'd16} : s = 330;
	{8'd97,8'd17} : s = 329;
	{8'd97,8'd18} : s = 440;
	{8'd97,8'd19} : s = 326;
	{8'd97,8'd20} : s = 436;
	{8'd97,8'd21} : s = 434;
	{8'd97,8'd22} : s = 497;
	{8'd97,8'd23} : s = 325;
	{8'd97,8'd24} : s = 433;
	{8'd97,8'd25} : s = 428;
	{8'd97,8'd26} : s = 492;
	{8'd97,8'd27} : s = 426;
	{8'd97,8'd28} : s = 490;
	{8'd97,8'd29} : s = 489;
	{8'd97,8'd30} : s = 508;
	{8'd97,8'd31} : s = 2;
	{8'd97,8'd32} : s = 48;
	{8'd97,8'd33} : s = 40;
	{8'd97,8'd34} : s = 168;
	{8'd97,8'd35} : s = 36;
	{8'd97,8'd36} : s = 164;
	{8'd97,8'd37} : s = 162;
	{8'd97,8'd38} : s = 323;
	{8'd97,8'd39} : s = 34;
	{8'd97,8'd40} : s = 161;
	{8'd97,8'd41} : s = 152;
	{8'd97,8'd42} : s = 312;
	{8'd97,8'd43} : s = 148;
	{8'd97,8'd44} : s = 308;
	{8'd97,8'd45} : s = 306;
	{8'd97,8'd46} : s = 425;
	{8'd97,8'd47} : s = 33;
	{8'd97,8'd48} : s = 146;
	{8'd97,8'd49} : s = 145;
	{8'd97,8'd50} : s = 305;
	{8'd97,8'd51} : s = 140;
	{8'd97,8'd52} : s = 300;
	{8'd97,8'd53} : s = 298;
	{8'd97,8'd54} : s = 422;
	{8'd97,8'd55} : s = 138;
	{8'd97,8'd56} : s = 297;
	{8'd97,8'd57} : s = 294;
	{8'd97,8'd58} : s = 421;
	{8'd97,8'd59} : s = 293;
	{8'd97,8'd60} : s = 419;
	{8'd97,8'd61} : s = 412;
	{8'd97,8'd62} : s = 486;
	{8'd97,8'd63} : s = 24;
	{8'd97,8'd64} : s = 137;
	{8'd97,8'd65} : s = 134;
	{8'd97,8'd66} : s = 291;
	{8'd97,8'd67} : s = 133;
	{8'd97,8'd68} : s = 284;
	{8'd97,8'd69} : s = 282;
	{8'd97,8'd70} : s = 410;
	{8'd97,8'd71} : s = 131;
	{8'd97,8'd72} : s = 281;
	{8'd97,8'd73} : s = 278;
	{8'd97,8'd74} : s = 409;
	{8'd97,8'd75} : s = 277;
	{8'd97,8'd76} : s = 406;
	{8'd97,8'd77} : s = 405;
	{8'd97,8'd78} : s = 485;
	{8'd97,8'd79} : s = 112;
	{8'd97,8'd80} : s = 275;
	{8'd97,8'd81} : s = 270;
	{8'd97,8'd82} : s = 403;
	{8'd97,8'd83} : s = 269;
	{8'd97,8'd84} : s = 398;
	{8'd97,8'd85} : s = 397;
	{8'd97,8'd86} : s = 483;
	{8'd97,8'd87} : s = 267;
	{8'd97,8'd88} : s = 395;
	{8'd97,8'd89} : s = 391;
	{8'd97,8'd90} : s = 476;
	{8'd97,8'd91} : s = 376;
	{8'd97,8'd92} : s = 474;
	{8'd97,8'd93} : s = 473;
	{8'd97,8'd94} : s = 506;
	{8'd97,8'd95} : s = 20;
	{8'd97,8'd96} : s = 104;
	{8'd97,8'd97} : s = 100;
	{8'd97,8'd98} : s = 263;
	{8'd97,8'd99} : s = 98;
	{8'd97,8'd100} : s = 240;
	{8'd97,8'd101} : s = 232;
	{8'd97,8'd102} : s = 372;
	{8'd97,8'd103} : s = 97;
	{8'd97,8'd104} : s = 228;
	{8'd97,8'd105} : s = 226;
	{8'd97,8'd106} : s = 370;
	{8'd97,8'd107} : s = 225;
	{8'd97,8'd108} : s = 369;
	{8'd97,8'd109} : s = 364;
	{8'd97,8'd110} : s = 470;
	{8'd97,8'd111} : s = 88;
	{8'd97,8'd112} : s = 216;
	{8'd97,8'd113} : s = 212;
	{8'd97,8'd114} : s = 362;
	{8'd97,8'd115} : s = 210;
	{8'd97,8'd116} : s = 361;
	{8'd97,8'd117} : s = 358;
	{8'd97,8'd118} : s = 469;
	{8'd97,8'd119} : s = 209;
	{8'd97,8'd120} : s = 357;
	{8'd97,8'd121} : s = 355;
	{8'd97,8'd122} : s = 467;
	{8'd97,8'd123} : s = 348;
	{8'd97,8'd124} : s = 462;
	{8'd97,8'd125} : s = 461;
	{8'd97,8'd126} : s = 505;
	{8'd97,8'd127} : s = 84;
	{8'd97,8'd128} : s = 204;
	{8'd97,8'd129} : s = 202;
	{8'd97,8'd130} : s = 346;
	{8'd97,8'd131} : s = 201;
	{8'd97,8'd132} : s = 345;
	{8'd97,8'd133} : s = 342;
	{8'd97,8'd134} : s = 459;
	{8'd97,8'd135} : s = 198;
	{8'd97,8'd136} : s = 341;
	{8'd97,8'd137} : s = 339;
	{8'd97,8'd138} : s = 455;
	{8'd97,8'd139} : s = 334;
	{8'd97,8'd140} : s = 444;
	{8'd97,8'd141} : s = 442;
	{8'd97,8'd142} : s = 502;
	{8'd97,8'd143} : s = 197;
	{8'd97,8'd144} : s = 333;
	{8'd97,8'd145} : s = 331;
	{8'd97,8'd146} : s = 441;
	{8'd97,8'd147} : s = 327;
	{8'd97,8'd148} : s = 438;
	{8'd97,8'd149} : s = 437;
	{8'd97,8'd150} : s = 501;
	{8'd97,8'd151} : s = 316;
	{8'd97,8'd152} : s = 435;
	{8'd97,8'd153} : s = 430;
	{8'd97,8'd154} : s = 499;
	{8'd97,8'd155} : s = 429;
	{8'd97,8'd156} : s = 494;
	{8'd97,8'd157} : s = 493;
	{8'd97,8'd158} : s = 510;
	{8'd97,8'd159} : s = 1;
	{8'd97,8'd160} : s = 18;
	{8'd97,8'd161} : s = 17;
	{8'd97,8'd162} : s = 82;
	{8'd97,8'd163} : s = 12;
	{8'd97,8'd164} : s = 81;
	{8'd97,8'd165} : s = 76;
	{8'd97,8'd166} : s = 195;
	{8'd97,8'd167} : s = 10;
	{8'd97,8'd168} : s = 74;
	{8'd97,8'd169} : s = 73;
	{8'd97,8'd170} : s = 184;
	{8'd97,8'd171} : s = 70;
	{8'd97,8'd172} : s = 180;
	{8'd97,8'd173} : s = 178;
	{8'd97,8'd174} : s = 314;
	{8'd97,8'd175} : s = 9;
	{8'd97,8'd176} : s = 69;
	{8'd97,8'd177} : s = 67;
	{8'd97,8'd178} : s = 177;
	{8'd97,8'd179} : s = 56;
	{8'd97,8'd180} : s = 172;
	{8'd97,8'd181} : s = 170;
	{8'd97,8'd182} : s = 313;
	{8'd97,8'd183} : s = 52;
	{8'd97,8'd184} : s = 169;
	{8'd97,8'd185} : s = 166;
	{8'd97,8'd186} : s = 310;
	{8'd97,8'd187} : s = 165;
	{8'd97,8'd188} : s = 309;
	{8'd97,8'd189} : s = 307;
	{8'd97,8'd190} : s = 427;
	{8'd97,8'd191} : s = 6;
	{8'd97,8'd192} : s = 50;
	{8'd97,8'd193} : s = 49;
	{8'd97,8'd194} : s = 163;
	{8'd97,8'd195} : s = 44;
	{8'd97,8'd196} : s = 156;
	{8'd97,8'd197} : s = 154;
	{8'd97,8'd198} : s = 302;
	{8'd97,8'd199} : s = 42;
	{8'd97,8'd200} : s = 153;
	{8'd97,8'd201} : s = 150;
	{8'd97,8'd202} : s = 301;
	{8'd97,8'd203} : s = 149;
	{8'd97,8'd204} : s = 299;
	{8'd97,8'd205} : s = 295;
	{8'd97,8'd206} : s = 423;
	{8'd97,8'd207} : s = 41;
	{8'd97,8'd208} : s = 147;
	{8'd97,8'd209} : s = 142;
	{8'd97,8'd210} : s = 286;
	{8'd97,8'd211} : s = 141;
	{8'd97,8'd212} : s = 285;
	{8'd97,8'd213} : s = 283;
	{8'd97,8'd214} : s = 414;
	{8'd97,8'd215} : s = 139;
	{8'd97,8'd216} : s = 279;
	{8'd97,8'd217} : s = 271;
	{8'd97,8'd218} : s = 413;
	{8'd97,8'd219} : s = 248;
	{8'd97,8'd220} : s = 411;
	{8'd97,8'd221} : s = 407;
	{8'd97,8'd222} : s = 491;
	{8'd97,8'd223} : s = 5;
	{8'd97,8'd224} : s = 38;
	{8'd97,8'd225} : s = 37;
	{8'd97,8'd226} : s = 135;
	{8'd97,8'd227} : s = 35;
	{8'd97,8'd228} : s = 120;
	{8'd97,8'd229} : s = 116;
	{8'd97,8'd230} : s = 244;
	{8'd97,8'd231} : s = 28;
	{8'd97,8'd232} : s = 114;
	{8'd97,8'd233} : s = 113;
	{8'd97,8'd234} : s = 242;
	{8'd97,8'd235} : s = 108;
	{8'd97,8'd236} : s = 241;
	{8'd97,8'd237} : s = 236;
	{8'd97,8'd238} : s = 399;
	{8'd97,8'd239} : s = 26;
	{8'd97,8'd240} : s = 106;
	{8'd97,8'd241} : s = 105;
	{8'd97,8'd242} : s = 234;
	{8'd97,8'd243} : s = 102;
	{8'd97,8'd244} : s = 233;
	{8'd97,8'd245} : s = 230;
	{8'd97,8'd246} : s = 380;
	{8'd97,8'd247} : s = 101;
	{8'd97,8'd248} : s = 229;
	{8'd97,8'd249} : s = 227;
	{8'd97,8'd250} : s = 378;
	{8'd97,8'd251} : s = 220;
	{8'd97,8'd252} : s = 377;
	{8'd97,8'd253} : s = 374;
	{8'd97,8'd254} : s = 487;
	{8'd97,8'd255} : s = 25;
	{8'd98,8'd0} : s = 196;
	{8'd98,8'd1} : s = 353;
	{8'd98,8'd2} : s = 194;
	{8'd98,8'd3} : s = 344;
	{8'd98,8'd4} : s = 340;
	{8'd98,8'd5} : s = 457;
	{8'd98,8'd6} : s = 193;
	{8'd98,8'd7} : s = 338;
	{8'd98,8'd8} : s = 337;
	{8'd98,8'd9} : s = 454;
	{8'd98,8'd10} : s = 332;
	{8'd98,8'd11} : s = 453;
	{8'd98,8'd12} : s = 451;
	{8'd98,8'd13} : s = 498;
	{8'd98,8'd14} : s = 176;
	{8'd98,8'd15} : s = 330;
	{8'd98,8'd16} : s = 329;
	{8'd98,8'd17} : s = 440;
	{8'd98,8'd18} : s = 326;
	{8'd98,8'd19} : s = 436;
	{8'd98,8'd20} : s = 434;
	{8'd98,8'd21} : s = 497;
	{8'd98,8'd22} : s = 325;
	{8'd98,8'd23} : s = 433;
	{8'd98,8'd24} : s = 428;
	{8'd98,8'd25} : s = 492;
	{8'd98,8'd26} : s = 426;
	{8'd98,8'd27} : s = 490;
	{8'd98,8'd28} : s = 489;
	{8'd98,8'd29} : s = 508;
	{8'd98,8'd30} : s = 2;
	{8'd98,8'd31} : s = 48;
	{8'd98,8'd32} : s = 40;
	{8'd98,8'd33} : s = 168;
	{8'd98,8'd34} : s = 36;
	{8'd98,8'd35} : s = 164;
	{8'd98,8'd36} : s = 162;
	{8'd98,8'd37} : s = 323;
	{8'd98,8'd38} : s = 34;
	{8'd98,8'd39} : s = 161;
	{8'd98,8'd40} : s = 152;
	{8'd98,8'd41} : s = 312;
	{8'd98,8'd42} : s = 148;
	{8'd98,8'd43} : s = 308;
	{8'd98,8'd44} : s = 306;
	{8'd98,8'd45} : s = 425;
	{8'd98,8'd46} : s = 33;
	{8'd98,8'd47} : s = 146;
	{8'd98,8'd48} : s = 145;
	{8'd98,8'd49} : s = 305;
	{8'd98,8'd50} : s = 140;
	{8'd98,8'd51} : s = 300;
	{8'd98,8'd52} : s = 298;
	{8'd98,8'd53} : s = 422;
	{8'd98,8'd54} : s = 138;
	{8'd98,8'd55} : s = 297;
	{8'd98,8'd56} : s = 294;
	{8'd98,8'd57} : s = 421;
	{8'd98,8'd58} : s = 293;
	{8'd98,8'd59} : s = 419;
	{8'd98,8'd60} : s = 412;
	{8'd98,8'd61} : s = 486;
	{8'd98,8'd62} : s = 24;
	{8'd98,8'd63} : s = 137;
	{8'd98,8'd64} : s = 134;
	{8'd98,8'd65} : s = 291;
	{8'd98,8'd66} : s = 133;
	{8'd98,8'd67} : s = 284;
	{8'd98,8'd68} : s = 282;
	{8'd98,8'd69} : s = 410;
	{8'd98,8'd70} : s = 131;
	{8'd98,8'd71} : s = 281;
	{8'd98,8'd72} : s = 278;
	{8'd98,8'd73} : s = 409;
	{8'd98,8'd74} : s = 277;
	{8'd98,8'd75} : s = 406;
	{8'd98,8'd76} : s = 405;
	{8'd98,8'd77} : s = 485;
	{8'd98,8'd78} : s = 112;
	{8'd98,8'd79} : s = 275;
	{8'd98,8'd80} : s = 270;
	{8'd98,8'd81} : s = 403;
	{8'd98,8'd82} : s = 269;
	{8'd98,8'd83} : s = 398;
	{8'd98,8'd84} : s = 397;
	{8'd98,8'd85} : s = 483;
	{8'd98,8'd86} : s = 267;
	{8'd98,8'd87} : s = 395;
	{8'd98,8'd88} : s = 391;
	{8'd98,8'd89} : s = 476;
	{8'd98,8'd90} : s = 376;
	{8'd98,8'd91} : s = 474;
	{8'd98,8'd92} : s = 473;
	{8'd98,8'd93} : s = 506;
	{8'd98,8'd94} : s = 20;
	{8'd98,8'd95} : s = 104;
	{8'd98,8'd96} : s = 100;
	{8'd98,8'd97} : s = 263;
	{8'd98,8'd98} : s = 98;
	{8'd98,8'd99} : s = 240;
	{8'd98,8'd100} : s = 232;
	{8'd98,8'd101} : s = 372;
	{8'd98,8'd102} : s = 97;
	{8'd98,8'd103} : s = 228;
	{8'd98,8'd104} : s = 226;
	{8'd98,8'd105} : s = 370;
	{8'd98,8'd106} : s = 225;
	{8'd98,8'd107} : s = 369;
	{8'd98,8'd108} : s = 364;
	{8'd98,8'd109} : s = 470;
	{8'd98,8'd110} : s = 88;
	{8'd98,8'd111} : s = 216;
	{8'd98,8'd112} : s = 212;
	{8'd98,8'd113} : s = 362;
	{8'd98,8'd114} : s = 210;
	{8'd98,8'd115} : s = 361;
	{8'd98,8'd116} : s = 358;
	{8'd98,8'd117} : s = 469;
	{8'd98,8'd118} : s = 209;
	{8'd98,8'd119} : s = 357;
	{8'd98,8'd120} : s = 355;
	{8'd98,8'd121} : s = 467;
	{8'd98,8'd122} : s = 348;
	{8'd98,8'd123} : s = 462;
	{8'd98,8'd124} : s = 461;
	{8'd98,8'd125} : s = 505;
	{8'd98,8'd126} : s = 84;
	{8'd98,8'd127} : s = 204;
	{8'd98,8'd128} : s = 202;
	{8'd98,8'd129} : s = 346;
	{8'd98,8'd130} : s = 201;
	{8'd98,8'd131} : s = 345;
	{8'd98,8'd132} : s = 342;
	{8'd98,8'd133} : s = 459;
	{8'd98,8'd134} : s = 198;
	{8'd98,8'd135} : s = 341;
	{8'd98,8'd136} : s = 339;
	{8'd98,8'd137} : s = 455;
	{8'd98,8'd138} : s = 334;
	{8'd98,8'd139} : s = 444;
	{8'd98,8'd140} : s = 442;
	{8'd98,8'd141} : s = 502;
	{8'd98,8'd142} : s = 197;
	{8'd98,8'd143} : s = 333;
	{8'd98,8'd144} : s = 331;
	{8'd98,8'd145} : s = 441;
	{8'd98,8'd146} : s = 327;
	{8'd98,8'd147} : s = 438;
	{8'd98,8'd148} : s = 437;
	{8'd98,8'd149} : s = 501;
	{8'd98,8'd150} : s = 316;
	{8'd98,8'd151} : s = 435;
	{8'd98,8'd152} : s = 430;
	{8'd98,8'd153} : s = 499;
	{8'd98,8'd154} : s = 429;
	{8'd98,8'd155} : s = 494;
	{8'd98,8'd156} : s = 493;
	{8'd98,8'd157} : s = 510;
	{8'd98,8'd158} : s = 1;
	{8'd98,8'd159} : s = 18;
	{8'd98,8'd160} : s = 17;
	{8'd98,8'd161} : s = 82;
	{8'd98,8'd162} : s = 12;
	{8'd98,8'd163} : s = 81;
	{8'd98,8'd164} : s = 76;
	{8'd98,8'd165} : s = 195;
	{8'd98,8'd166} : s = 10;
	{8'd98,8'd167} : s = 74;
	{8'd98,8'd168} : s = 73;
	{8'd98,8'd169} : s = 184;
	{8'd98,8'd170} : s = 70;
	{8'd98,8'd171} : s = 180;
	{8'd98,8'd172} : s = 178;
	{8'd98,8'd173} : s = 314;
	{8'd98,8'd174} : s = 9;
	{8'd98,8'd175} : s = 69;
	{8'd98,8'd176} : s = 67;
	{8'd98,8'd177} : s = 177;
	{8'd98,8'd178} : s = 56;
	{8'd98,8'd179} : s = 172;
	{8'd98,8'd180} : s = 170;
	{8'd98,8'd181} : s = 313;
	{8'd98,8'd182} : s = 52;
	{8'd98,8'd183} : s = 169;
	{8'd98,8'd184} : s = 166;
	{8'd98,8'd185} : s = 310;
	{8'd98,8'd186} : s = 165;
	{8'd98,8'd187} : s = 309;
	{8'd98,8'd188} : s = 307;
	{8'd98,8'd189} : s = 427;
	{8'd98,8'd190} : s = 6;
	{8'd98,8'd191} : s = 50;
	{8'd98,8'd192} : s = 49;
	{8'd98,8'd193} : s = 163;
	{8'd98,8'd194} : s = 44;
	{8'd98,8'd195} : s = 156;
	{8'd98,8'd196} : s = 154;
	{8'd98,8'd197} : s = 302;
	{8'd98,8'd198} : s = 42;
	{8'd98,8'd199} : s = 153;
	{8'd98,8'd200} : s = 150;
	{8'd98,8'd201} : s = 301;
	{8'd98,8'd202} : s = 149;
	{8'd98,8'd203} : s = 299;
	{8'd98,8'd204} : s = 295;
	{8'd98,8'd205} : s = 423;
	{8'd98,8'd206} : s = 41;
	{8'd98,8'd207} : s = 147;
	{8'd98,8'd208} : s = 142;
	{8'd98,8'd209} : s = 286;
	{8'd98,8'd210} : s = 141;
	{8'd98,8'd211} : s = 285;
	{8'd98,8'd212} : s = 283;
	{8'd98,8'd213} : s = 414;
	{8'd98,8'd214} : s = 139;
	{8'd98,8'd215} : s = 279;
	{8'd98,8'd216} : s = 271;
	{8'd98,8'd217} : s = 413;
	{8'd98,8'd218} : s = 248;
	{8'd98,8'd219} : s = 411;
	{8'd98,8'd220} : s = 407;
	{8'd98,8'd221} : s = 491;
	{8'd98,8'd222} : s = 5;
	{8'd98,8'd223} : s = 38;
	{8'd98,8'd224} : s = 37;
	{8'd98,8'd225} : s = 135;
	{8'd98,8'd226} : s = 35;
	{8'd98,8'd227} : s = 120;
	{8'd98,8'd228} : s = 116;
	{8'd98,8'd229} : s = 244;
	{8'd98,8'd230} : s = 28;
	{8'd98,8'd231} : s = 114;
	{8'd98,8'd232} : s = 113;
	{8'd98,8'd233} : s = 242;
	{8'd98,8'd234} : s = 108;
	{8'd98,8'd235} : s = 241;
	{8'd98,8'd236} : s = 236;
	{8'd98,8'd237} : s = 399;
	{8'd98,8'd238} : s = 26;
	{8'd98,8'd239} : s = 106;
	{8'd98,8'd240} : s = 105;
	{8'd98,8'd241} : s = 234;
	{8'd98,8'd242} : s = 102;
	{8'd98,8'd243} : s = 233;
	{8'd98,8'd244} : s = 230;
	{8'd98,8'd245} : s = 380;
	{8'd98,8'd246} : s = 101;
	{8'd98,8'd247} : s = 229;
	{8'd98,8'd248} : s = 227;
	{8'd98,8'd249} : s = 378;
	{8'd98,8'd250} : s = 220;
	{8'd98,8'd251} : s = 377;
	{8'd98,8'd252} : s = 374;
	{8'd98,8'd253} : s = 487;
	{8'd98,8'd254} : s = 25;
	{8'd98,8'd255} : s = 99;
	{8'd99,8'd0} : s = 353;
	{8'd99,8'd1} : s = 194;
	{8'd99,8'd2} : s = 344;
	{8'd99,8'd3} : s = 340;
	{8'd99,8'd4} : s = 457;
	{8'd99,8'd5} : s = 193;
	{8'd99,8'd6} : s = 338;
	{8'd99,8'd7} : s = 337;
	{8'd99,8'd8} : s = 454;
	{8'd99,8'd9} : s = 332;
	{8'd99,8'd10} : s = 453;
	{8'd99,8'd11} : s = 451;
	{8'd99,8'd12} : s = 498;
	{8'd99,8'd13} : s = 176;
	{8'd99,8'd14} : s = 330;
	{8'd99,8'd15} : s = 329;
	{8'd99,8'd16} : s = 440;
	{8'd99,8'd17} : s = 326;
	{8'd99,8'd18} : s = 436;
	{8'd99,8'd19} : s = 434;
	{8'd99,8'd20} : s = 497;
	{8'd99,8'd21} : s = 325;
	{8'd99,8'd22} : s = 433;
	{8'd99,8'd23} : s = 428;
	{8'd99,8'd24} : s = 492;
	{8'd99,8'd25} : s = 426;
	{8'd99,8'd26} : s = 490;
	{8'd99,8'd27} : s = 489;
	{8'd99,8'd28} : s = 508;
	{8'd99,8'd29} : s = 2;
	{8'd99,8'd30} : s = 48;
	{8'd99,8'd31} : s = 40;
	{8'd99,8'd32} : s = 168;
	{8'd99,8'd33} : s = 36;
	{8'd99,8'd34} : s = 164;
	{8'd99,8'd35} : s = 162;
	{8'd99,8'd36} : s = 323;
	{8'd99,8'd37} : s = 34;
	{8'd99,8'd38} : s = 161;
	{8'd99,8'd39} : s = 152;
	{8'd99,8'd40} : s = 312;
	{8'd99,8'd41} : s = 148;
	{8'd99,8'd42} : s = 308;
	{8'd99,8'd43} : s = 306;
	{8'd99,8'd44} : s = 425;
	{8'd99,8'd45} : s = 33;
	{8'd99,8'd46} : s = 146;
	{8'd99,8'd47} : s = 145;
	{8'd99,8'd48} : s = 305;
	{8'd99,8'd49} : s = 140;
	{8'd99,8'd50} : s = 300;
	{8'd99,8'd51} : s = 298;
	{8'd99,8'd52} : s = 422;
	{8'd99,8'd53} : s = 138;
	{8'd99,8'd54} : s = 297;
	{8'd99,8'd55} : s = 294;
	{8'd99,8'd56} : s = 421;
	{8'd99,8'd57} : s = 293;
	{8'd99,8'd58} : s = 419;
	{8'd99,8'd59} : s = 412;
	{8'd99,8'd60} : s = 486;
	{8'd99,8'd61} : s = 24;
	{8'd99,8'd62} : s = 137;
	{8'd99,8'd63} : s = 134;
	{8'd99,8'd64} : s = 291;
	{8'd99,8'd65} : s = 133;
	{8'd99,8'd66} : s = 284;
	{8'd99,8'd67} : s = 282;
	{8'd99,8'd68} : s = 410;
	{8'd99,8'd69} : s = 131;
	{8'd99,8'd70} : s = 281;
	{8'd99,8'd71} : s = 278;
	{8'd99,8'd72} : s = 409;
	{8'd99,8'd73} : s = 277;
	{8'd99,8'd74} : s = 406;
	{8'd99,8'd75} : s = 405;
	{8'd99,8'd76} : s = 485;
	{8'd99,8'd77} : s = 112;
	{8'd99,8'd78} : s = 275;
	{8'd99,8'd79} : s = 270;
	{8'd99,8'd80} : s = 403;
	{8'd99,8'd81} : s = 269;
	{8'd99,8'd82} : s = 398;
	{8'd99,8'd83} : s = 397;
	{8'd99,8'd84} : s = 483;
	{8'd99,8'd85} : s = 267;
	{8'd99,8'd86} : s = 395;
	{8'd99,8'd87} : s = 391;
	{8'd99,8'd88} : s = 476;
	{8'd99,8'd89} : s = 376;
	{8'd99,8'd90} : s = 474;
	{8'd99,8'd91} : s = 473;
	{8'd99,8'd92} : s = 506;
	{8'd99,8'd93} : s = 20;
	{8'd99,8'd94} : s = 104;
	{8'd99,8'd95} : s = 100;
	{8'd99,8'd96} : s = 263;
	{8'd99,8'd97} : s = 98;
	{8'd99,8'd98} : s = 240;
	{8'd99,8'd99} : s = 232;
	{8'd99,8'd100} : s = 372;
	{8'd99,8'd101} : s = 97;
	{8'd99,8'd102} : s = 228;
	{8'd99,8'd103} : s = 226;
	{8'd99,8'd104} : s = 370;
	{8'd99,8'd105} : s = 225;
	{8'd99,8'd106} : s = 369;
	{8'd99,8'd107} : s = 364;
	{8'd99,8'd108} : s = 470;
	{8'd99,8'd109} : s = 88;
	{8'd99,8'd110} : s = 216;
	{8'd99,8'd111} : s = 212;
	{8'd99,8'd112} : s = 362;
	{8'd99,8'd113} : s = 210;
	{8'd99,8'd114} : s = 361;
	{8'd99,8'd115} : s = 358;
	{8'd99,8'd116} : s = 469;
	{8'd99,8'd117} : s = 209;
	{8'd99,8'd118} : s = 357;
	{8'd99,8'd119} : s = 355;
	{8'd99,8'd120} : s = 467;
	{8'd99,8'd121} : s = 348;
	{8'd99,8'd122} : s = 462;
	{8'd99,8'd123} : s = 461;
	{8'd99,8'd124} : s = 505;
	{8'd99,8'd125} : s = 84;
	{8'd99,8'd126} : s = 204;
	{8'd99,8'd127} : s = 202;
	{8'd99,8'd128} : s = 346;
	{8'd99,8'd129} : s = 201;
	{8'd99,8'd130} : s = 345;
	{8'd99,8'd131} : s = 342;
	{8'd99,8'd132} : s = 459;
	{8'd99,8'd133} : s = 198;
	{8'd99,8'd134} : s = 341;
	{8'd99,8'd135} : s = 339;
	{8'd99,8'd136} : s = 455;
	{8'd99,8'd137} : s = 334;
	{8'd99,8'd138} : s = 444;
	{8'd99,8'd139} : s = 442;
	{8'd99,8'd140} : s = 502;
	{8'd99,8'd141} : s = 197;
	{8'd99,8'd142} : s = 333;
	{8'd99,8'd143} : s = 331;
	{8'd99,8'd144} : s = 441;
	{8'd99,8'd145} : s = 327;
	{8'd99,8'd146} : s = 438;
	{8'd99,8'd147} : s = 437;
	{8'd99,8'd148} : s = 501;
	{8'd99,8'd149} : s = 316;
	{8'd99,8'd150} : s = 435;
	{8'd99,8'd151} : s = 430;
	{8'd99,8'd152} : s = 499;
	{8'd99,8'd153} : s = 429;
	{8'd99,8'd154} : s = 494;
	{8'd99,8'd155} : s = 493;
	{8'd99,8'd156} : s = 510;
	{8'd99,8'd157} : s = 1;
	{8'd99,8'd158} : s = 18;
	{8'd99,8'd159} : s = 17;
	{8'd99,8'd160} : s = 82;
	{8'd99,8'd161} : s = 12;
	{8'd99,8'd162} : s = 81;
	{8'd99,8'd163} : s = 76;
	{8'd99,8'd164} : s = 195;
	{8'd99,8'd165} : s = 10;
	{8'd99,8'd166} : s = 74;
	{8'd99,8'd167} : s = 73;
	{8'd99,8'd168} : s = 184;
	{8'd99,8'd169} : s = 70;
	{8'd99,8'd170} : s = 180;
	{8'd99,8'd171} : s = 178;
	{8'd99,8'd172} : s = 314;
	{8'd99,8'd173} : s = 9;
	{8'd99,8'd174} : s = 69;
	{8'd99,8'd175} : s = 67;
	{8'd99,8'd176} : s = 177;
	{8'd99,8'd177} : s = 56;
	{8'd99,8'd178} : s = 172;
	{8'd99,8'd179} : s = 170;
	{8'd99,8'd180} : s = 313;
	{8'd99,8'd181} : s = 52;
	{8'd99,8'd182} : s = 169;
	{8'd99,8'd183} : s = 166;
	{8'd99,8'd184} : s = 310;
	{8'd99,8'd185} : s = 165;
	{8'd99,8'd186} : s = 309;
	{8'd99,8'd187} : s = 307;
	{8'd99,8'd188} : s = 427;
	{8'd99,8'd189} : s = 6;
	{8'd99,8'd190} : s = 50;
	{8'd99,8'd191} : s = 49;
	{8'd99,8'd192} : s = 163;
	{8'd99,8'd193} : s = 44;
	{8'd99,8'd194} : s = 156;
	{8'd99,8'd195} : s = 154;
	{8'd99,8'd196} : s = 302;
	{8'd99,8'd197} : s = 42;
	{8'd99,8'd198} : s = 153;
	{8'd99,8'd199} : s = 150;
	{8'd99,8'd200} : s = 301;
	{8'd99,8'd201} : s = 149;
	{8'd99,8'd202} : s = 299;
	{8'd99,8'd203} : s = 295;
	{8'd99,8'd204} : s = 423;
	{8'd99,8'd205} : s = 41;
	{8'd99,8'd206} : s = 147;
	{8'd99,8'd207} : s = 142;
	{8'd99,8'd208} : s = 286;
	{8'd99,8'd209} : s = 141;
	{8'd99,8'd210} : s = 285;
	{8'd99,8'd211} : s = 283;
	{8'd99,8'd212} : s = 414;
	{8'd99,8'd213} : s = 139;
	{8'd99,8'd214} : s = 279;
	{8'd99,8'd215} : s = 271;
	{8'd99,8'd216} : s = 413;
	{8'd99,8'd217} : s = 248;
	{8'd99,8'd218} : s = 411;
	{8'd99,8'd219} : s = 407;
	{8'd99,8'd220} : s = 491;
	{8'd99,8'd221} : s = 5;
	{8'd99,8'd222} : s = 38;
	{8'd99,8'd223} : s = 37;
	{8'd99,8'd224} : s = 135;
	{8'd99,8'd225} : s = 35;
	{8'd99,8'd226} : s = 120;
	{8'd99,8'd227} : s = 116;
	{8'd99,8'd228} : s = 244;
	{8'd99,8'd229} : s = 28;
	{8'd99,8'd230} : s = 114;
	{8'd99,8'd231} : s = 113;
	{8'd99,8'd232} : s = 242;
	{8'd99,8'd233} : s = 108;
	{8'd99,8'd234} : s = 241;
	{8'd99,8'd235} : s = 236;
	{8'd99,8'd236} : s = 399;
	{8'd99,8'd237} : s = 26;
	{8'd99,8'd238} : s = 106;
	{8'd99,8'd239} : s = 105;
	{8'd99,8'd240} : s = 234;
	{8'd99,8'd241} : s = 102;
	{8'd99,8'd242} : s = 233;
	{8'd99,8'd243} : s = 230;
	{8'd99,8'd244} : s = 380;
	{8'd99,8'd245} : s = 101;
	{8'd99,8'd246} : s = 229;
	{8'd99,8'd247} : s = 227;
	{8'd99,8'd248} : s = 378;
	{8'd99,8'd249} : s = 220;
	{8'd99,8'd250} : s = 377;
	{8'd99,8'd251} : s = 374;
	{8'd99,8'd252} : s = 487;
	{8'd99,8'd253} : s = 25;
	{8'd99,8'd254} : s = 99;
	{8'd99,8'd255} : s = 92;
	{8'd100,8'd0} : s = 194;
	{8'd100,8'd1} : s = 344;
	{8'd100,8'd2} : s = 340;
	{8'd100,8'd3} : s = 457;
	{8'd100,8'd4} : s = 193;
	{8'd100,8'd5} : s = 338;
	{8'd100,8'd6} : s = 337;
	{8'd100,8'd7} : s = 454;
	{8'd100,8'd8} : s = 332;
	{8'd100,8'd9} : s = 453;
	{8'd100,8'd10} : s = 451;
	{8'd100,8'd11} : s = 498;
	{8'd100,8'd12} : s = 176;
	{8'd100,8'd13} : s = 330;
	{8'd100,8'd14} : s = 329;
	{8'd100,8'd15} : s = 440;
	{8'd100,8'd16} : s = 326;
	{8'd100,8'd17} : s = 436;
	{8'd100,8'd18} : s = 434;
	{8'd100,8'd19} : s = 497;
	{8'd100,8'd20} : s = 325;
	{8'd100,8'd21} : s = 433;
	{8'd100,8'd22} : s = 428;
	{8'd100,8'd23} : s = 492;
	{8'd100,8'd24} : s = 426;
	{8'd100,8'd25} : s = 490;
	{8'd100,8'd26} : s = 489;
	{8'd100,8'd27} : s = 508;
	{8'd100,8'd28} : s = 2;
	{8'd100,8'd29} : s = 48;
	{8'd100,8'd30} : s = 40;
	{8'd100,8'd31} : s = 168;
	{8'd100,8'd32} : s = 36;
	{8'd100,8'd33} : s = 164;
	{8'd100,8'd34} : s = 162;
	{8'd100,8'd35} : s = 323;
	{8'd100,8'd36} : s = 34;
	{8'd100,8'd37} : s = 161;
	{8'd100,8'd38} : s = 152;
	{8'd100,8'd39} : s = 312;
	{8'd100,8'd40} : s = 148;
	{8'd100,8'd41} : s = 308;
	{8'd100,8'd42} : s = 306;
	{8'd100,8'd43} : s = 425;
	{8'd100,8'd44} : s = 33;
	{8'd100,8'd45} : s = 146;
	{8'd100,8'd46} : s = 145;
	{8'd100,8'd47} : s = 305;
	{8'd100,8'd48} : s = 140;
	{8'd100,8'd49} : s = 300;
	{8'd100,8'd50} : s = 298;
	{8'd100,8'd51} : s = 422;
	{8'd100,8'd52} : s = 138;
	{8'd100,8'd53} : s = 297;
	{8'd100,8'd54} : s = 294;
	{8'd100,8'd55} : s = 421;
	{8'd100,8'd56} : s = 293;
	{8'd100,8'd57} : s = 419;
	{8'd100,8'd58} : s = 412;
	{8'd100,8'd59} : s = 486;
	{8'd100,8'd60} : s = 24;
	{8'd100,8'd61} : s = 137;
	{8'd100,8'd62} : s = 134;
	{8'd100,8'd63} : s = 291;
	{8'd100,8'd64} : s = 133;
	{8'd100,8'd65} : s = 284;
	{8'd100,8'd66} : s = 282;
	{8'd100,8'd67} : s = 410;
	{8'd100,8'd68} : s = 131;
	{8'd100,8'd69} : s = 281;
	{8'd100,8'd70} : s = 278;
	{8'd100,8'd71} : s = 409;
	{8'd100,8'd72} : s = 277;
	{8'd100,8'd73} : s = 406;
	{8'd100,8'd74} : s = 405;
	{8'd100,8'd75} : s = 485;
	{8'd100,8'd76} : s = 112;
	{8'd100,8'd77} : s = 275;
	{8'd100,8'd78} : s = 270;
	{8'd100,8'd79} : s = 403;
	{8'd100,8'd80} : s = 269;
	{8'd100,8'd81} : s = 398;
	{8'd100,8'd82} : s = 397;
	{8'd100,8'd83} : s = 483;
	{8'd100,8'd84} : s = 267;
	{8'd100,8'd85} : s = 395;
	{8'd100,8'd86} : s = 391;
	{8'd100,8'd87} : s = 476;
	{8'd100,8'd88} : s = 376;
	{8'd100,8'd89} : s = 474;
	{8'd100,8'd90} : s = 473;
	{8'd100,8'd91} : s = 506;
	{8'd100,8'd92} : s = 20;
	{8'd100,8'd93} : s = 104;
	{8'd100,8'd94} : s = 100;
	{8'd100,8'd95} : s = 263;
	{8'd100,8'd96} : s = 98;
	{8'd100,8'd97} : s = 240;
	{8'd100,8'd98} : s = 232;
	{8'd100,8'd99} : s = 372;
	{8'd100,8'd100} : s = 97;
	{8'd100,8'd101} : s = 228;
	{8'd100,8'd102} : s = 226;
	{8'd100,8'd103} : s = 370;
	{8'd100,8'd104} : s = 225;
	{8'd100,8'd105} : s = 369;
	{8'd100,8'd106} : s = 364;
	{8'd100,8'd107} : s = 470;
	{8'd100,8'd108} : s = 88;
	{8'd100,8'd109} : s = 216;
	{8'd100,8'd110} : s = 212;
	{8'd100,8'd111} : s = 362;
	{8'd100,8'd112} : s = 210;
	{8'd100,8'd113} : s = 361;
	{8'd100,8'd114} : s = 358;
	{8'd100,8'd115} : s = 469;
	{8'd100,8'd116} : s = 209;
	{8'd100,8'd117} : s = 357;
	{8'd100,8'd118} : s = 355;
	{8'd100,8'd119} : s = 467;
	{8'd100,8'd120} : s = 348;
	{8'd100,8'd121} : s = 462;
	{8'd100,8'd122} : s = 461;
	{8'd100,8'd123} : s = 505;
	{8'd100,8'd124} : s = 84;
	{8'd100,8'd125} : s = 204;
	{8'd100,8'd126} : s = 202;
	{8'd100,8'd127} : s = 346;
	{8'd100,8'd128} : s = 201;
	{8'd100,8'd129} : s = 345;
	{8'd100,8'd130} : s = 342;
	{8'd100,8'd131} : s = 459;
	{8'd100,8'd132} : s = 198;
	{8'd100,8'd133} : s = 341;
	{8'd100,8'd134} : s = 339;
	{8'd100,8'd135} : s = 455;
	{8'd100,8'd136} : s = 334;
	{8'd100,8'd137} : s = 444;
	{8'd100,8'd138} : s = 442;
	{8'd100,8'd139} : s = 502;
	{8'd100,8'd140} : s = 197;
	{8'd100,8'd141} : s = 333;
	{8'd100,8'd142} : s = 331;
	{8'd100,8'd143} : s = 441;
	{8'd100,8'd144} : s = 327;
	{8'd100,8'd145} : s = 438;
	{8'd100,8'd146} : s = 437;
	{8'd100,8'd147} : s = 501;
	{8'd100,8'd148} : s = 316;
	{8'd100,8'd149} : s = 435;
	{8'd100,8'd150} : s = 430;
	{8'd100,8'd151} : s = 499;
	{8'd100,8'd152} : s = 429;
	{8'd100,8'd153} : s = 494;
	{8'd100,8'd154} : s = 493;
	{8'd100,8'd155} : s = 510;
	{8'd100,8'd156} : s = 1;
	{8'd100,8'd157} : s = 18;
	{8'd100,8'd158} : s = 17;
	{8'd100,8'd159} : s = 82;
	{8'd100,8'd160} : s = 12;
	{8'd100,8'd161} : s = 81;
	{8'd100,8'd162} : s = 76;
	{8'd100,8'd163} : s = 195;
	{8'd100,8'd164} : s = 10;
	{8'd100,8'd165} : s = 74;
	{8'd100,8'd166} : s = 73;
	{8'd100,8'd167} : s = 184;
	{8'd100,8'd168} : s = 70;
	{8'd100,8'd169} : s = 180;
	{8'd100,8'd170} : s = 178;
	{8'd100,8'd171} : s = 314;
	{8'd100,8'd172} : s = 9;
	{8'd100,8'd173} : s = 69;
	{8'd100,8'd174} : s = 67;
	{8'd100,8'd175} : s = 177;
	{8'd100,8'd176} : s = 56;
	{8'd100,8'd177} : s = 172;
	{8'd100,8'd178} : s = 170;
	{8'd100,8'd179} : s = 313;
	{8'd100,8'd180} : s = 52;
	{8'd100,8'd181} : s = 169;
	{8'd100,8'd182} : s = 166;
	{8'd100,8'd183} : s = 310;
	{8'd100,8'd184} : s = 165;
	{8'd100,8'd185} : s = 309;
	{8'd100,8'd186} : s = 307;
	{8'd100,8'd187} : s = 427;
	{8'd100,8'd188} : s = 6;
	{8'd100,8'd189} : s = 50;
	{8'd100,8'd190} : s = 49;
	{8'd100,8'd191} : s = 163;
	{8'd100,8'd192} : s = 44;
	{8'd100,8'd193} : s = 156;
	{8'd100,8'd194} : s = 154;
	{8'd100,8'd195} : s = 302;
	{8'd100,8'd196} : s = 42;
	{8'd100,8'd197} : s = 153;
	{8'd100,8'd198} : s = 150;
	{8'd100,8'd199} : s = 301;
	{8'd100,8'd200} : s = 149;
	{8'd100,8'd201} : s = 299;
	{8'd100,8'd202} : s = 295;
	{8'd100,8'd203} : s = 423;
	{8'd100,8'd204} : s = 41;
	{8'd100,8'd205} : s = 147;
	{8'd100,8'd206} : s = 142;
	{8'd100,8'd207} : s = 286;
	{8'd100,8'd208} : s = 141;
	{8'd100,8'd209} : s = 285;
	{8'd100,8'd210} : s = 283;
	{8'd100,8'd211} : s = 414;
	{8'd100,8'd212} : s = 139;
	{8'd100,8'd213} : s = 279;
	{8'd100,8'd214} : s = 271;
	{8'd100,8'd215} : s = 413;
	{8'd100,8'd216} : s = 248;
	{8'd100,8'd217} : s = 411;
	{8'd100,8'd218} : s = 407;
	{8'd100,8'd219} : s = 491;
	{8'd100,8'd220} : s = 5;
	{8'd100,8'd221} : s = 38;
	{8'd100,8'd222} : s = 37;
	{8'd100,8'd223} : s = 135;
	{8'd100,8'd224} : s = 35;
	{8'd100,8'd225} : s = 120;
	{8'd100,8'd226} : s = 116;
	{8'd100,8'd227} : s = 244;
	{8'd100,8'd228} : s = 28;
	{8'd100,8'd229} : s = 114;
	{8'd100,8'd230} : s = 113;
	{8'd100,8'd231} : s = 242;
	{8'd100,8'd232} : s = 108;
	{8'd100,8'd233} : s = 241;
	{8'd100,8'd234} : s = 236;
	{8'd100,8'd235} : s = 399;
	{8'd100,8'd236} : s = 26;
	{8'd100,8'd237} : s = 106;
	{8'd100,8'd238} : s = 105;
	{8'd100,8'd239} : s = 234;
	{8'd100,8'd240} : s = 102;
	{8'd100,8'd241} : s = 233;
	{8'd100,8'd242} : s = 230;
	{8'd100,8'd243} : s = 380;
	{8'd100,8'd244} : s = 101;
	{8'd100,8'd245} : s = 229;
	{8'd100,8'd246} : s = 227;
	{8'd100,8'd247} : s = 378;
	{8'd100,8'd248} : s = 220;
	{8'd100,8'd249} : s = 377;
	{8'd100,8'd250} : s = 374;
	{8'd100,8'd251} : s = 487;
	{8'd100,8'd252} : s = 25;
	{8'd100,8'd253} : s = 99;
	{8'd100,8'd254} : s = 92;
	{8'd100,8'd255} : s = 218;
	{8'd101,8'd0} : s = 344;
	{8'd101,8'd1} : s = 340;
	{8'd101,8'd2} : s = 457;
	{8'd101,8'd3} : s = 193;
	{8'd101,8'd4} : s = 338;
	{8'd101,8'd5} : s = 337;
	{8'd101,8'd6} : s = 454;
	{8'd101,8'd7} : s = 332;
	{8'd101,8'd8} : s = 453;
	{8'd101,8'd9} : s = 451;
	{8'd101,8'd10} : s = 498;
	{8'd101,8'd11} : s = 176;
	{8'd101,8'd12} : s = 330;
	{8'd101,8'd13} : s = 329;
	{8'd101,8'd14} : s = 440;
	{8'd101,8'd15} : s = 326;
	{8'd101,8'd16} : s = 436;
	{8'd101,8'd17} : s = 434;
	{8'd101,8'd18} : s = 497;
	{8'd101,8'd19} : s = 325;
	{8'd101,8'd20} : s = 433;
	{8'd101,8'd21} : s = 428;
	{8'd101,8'd22} : s = 492;
	{8'd101,8'd23} : s = 426;
	{8'd101,8'd24} : s = 490;
	{8'd101,8'd25} : s = 489;
	{8'd101,8'd26} : s = 508;
	{8'd101,8'd27} : s = 2;
	{8'd101,8'd28} : s = 48;
	{8'd101,8'd29} : s = 40;
	{8'd101,8'd30} : s = 168;
	{8'd101,8'd31} : s = 36;
	{8'd101,8'd32} : s = 164;
	{8'd101,8'd33} : s = 162;
	{8'd101,8'd34} : s = 323;
	{8'd101,8'd35} : s = 34;
	{8'd101,8'd36} : s = 161;
	{8'd101,8'd37} : s = 152;
	{8'd101,8'd38} : s = 312;
	{8'd101,8'd39} : s = 148;
	{8'd101,8'd40} : s = 308;
	{8'd101,8'd41} : s = 306;
	{8'd101,8'd42} : s = 425;
	{8'd101,8'd43} : s = 33;
	{8'd101,8'd44} : s = 146;
	{8'd101,8'd45} : s = 145;
	{8'd101,8'd46} : s = 305;
	{8'd101,8'd47} : s = 140;
	{8'd101,8'd48} : s = 300;
	{8'd101,8'd49} : s = 298;
	{8'd101,8'd50} : s = 422;
	{8'd101,8'd51} : s = 138;
	{8'd101,8'd52} : s = 297;
	{8'd101,8'd53} : s = 294;
	{8'd101,8'd54} : s = 421;
	{8'd101,8'd55} : s = 293;
	{8'd101,8'd56} : s = 419;
	{8'd101,8'd57} : s = 412;
	{8'd101,8'd58} : s = 486;
	{8'd101,8'd59} : s = 24;
	{8'd101,8'd60} : s = 137;
	{8'd101,8'd61} : s = 134;
	{8'd101,8'd62} : s = 291;
	{8'd101,8'd63} : s = 133;
	{8'd101,8'd64} : s = 284;
	{8'd101,8'd65} : s = 282;
	{8'd101,8'd66} : s = 410;
	{8'd101,8'd67} : s = 131;
	{8'd101,8'd68} : s = 281;
	{8'd101,8'd69} : s = 278;
	{8'd101,8'd70} : s = 409;
	{8'd101,8'd71} : s = 277;
	{8'd101,8'd72} : s = 406;
	{8'd101,8'd73} : s = 405;
	{8'd101,8'd74} : s = 485;
	{8'd101,8'd75} : s = 112;
	{8'd101,8'd76} : s = 275;
	{8'd101,8'd77} : s = 270;
	{8'd101,8'd78} : s = 403;
	{8'd101,8'd79} : s = 269;
	{8'd101,8'd80} : s = 398;
	{8'd101,8'd81} : s = 397;
	{8'd101,8'd82} : s = 483;
	{8'd101,8'd83} : s = 267;
	{8'd101,8'd84} : s = 395;
	{8'd101,8'd85} : s = 391;
	{8'd101,8'd86} : s = 476;
	{8'd101,8'd87} : s = 376;
	{8'd101,8'd88} : s = 474;
	{8'd101,8'd89} : s = 473;
	{8'd101,8'd90} : s = 506;
	{8'd101,8'd91} : s = 20;
	{8'd101,8'd92} : s = 104;
	{8'd101,8'd93} : s = 100;
	{8'd101,8'd94} : s = 263;
	{8'd101,8'd95} : s = 98;
	{8'd101,8'd96} : s = 240;
	{8'd101,8'd97} : s = 232;
	{8'd101,8'd98} : s = 372;
	{8'd101,8'd99} : s = 97;
	{8'd101,8'd100} : s = 228;
	{8'd101,8'd101} : s = 226;
	{8'd101,8'd102} : s = 370;
	{8'd101,8'd103} : s = 225;
	{8'd101,8'd104} : s = 369;
	{8'd101,8'd105} : s = 364;
	{8'd101,8'd106} : s = 470;
	{8'd101,8'd107} : s = 88;
	{8'd101,8'd108} : s = 216;
	{8'd101,8'd109} : s = 212;
	{8'd101,8'd110} : s = 362;
	{8'd101,8'd111} : s = 210;
	{8'd101,8'd112} : s = 361;
	{8'd101,8'd113} : s = 358;
	{8'd101,8'd114} : s = 469;
	{8'd101,8'd115} : s = 209;
	{8'd101,8'd116} : s = 357;
	{8'd101,8'd117} : s = 355;
	{8'd101,8'd118} : s = 467;
	{8'd101,8'd119} : s = 348;
	{8'd101,8'd120} : s = 462;
	{8'd101,8'd121} : s = 461;
	{8'd101,8'd122} : s = 505;
	{8'd101,8'd123} : s = 84;
	{8'd101,8'd124} : s = 204;
	{8'd101,8'd125} : s = 202;
	{8'd101,8'd126} : s = 346;
	{8'd101,8'd127} : s = 201;
	{8'd101,8'd128} : s = 345;
	{8'd101,8'd129} : s = 342;
	{8'd101,8'd130} : s = 459;
	{8'd101,8'd131} : s = 198;
	{8'd101,8'd132} : s = 341;
	{8'd101,8'd133} : s = 339;
	{8'd101,8'd134} : s = 455;
	{8'd101,8'd135} : s = 334;
	{8'd101,8'd136} : s = 444;
	{8'd101,8'd137} : s = 442;
	{8'd101,8'd138} : s = 502;
	{8'd101,8'd139} : s = 197;
	{8'd101,8'd140} : s = 333;
	{8'd101,8'd141} : s = 331;
	{8'd101,8'd142} : s = 441;
	{8'd101,8'd143} : s = 327;
	{8'd101,8'd144} : s = 438;
	{8'd101,8'd145} : s = 437;
	{8'd101,8'd146} : s = 501;
	{8'd101,8'd147} : s = 316;
	{8'd101,8'd148} : s = 435;
	{8'd101,8'd149} : s = 430;
	{8'd101,8'd150} : s = 499;
	{8'd101,8'd151} : s = 429;
	{8'd101,8'd152} : s = 494;
	{8'd101,8'd153} : s = 493;
	{8'd101,8'd154} : s = 510;
	{8'd101,8'd155} : s = 1;
	{8'd101,8'd156} : s = 18;
	{8'd101,8'd157} : s = 17;
	{8'd101,8'd158} : s = 82;
	{8'd101,8'd159} : s = 12;
	{8'd101,8'd160} : s = 81;
	{8'd101,8'd161} : s = 76;
	{8'd101,8'd162} : s = 195;
	{8'd101,8'd163} : s = 10;
	{8'd101,8'd164} : s = 74;
	{8'd101,8'd165} : s = 73;
	{8'd101,8'd166} : s = 184;
	{8'd101,8'd167} : s = 70;
	{8'd101,8'd168} : s = 180;
	{8'd101,8'd169} : s = 178;
	{8'd101,8'd170} : s = 314;
	{8'd101,8'd171} : s = 9;
	{8'd101,8'd172} : s = 69;
	{8'd101,8'd173} : s = 67;
	{8'd101,8'd174} : s = 177;
	{8'd101,8'd175} : s = 56;
	{8'd101,8'd176} : s = 172;
	{8'd101,8'd177} : s = 170;
	{8'd101,8'd178} : s = 313;
	{8'd101,8'd179} : s = 52;
	{8'd101,8'd180} : s = 169;
	{8'd101,8'd181} : s = 166;
	{8'd101,8'd182} : s = 310;
	{8'd101,8'd183} : s = 165;
	{8'd101,8'd184} : s = 309;
	{8'd101,8'd185} : s = 307;
	{8'd101,8'd186} : s = 427;
	{8'd101,8'd187} : s = 6;
	{8'd101,8'd188} : s = 50;
	{8'd101,8'd189} : s = 49;
	{8'd101,8'd190} : s = 163;
	{8'd101,8'd191} : s = 44;
	{8'd101,8'd192} : s = 156;
	{8'd101,8'd193} : s = 154;
	{8'd101,8'd194} : s = 302;
	{8'd101,8'd195} : s = 42;
	{8'd101,8'd196} : s = 153;
	{8'd101,8'd197} : s = 150;
	{8'd101,8'd198} : s = 301;
	{8'd101,8'd199} : s = 149;
	{8'd101,8'd200} : s = 299;
	{8'd101,8'd201} : s = 295;
	{8'd101,8'd202} : s = 423;
	{8'd101,8'd203} : s = 41;
	{8'd101,8'd204} : s = 147;
	{8'd101,8'd205} : s = 142;
	{8'd101,8'd206} : s = 286;
	{8'd101,8'd207} : s = 141;
	{8'd101,8'd208} : s = 285;
	{8'd101,8'd209} : s = 283;
	{8'd101,8'd210} : s = 414;
	{8'd101,8'd211} : s = 139;
	{8'd101,8'd212} : s = 279;
	{8'd101,8'd213} : s = 271;
	{8'd101,8'd214} : s = 413;
	{8'd101,8'd215} : s = 248;
	{8'd101,8'd216} : s = 411;
	{8'd101,8'd217} : s = 407;
	{8'd101,8'd218} : s = 491;
	{8'd101,8'd219} : s = 5;
	{8'd101,8'd220} : s = 38;
	{8'd101,8'd221} : s = 37;
	{8'd101,8'd222} : s = 135;
	{8'd101,8'd223} : s = 35;
	{8'd101,8'd224} : s = 120;
	{8'd101,8'd225} : s = 116;
	{8'd101,8'd226} : s = 244;
	{8'd101,8'd227} : s = 28;
	{8'd101,8'd228} : s = 114;
	{8'd101,8'd229} : s = 113;
	{8'd101,8'd230} : s = 242;
	{8'd101,8'd231} : s = 108;
	{8'd101,8'd232} : s = 241;
	{8'd101,8'd233} : s = 236;
	{8'd101,8'd234} : s = 399;
	{8'd101,8'd235} : s = 26;
	{8'd101,8'd236} : s = 106;
	{8'd101,8'd237} : s = 105;
	{8'd101,8'd238} : s = 234;
	{8'd101,8'd239} : s = 102;
	{8'd101,8'd240} : s = 233;
	{8'd101,8'd241} : s = 230;
	{8'd101,8'd242} : s = 380;
	{8'd101,8'd243} : s = 101;
	{8'd101,8'd244} : s = 229;
	{8'd101,8'd245} : s = 227;
	{8'd101,8'd246} : s = 378;
	{8'd101,8'd247} : s = 220;
	{8'd101,8'd248} : s = 377;
	{8'd101,8'd249} : s = 374;
	{8'd101,8'd250} : s = 487;
	{8'd101,8'd251} : s = 25;
	{8'd101,8'd252} : s = 99;
	{8'd101,8'd253} : s = 92;
	{8'd101,8'd254} : s = 218;
	{8'd101,8'd255} : s = 90;
	{8'd102,8'd0} : s = 340;
	{8'd102,8'd1} : s = 457;
	{8'd102,8'd2} : s = 193;
	{8'd102,8'd3} : s = 338;
	{8'd102,8'd4} : s = 337;
	{8'd102,8'd5} : s = 454;
	{8'd102,8'd6} : s = 332;
	{8'd102,8'd7} : s = 453;
	{8'd102,8'd8} : s = 451;
	{8'd102,8'd9} : s = 498;
	{8'd102,8'd10} : s = 176;
	{8'd102,8'd11} : s = 330;
	{8'd102,8'd12} : s = 329;
	{8'd102,8'd13} : s = 440;
	{8'd102,8'd14} : s = 326;
	{8'd102,8'd15} : s = 436;
	{8'd102,8'd16} : s = 434;
	{8'd102,8'd17} : s = 497;
	{8'd102,8'd18} : s = 325;
	{8'd102,8'd19} : s = 433;
	{8'd102,8'd20} : s = 428;
	{8'd102,8'd21} : s = 492;
	{8'd102,8'd22} : s = 426;
	{8'd102,8'd23} : s = 490;
	{8'd102,8'd24} : s = 489;
	{8'd102,8'd25} : s = 508;
	{8'd102,8'd26} : s = 2;
	{8'd102,8'd27} : s = 48;
	{8'd102,8'd28} : s = 40;
	{8'd102,8'd29} : s = 168;
	{8'd102,8'd30} : s = 36;
	{8'd102,8'd31} : s = 164;
	{8'd102,8'd32} : s = 162;
	{8'd102,8'd33} : s = 323;
	{8'd102,8'd34} : s = 34;
	{8'd102,8'd35} : s = 161;
	{8'd102,8'd36} : s = 152;
	{8'd102,8'd37} : s = 312;
	{8'd102,8'd38} : s = 148;
	{8'd102,8'd39} : s = 308;
	{8'd102,8'd40} : s = 306;
	{8'd102,8'd41} : s = 425;
	{8'd102,8'd42} : s = 33;
	{8'd102,8'd43} : s = 146;
	{8'd102,8'd44} : s = 145;
	{8'd102,8'd45} : s = 305;
	{8'd102,8'd46} : s = 140;
	{8'd102,8'd47} : s = 300;
	{8'd102,8'd48} : s = 298;
	{8'd102,8'd49} : s = 422;
	{8'd102,8'd50} : s = 138;
	{8'd102,8'd51} : s = 297;
	{8'd102,8'd52} : s = 294;
	{8'd102,8'd53} : s = 421;
	{8'd102,8'd54} : s = 293;
	{8'd102,8'd55} : s = 419;
	{8'd102,8'd56} : s = 412;
	{8'd102,8'd57} : s = 486;
	{8'd102,8'd58} : s = 24;
	{8'd102,8'd59} : s = 137;
	{8'd102,8'd60} : s = 134;
	{8'd102,8'd61} : s = 291;
	{8'd102,8'd62} : s = 133;
	{8'd102,8'd63} : s = 284;
	{8'd102,8'd64} : s = 282;
	{8'd102,8'd65} : s = 410;
	{8'd102,8'd66} : s = 131;
	{8'd102,8'd67} : s = 281;
	{8'd102,8'd68} : s = 278;
	{8'd102,8'd69} : s = 409;
	{8'd102,8'd70} : s = 277;
	{8'd102,8'd71} : s = 406;
	{8'd102,8'd72} : s = 405;
	{8'd102,8'd73} : s = 485;
	{8'd102,8'd74} : s = 112;
	{8'd102,8'd75} : s = 275;
	{8'd102,8'd76} : s = 270;
	{8'd102,8'd77} : s = 403;
	{8'd102,8'd78} : s = 269;
	{8'd102,8'd79} : s = 398;
	{8'd102,8'd80} : s = 397;
	{8'd102,8'd81} : s = 483;
	{8'd102,8'd82} : s = 267;
	{8'd102,8'd83} : s = 395;
	{8'd102,8'd84} : s = 391;
	{8'd102,8'd85} : s = 476;
	{8'd102,8'd86} : s = 376;
	{8'd102,8'd87} : s = 474;
	{8'd102,8'd88} : s = 473;
	{8'd102,8'd89} : s = 506;
	{8'd102,8'd90} : s = 20;
	{8'd102,8'd91} : s = 104;
	{8'd102,8'd92} : s = 100;
	{8'd102,8'd93} : s = 263;
	{8'd102,8'd94} : s = 98;
	{8'd102,8'd95} : s = 240;
	{8'd102,8'd96} : s = 232;
	{8'd102,8'd97} : s = 372;
	{8'd102,8'd98} : s = 97;
	{8'd102,8'd99} : s = 228;
	{8'd102,8'd100} : s = 226;
	{8'd102,8'd101} : s = 370;
	{8'd102,8'd102} : s = 225;
	{8'd102,8'd103} : s = 369;
	{8'd102,8'd104} : s = 364;
	{8'd102,8'd105} : s = 470;
	{8'd102,8'd106} : s = 88;
	{8'd102,8'd107} : s = 216;
	{8'd102,8'd108} : s = 212;
	{8'd102,8'd109} : s = 362;
	{8'd102,8'd110} : s = 210;
	{8'd102,8'd111} : s = 361;
	{8'd102,8'd112} : s = 358;
	{8'd102,8'd113} : s = 469;
	{8'd102,8'd114} : s = 209;
	{8'd102,8'd115} : s = 357;
	{8'd102,8'd116} : s = 355;
	{8'd102,8'd117} : s = 467;
	{8'd102,8'd118} : s = 348;
	{8'd102,8'd119} : s = 462;
	{8'd102,8'd120} : s = 461;
	{8'd102,8'd121} : s = 505;
	{8'd102,8'd122} : s = 84;
	{8'd102,8'd123} : s = 204;
	{8'd102,8'd124} : s = 202;
	{8'd102,8'd125} : s = 346;
	{8'd102,8'd126} : s = 201;
	{8'd102,8'd127} : s = 345;
	{8'd102,8'd128} : s = 342;
	{8'd102,8'd129} : s = 459;
	{8'd102,8'd130} : s = 198;
	{8'd102,8'd131} : s = 341;
	{8'd102,8'd132} : s = 339;
	{8'd102,8'd133} : s = 455;
	{8'd102,8'd134} : s = 334;
	{8'd102,8'd135} : s = 444;
	{8'd102,8'd136} : s = 442;
	{8'd102,8'd137} : s = 502;
	{8'd102,8'd138} : s = 197;
	{8'd102,8'd139} : s = 333;
	{8'd102,8'd140} : s = 331;
	{8'd102,8'd141} : s = 441;
	{8'd102,8'd142} : s = 327;
	{8'd102,8'd143} : s = 438;
	{8'd102,8'd144} : s = 437;
	{8'd102,8'd145} : s = 501;
	{8'd102,8'd146} : s = 316;
	{8'd102,8'd147} : s = 435;
	{8'd102,8'd148} : s = 430;
	{8'd102,8'd149} : s = 499;
	{8'd102,8'd150} : s = 429;
	{8'd102,8'd151} : s = 494;
	{8'd102,8'd152} : s = 493;
	{8'd102,8'd153} : s = 510;
	{8'd102,8'd154} : s = 1;
	{8'd102,8'd155} : s = 18;
	{8'd102,8'd156} : s = 17;
	{8'd102,8'd157} : s = 82;
	{8'd102,8'd158} : s = 12;
	{8'd102,8'd159} : s = 81;
	{8'd102,8'd160} : s = 76;
	{8'd102,8'd161} : s = 195;
	{8'd102,8'd162} : s = 10;
	{8'd102,8'd163} : s = 74;
	{8'd102,8'd164} : s = 73;
	{8'd102,8'd165} : s = 184;
	{8'd102,8'd166} : s = 70;
	{8'd102,8'd167} : s = 180;
	{8'd102,8'd168} : s = 178;
	{8'd102,8'd169} : s = 314;
	{8'd102,8'd170} : s = 9;
	{8'd102,8'd171} : s = 69;
	{8'd102,8'd172} : s = 67;
	{8'd102,8'd173} : s = 177;
	{8'd102,8'd174} : s = 56;
	{8'd102,8'd175} : s = 172;
	{8'd102,8'd176} : s = 170;
	{8'd102,8'd177} : s = 313;
	{8'd102,8'd178} : s = 52;
	{8'd102,8'd179} : s = 169;
	{8'd102,8'd180} : s = 166;
	{8'd102,8'd181} : s = 310;
	{8'd102,8'd182} : s = 165;
	{8'd102,8'd183} : s = 309;
	{8'd102,8'd184} : s = 307;
	{8'd102,8'd185} : s = 427;
	{8'd102,8'd186} : s = 6;
	{8'd102,8'd187} : s = 50;
	{8'd102,8'd188} : s = 49;
	{8'd102,8'd189} : s = 163;
	{8'd102,8'd190} : s = 44;
	{8'd102,8'd191} : s = 156;
	{8'd102,8'd192} : s = 154;
	{8'd102,8'd193} : s = 302;
	{8'd102,8'd194} : s = 42;
	{8'd102,8'd195} : s = 153;
	{8'd102,8'd196} : s = 150;
	{8'd102,8'd197} : s = 301;
	{8'd102,8'd198} : s = 149;
	{8'd102,8'd199} : s = 299;
	{8'd102,8'd200} : s = 295;
	{8'd102,8'd201} : s = 423;
	{8'd102,8'd202} : s = 41;
	{8'd102,8'd203} : s = 147;
	{8'd102,8'd204} : s = 142;
	{8'd102,8'd205} : s = 286;
	{8'd102,8'd206} : s = 141;
	{8'd102,8'd207} : s = 285;
	{8'd102,8'd208} : s = 283;
	{8'd102,8'd209} : s = 414;
	{8'd102,8'd210} : s = 139;
	{8'd102,8'd211} : s = 279;
	{8'd102,8'd212} : s = 271;
	{8'd102,8'd213} : s = 413;
	{8'd102,8'd214} : s = 248;
	{8'd102,8'd215} : s = 411;
	{8'd102,8'd216} : s = 407;
	{8'd102,8'd217} : s = 491;
	{8'd102,8'd218} : s = 5;
	{8'd102,8'd219} : s = 38;
	{8'd102,8'd220} : s = 37;
	{8'd102,8'd221} : s = 135;
	{8'd102,8'd222} : s = 35;
	{8'd102,8'd223} : s = 120;
	{8'd102,8'd224} : s = 116;
	{8'd102,8'd225} : s = 244;
	{8'd102,8'd226} : s = 28;
	{8'd102,8'd227} : s = 114;
	{8'd102,8'd228} : s = 113;
	{8'd102,8'd229} : s = 242;
	{8'd102,8'd230} : s = 108;
	{8'd102,8'd231} : s = 241;
	{8'd102,8'd232} : s = 236;
	{8'd102,8'd233} : s = 399;
	{8'd102,8'd234} : s = 26;
	{8'd102,8'd235} : s = 106;
	{8'd102,8'd236} : s = 105;
	{8'd102,8'd237} : s = 234;
	{8'd102,8'd238} : s = 102;
	{8'd102,8'd239} : s = 233;
	{8'd102,8'd240} : s = 230;
	{8'd102,8'd241} : s = 380;
	{8'd102,8'd242} : s = 101;
	{8'd102,8'd243} : s = 229;
	{8'd102,8'd244} : s = 227;
	{8'd102,8'd245} : s = 378;
	{8'd102,8'd246} : s = 220;
	{8'd102,8'd247} : s = 377;
	{8'd102,8'd248} : s = 374;
	{8'd102,8'd249} : s = 487;
	{8'd102,8'd250} : s = 25;
	{8'd102,8'd251} : s = 99;
	{8'd102,8'd252} : s = 92;
	{8'd102,8'd253} : s = 218;
	{8'd102,8'd254} : s = 90;
	{8'd102,8'd255} : s = 217;
	{8'd103,8'd0} : s = 457;
	{8'd103,8'd1} : s = 193;
	{8'd103,8'd2} : s = 338;
	{8'd103,8'd3} : s = 337;
	{8'd103,8'd4} : s = 454;
	{8'd103,8'd5} : s = 332;
	{8'd103,8'd6} : s = 453;
	{8'd103,8'd7} : s = 451;
	{8'd103,8'd8} : s = 498;
	{8'd103,8'd9} : s = 176;
	{8'd103,8'd10} : s = 330;
	{8'd103,8'd11} : s = 329;
	{8'd103,8'd12} : s = 440;
	{8'd103,8'd13} : s = 326;
	{8'd103,8'd14} : s = 436;
	{8'd103,8'd15} : s = 434;
	{8'd103,8'd16} : s = 497;
	{8'd103,8'd17} : s = 325;
	{8'd103,8'd18} : s = 433;
	{8'd103,8'd19} : s = 428;
	{8'd103,8'd20} : s = 492;
	{8'd103,8'd21} : s = 426;
	{8'd103,8'd22} : s = 490;
	{8'd103,8'd23} : s = 489;
	{8'd103,8'd24} : s = 508;
	{8'd103,8'd25} : s = 2;
	{8'd103,8'd26} : s = 48;
	{8'd103,8'd27} : s = 40;
	{8'd103,8'd28} : s = 168;
	{8'd103,8'd29} : s = 36;
	{8'd103,8'd30} : s = 164;
	{8'd103,8'd31} : s = 162;
	{8'd103,8'd32} : s = 323;
	{8'd103,8'd33} : s = 34;
	{8'd103,8'd34} : s = 161;
	{8'd103,8'd35} : s = 152;
	{8'd103,8'd36} : s = 312;
	{8'd103,8'd37} : s = 148;
	{8'd103,8'd38} : s = 308;
	{8'd103,8'd39} : s = 306;
	{8'd103,8'd40} : s = 425;
	{8'd103,8'd41} : s = 33;
	{8'd103,8'd42} : s = 146;
	{8'd103,8'd43} : s = 145;
	{8'd103,8'd44} : s = 305;
	{8'd103,8'd45} : s = 140;
	{8'd103,8'd46} : s = 300;
	{8'd103,8'd47} : s = 298;
	{8'd103,8'd48} : s = 422;
	{8'd103,8'd49} : s = 138;
	{8'd103,8'd50} : s = 297;
	{8'd103,8'd51} : s = 294;
	{8'd103,8'd52} : s = 421;
	{8'd103,8'd53} : s = 293;
	{8'd103,8'd54} : s = 419;
	{8'd103,8'd55} : s = 412;
	{8'd103,8'd56} : s = 486;
	{8'd103,8'd57} : s = 24;
	{8'd103,8'd58} : s = 137;
	{8'd103,8'd59} : s = 134;
	{8'd103,8'd60} : s = 291;
	{8'd103,8'd61} : s = 133;
	{8'd103,8'd62} : s = 284;
	{8'd103,8'd63} : s = 282;
	{8'd103,8'd64} : s = 410;
	{8'd103,8'd65} : s = 131;
	{8'd103,8'd66} : s = 281;
	{8'd103,8'd67} : s = 278;
	{8'd103,8'd68} : s = 409;
	{8'd103,8'd69} : s = 277;
	{8'd103,8'd70} : s = 406;
	{8'd103,8'd71} : s = 405;
	{8'd103,8'd72} : s = 485;
	{8'd103,8'd73} : s = 112;
	{8'd103,8'd74} : s = 275;
	{8'd103,8'd75} : s = 270;
	{8'd103,8'd76} : s = 403;
	{8'd103,8'd77} : s = 269;
	{8'd103,8'd78} : s = 398;
	{8'd103,8'd79} : s = 397;
	{8'd103,8'd80} : s = 483;
	{8'd103,8'd81} : s = 267;
	{8'd103,8'd82} : s = 395;
	{8'd103,8'd83} : s = 391;
	{8'd103,8'd84} : s = 476;
	{8'd103,8'd85} : s = 376;
	{8'd103,8'd86} : s = 474;
	{8'd103,8'd87} : s = 473;
	{8'd103,8'd88} : s = 506;
	{8'd103,8'd89} : s = 20;
	{8'd103,8'd90} : s = 104;
	{8'd103,8'd91} : s = 100;
	{8'd103,8'd92} : s = 263;
	{8'd103,8'd93} : s = 98;
	{8'd103,8'd94} : s = 240;
	{8'd103,8'd95} : s = 232;
	{8'd103,8'd96} : s = 372;
	{8'd103,8'd97} : s = 97;
	{8'd103,8'd98} : s = 228;
	{8'd103,8'd99} : s = 226;
	{8'd103,8'd100} : s = 370;
	{8'd103,8'd101} : s = 225;
	{8'd103,8'd102} : s = 369;
	{8'd103,8'd103} : s = 364;
	{8'd103,8'd104} : s = 470;
	{8'd103,8'd105} : s = 88;
	{8'd103,8'd106} : s = 216;
	{8'd103,8'd107} : s = 212;
	{8'd103,8'd108} : s = 362;
	{8'd103,8'd109} : s = 210;
	{8'd103,8'd110} : s = 361;
	{8'd103,8'd111} : s = 358;
	{8'd103,8'd112} : s = 469;
	{8'd103,8'd113} : s = 209;
	{8'd103,8'd114} : s = 357;
	{8'd103,8'd115} : s = 355;
	{8'd103,8'd116} : s = 467;
	{8'd103,8'd117} : s = 348;
	{8'd103,8'd118} : s = 462;
	{8'd103,8'd119} : s = 461;
	{8'd103,8'd120} : s = 505;
	{8'd103,8'd121} : s = 84;
	{8'd103,8'd122} : s = 204;
	{8'd103,8'd123} : s = 202;
	{8'd103,8'd124} : s = 346;
	{8'd103,8'd125} : s = 201;
	{8'd103,8'd126} : s = 345;
	{8'd103,8'd127} : s = 342;
	{8'd103,8'd128} : s = 459;
	{8'd103,8'd129} : s = 198;
	{8'd103,8'd130} : s = 341;
	{8'd103,8'd131} : s = 339;
	{8'd103,8'd132} : s = 455;
	{8'd103,8'd133} : s = 334;
	{8'd103,8'd134} : s = 444;
	{8'd103,8'd135} : s = 442;
	{8'd103,8'd136} : s = 502;
	{8'd103,8'd137} : s = 197;
	{8'd103,8'd138} : s = 333;
	{8'd103,8'd139} : s = 331;
	{8'd103,8'd140} : s = 441;
	{8'd103,8'd141} : s = 327;
	{8'd103,8'd142} : s = 438;
	{8'd103,8'd143} : s = 437;
	{8'd103,8'd144} : s = 501;
	{8'd103,8'd145} : s = 316;
	{8'd103,8'd146} : s = 435;
	{8'd103,8'd147} : s = 430;
	{8'd103,8'd148} : s = 499;
	{8'd103,8'd149} : s = 429;
	{8'd103,8'd150} : s = 494;
	{8'd103,8'd151} : s = 493;
	{8'd103,8'd152} : s = 510;
	{8'd103,8'd153} : s = 1;
	{8'd103,8'd154} : s = 18;
	{8'd103,8'd155} : s = 17;
	{8'd103,8'd156} : s = 82;
	{8'd103,8'd157} : s = 12;
	{8'd103,8'd158} : s = 81;
	{8'd103,8'd159} : s = 76;
	{8'd103,8'd160} : s = 195;
	{8'd103,8'd161} : s = 10;
	{8'd103,8'd162} : s = 74;
	{8'd103,8'd163} : s = 73;
	{8'd103,8'd164} : s = 184;
	{8'd103,8'd165} : s = 70;
	{8'd103,8'd166} : s = 180;
	{8'd103,8'd167} : s = 178;
	{8'd103,8'd168} : s = 314;
	{8'd103,8'd169} : s = 9;
	{8'd103,8'd170} : s = 69;
	{8'd103,8'd171} : s = 67;
	{8'd103,8'd172} : s = 177;
	{8'd103,8'd173} : s = 56;
	{8'd103,8'd174} : s = 172;
	{8'd103,8'd175} : s = 170;
	{8'd103,8'd176} : s = 313;
	{8'd103,8'd177} : s = 52;
	{8'd103,8'd178} : s = 169;
	{8'd103,8'd179} : s = 166;
	{8'd103,8'd180} : s = 310;
	{8'd103,8'd181} : s = 165;
	{8'd103,8'd182} : s = 309;
	{8'd103,8'd183} : s = 307;
	{8'd103,8'd184} : s = 427;
	{8'd103,8'd185} : s = 6;
	{8'd103,8'd186} : s = 50;
	{8'd103,8'd187} : s = 49;
	{8'd103,8'd188} : s = 163;
	{8'd103,8'd189} : s = 44;
	{8'd103,8'd190} : s = 156;
	{8'd103,8'd191} : s = 154;
	{8'd103,8'd192} : s = 302;
	{8'd103,8'd193} : s = 42;
	{8'd103,8'd194} : s = 153;
	{8'd103,8'd195} : s = 150;
	{8'd103,8'd196} : s = 301;
	{8'd103,8'd197} : s = 149;
	{8'd103,8'd198} : s = 299;
	{8'd103,8'd199} : s = 295;
	{8'd103,8'd200} : s = 423;
	{8'd103,8'd201} : s = 41;
	{8'd103,8'd202} : s = 147;
	{8'd103,8'd203} : s = 142;
	{8'd103,8'd204} : s = 286;
	{8'd103,8'd205} : s = 141;
	{8'd103,8'd206} : s = 285;
	{8'd103,8'd207} : s = 283;
	{8'd103,8'd208} : s = 414;
	{8'd103,8'd209} : s = 139;
	{8'd103,8'd210} : s = 279;
	{8'd103,8'd211} : s = 271;
	{8'd103,8'd212} : s = 413;
	{8'd103,8'd213} : s = 248;
	{8'd103,8'd214} : s = 411;
	{8'd103,8'd215} : s = 407;
	{8'd103,8'd216} : s = 491;
	{8'd103,8'd217} : s = 5;
	{8'd103,8'd218} : s = 38;
	{8'd103,8'd219} : s = 37;
	{8'd103,8'd220} : s = 135;
	{8'd103,8'd221} : s = 35;
	{8'd103,8'd222} : s = 120;
	{8'd103,8'd223} : s = 116;
	{8'd103,8'd224} : s = 244;
	{8'd103,8'd225} : s = 28;
	{8'd103,8'd226} : s = 114;
	{8'd103,8'd227} : s = 113;
	{8'd103,8'd228} : s = 242;
	{8'd103,8'd229} : s = 108;
	{8'd103,8'd230} : s = 241;
	{8'd103,8'd231} : s = 236;
	{8'd103,8'd232} : s = 399;
	{8'd103,8'd233} : s = 26;
	{8'd103,8'd234} : s = 106;
	{8'd103,8'd235} : s = 105;
	{8'd103,8'd236} : s = 234;
	{8'd103,8'd237} : s = 102;
	{8'd103,8'd238} : s = 233;
	{8'd103,8'd239} : s = 230;
	{8'd103,8'd240} : s = 380;
	{8'd103,8'd241} : s = 101;
	{8'd103,8'd242} : s = 229;
	{8'd103,8'd243} : s = 227;
	{8'd103,8'd244} : s = 378;
	{8'd103,8'd245} : s = 220;
	{8'd103,8'd246} : s = 377;
	{8'd103,8'd247} : s = 374;
	{8'd103,8'd248} : s = 487;
	{8'd103,8'd249} : s = 25;
	{8'd103,8'd250} : s = 99;
	{8'd103,8'd251} : s = 92;
	{8'd103,8'd252} : s = 218;
	{8'd103,8'd253} : s = 90;
	{8'd103,8'd254} : s = 217;
	{8'd103,8'd255} : s = 214;
	{8'd104,8'd0} : s = 193;
	{8'd104,8'd1} : s = 338;
	{8'd104,8'd2} : s = 337;
	{8'd104,8'd3} : s = 454;
	{8'd104,8'd4} : s = 332;
	{8'd104,8'd5} : s = 453;
	{8'd104,8'd6} : s = 451;
	{8'd104,8'd7} : s = 498;
	{8'd104,8'd8} : s = 176;
	{8'd104,8'd9} : s = 330;
	{8'd104,8'd10} : s = 329;
	{8'd104,8'd11} : s = 440;
	{8'd104,8'd12} : s = 326;
	{8'd104,8'd13} : s = 436;
	{8'd104,8'd14} : s = 434;
	{8'd104,8'd15} : s = 497;
	{8'd104,8'd16} : s = 325;
	{8'd104,8'd17} : s = 433;
	{8'd104,8'd18} : s = 428;
	{8'd104,8'd19} : s = 492;
	{8'd104,8'd20} : s = 426;
	{8'd104,8'd21} : s = 490;
	{8'd104,8'd22} : s = 489;
	{8'd104,8'd23} : s = 508;
	{8'd104,8'd24} : s = 2;
	{8'd104,8'd25} : s = 48;
	{8'd104,8'd26} : s = 40;
	{8'd104,8'd27} : s = 168;
	{8'd104,8'd28} : s = 36;
	{8'd104,8'd29} : s = 164;
	{8'd104,8'd30} : s = 162;
	{8'd104,8'd31} : s = 323;
	{8'd104,8'd32} : s = 34;
	{8'd104,8'd33} : s = 161;
	{8'd104,8'd34} : s = 152;
	{8'd104,8'd35} : s = 312;
	{8'd104,8'd36} : s = 148;
	{8'd104,8'd37} : s = 308;
	{8'd104,8'd38} : s = 306;
	{8'd104,8'd39} : s = 425;
	{8'd104,8'd40} : s = 33;
	{8'd104,8'd41} : s = 146;
	{8'd104,8'd42} : s = 145;
	{8'd104,8'd43} : s = 305;
	{8'd104,8'd44} : s = 140;
	{8'd104,8'd45} : s = 300;
	{8'd104,8'd46} : s = 298;
	{8'd104,8'd47} : s = 422;
	{8'd104,8'd48} : s = 138;
	{8'd104,8'd49} : s = 297;
	{8'd104,8'd50} : s = 294;
	{8'd104,8'd51} : s = 421;
	{8'd104,8'd52} : s = 293;
	{8'd104,8'd53} : s = 419;
	{8'd104,8'd54} : s = 412;
	{8'd104,8'd55} : s = 486;
	{8'd104,8'd56} : s = 24;
	{8'd104,8'd57} : s = 137;
	{8'd104,8'd58} : s = 134;
	{8'd104,8'd59} : s = 291;
	{8'd104,8'd60} : s = 133;
	{8'd104,8'd61} : s = 284;
	{8'd104,8'd62} : s = 282;
	{8'd104,8'd63} : s = 410;
	{8'd104,8'd64} : s = 131;
	{8'd104,8'd65} : s = 281;
	{8'd104,8'd66} : s = 278;
	{8'd104,8'd67} : s = 409;
	{8'd104,8'd68} : s = 277;
	{8'd104,8'd69} : s = 406;
	{8'd104,8'd70} : s = 405;
	{8'd104,8'd71} : s = 485;
	{8'd104,8'd72} : s = 112;
	{8'd104,8'd73} : s = 275;
	{8'd104,8'd74} : s = 270;
	{8'd104,8'd75} : s = 403;
	{8'd104,8'd76} : s = 269;
	{8'd104,8'd77} : s = 398;
	{8'd104,8'd78} : s = 397;
	{8'd104,8'd79} : s = 483;
	{8'd104,8'd80} : s = 267;
	{8'd104,8'd81} : s = 395;
	{8'd104,8'd82} : s = 391;
	{8'd104,8'd83} : s = 476;
	{8'd104,8'd84} : s = 376;
	{8'd104,8'd85} : s = 474;
	{8'd104,8'd86} : s = 473;
	{8'd104,8'd87} : s = 506;
	{8'd104,8'd88} : s = 20;
	{8'd104,8'd89} : s = 104;
	{8'd104,8'd90} : s = 100;
	{8'd104,8'd91} : s = 263;
	{8'd104,8'd92} : s = 98;
	{8'd104,8'd93} : s = 240;
	{8'd104,8'd94} : s = 232;
	{8'd104,8'd95} : s = 372;
	{8'd104,8'd96} : s = 97;
	{8'd104,8'd97} : s = 228;
	{8'd104,8'd98} : s = 226;
	{8'd104,8'd99} : s = 370;
	{8'd104,8'd100} : s = 225;
	{8'd104,8'd101} : s = 369;
	{8'd104,8'd102} : s = 364;
	{8'd104,8'd103} : s = 470;
	{8'd104,8'd104} : s = 88;
	{8'd104,8'd105} : s = 216;
	{8'd104,8'd106} : s = 212;
	{8'd104,8'd107} : s = 362;
	{8'd104,8'd108} : s = 210;
	{8'd104,8'd109} : s = 361;
	{8'd104,8'd110} : s = 358;
	{8'd104,8'd111} : s = 469;
	{8'd104,8'd112} : s = 209;
	{8'd104,8'd113} : s = 357;
	{8'd104,8'd114} : s = 355;
	{8'd104,8'd115} : s = 467;
	{8'd104,8'd116} : s = 348;
	{8'd104,8'd117} : s = 462;
	{8'd104,8'd118} : s = 461;
	{8'd104,8'd119} : s = 505;
	{8'd104,8'd120} : s = 84;
	{8'd104,8'd121} : s = 204;
	{8'd104,8'd122} : s = 202;
	{8'd104,8'd123} : s = 346;
	{8'd104,8'd124} : s = 201;
	{8'd104,8'd125} : s = 345;
	{8'd104,8'd126} : s = 342;
	{8'd104,8'd127} : s = 459;
	{8'd104,8'd128} : s = 198;
	{8'd104,8'd129} : s = 341;
	{8'd104,8'd130} : s = 339;
	{8'd104,8'd131} : s = 455;
	{8'd104,8'd132} : s = 334;
	{8'd104,8'd133} : s = 444;
	{8'd104,8'd134} : s = 442;
	{8'd104,8'd135} : s = 502;
	{8'd104,8'd136} : s = 197;
	{8'd104,8'd137} : s = 333;
	{8'd104,8'd138} : s = 331;
	{8'd104,8'd139} : s = 441;
	{8'd104,8'd140} : s = 327;
	{8'd104,8'd141} : s = 438;
	{8'd104,8'd142} : s = 437;
	{8'd104,8'd143} : s = 501;
	{8'd104,8'd144} : s = 316;
	{8'd104,8'd145} : s = 435;
	{8'd104,8'd146} : s = 430;
	{8'd104,8'd147} : s = 499;
	{8'd104,8'd148} : s = 429;
	{8'd104,8'd149} : s = 494;
	{8'd104,8'd150} : s = 493;
	{8'd104,8'd151} : s = 510;
	{8'd104,8'd152} : s = 1;
	{8'd104,8'd153} : s = 18;
	{8'd104,8'd154} : s = 17;
	{8'd104,8'd155} : s = 82;
	{8'd104,8'd156} : s = 12;
	{8'd104,8'd157} : s = 81;
	{8'd104,8'd158} : s = 76;
	{8'd104,8'd159} : s = 195;
	{8'd104,8'd160} : s = 10;
	{8'd104,8'd161} : s = 74;
	{8'd104,8'd162} : s = 73;
	{8'd104,8'd163} : s = 184;
	{8'd104,8'd164} : s = 70;
	{8'd104,8'd165} : s = 180;
	{8'd104,8'd166} : s = 178;
	{8'd104,8'd167} : s = 314;
	{8'd104,8'd168} : s = 9;
	{8'd104,8'd169} : s = 69;
	{8'd104,8'd170} : s = 67;
	{8'd104,8'd171} : s = 177;
	{8'd104,8'd172} : s = 56;
	{8'd104,8'd173} : s = 172;
	{8'd104,8'd174} : s = 170;
	{8'd104,8'd175} : s = 313;
	{8'd104,8'd176} : s = 52;
	{8'd104,8'd177} : s = 169;
	{8'd104,8'd178} : s = 166;
	{8'd104,8'd179} : s = 310;
	{8'd104,8'd180} : s = 165;
	{8'd104,8'd181} : s = 309;
	{8'd104,8'd182} : s = 307;
	{8'd104,8'd183} : s = 427;
	{8'd104,8'd184} : s = 6;
	{8'd104,8'd185} : s = 50;
	{8'd104,8'd186} : s = 49;
	{8'd104,8'd187} : s = 163;
	{8'd104,8'd188} : s = 44;
	{8'd104,8'd189} : s = 156;
	{8'd104,8'd190} : s = 154;
	{8'd104,8'd191} : s = 302;
	{8'd104,8'd192} : s = 42;
	{8'd104,8'd193} : s = 153;
	{8'd104,8'd194} : s = 150;
	{8'd104,8'd195} : s = 301;
	{8'd104,8'd196} : s = 149;
	{8'd104,8'd197} : s = 299;
	{8'd104,8'd198} : s = 295;
	{8'd104,8'd199} : s = 423;
	{8'd104,8'd200} : s = 41;
	{8'd104,8'd201} : s = 147;
	{8'd104,8'd202} : s = 142;
	{8'd104,8'd203} : s = 286;
	{8'd104,8'd204} : s = 141;
	{8'd104,8'd205} : s = 285;
	{8'd104,8'd206} : s = 283;
	{8'd104,8'd207} : s = 414;
	{8'd104,8'd208} : s = 139;
	{8'd104,8'd209} : s = 279;
	{8'd104,8'd210} : s = 271;
	{8'd104,8'd211} : s = 413;
	{8'd104,8'd212} : s = 248;
	{8'd104,8'd213} : s = 411;
	{8'd104,8'd214} : s = 407;
	{8'd104,8'd215} : s = 491;
	{8'd104,8'd216} : s = 5;
	{8'd104,8'd217} : s = 38;
	{8'd104,8'd218} : s = 37;
	{8'd104,8'd219} : s = 135;
	{8'd104,8'd220} : s = 35;
	{8'd104,8'd221} : s = 120;
	{8'd104,8'd222} : s = 116;
	{8'd104,8'd223} : s = 244;
	{8'd104,8'd224} : s = 28;
	{8'd104,8'd225} : s = 114;
	{8'd104,8'd226} : s = 113;
	{8'd104,8'd227} : s = 242;
	{8'd104,8'd228} : s = 108;
	{8'd104,8'd229} : s = 241;
	{8'd104,8'd230} : s = 236;
	{8'd104,8'd231} : s = 399;
	{8'd104,8'd232} : s = 26;
	{8'd104,8'd233} : s = 106;
	{8'd104,8'd234} : s = 105;
	{8'd104,8'd235} : s = 234;
	{8'd104,8'd236} : s = 102;
	{8'd104,8'd237} : s = 233;
	{8'd104,8'd238} : s = 230;
	{8'd104,8'd239} : s = 380;
	{8'd104,8'd240} : s = 101;
	{8'd104,8'd241} : s = 229;
	{8'd104,8'd242} : s = 227;
	{8'd104,8'd243} : s = 378;
	{8'd104,8'd244} : s = 220;
	{8'd104,8'd245} : s = 377;
	{8'd104,8'd246} : s = 374;
	{8'd104,8'd247} : s = 487;
	{8'd104,8'd248} : s = 25;
	{8'd104,8'd249} : s = 99;
	{8'd104,8'd250} : s = 92;
	{8'd104,8'd251} : s = 218;
	{8'd104,8'd252} : s = 90;
	{8'd104,8'd253} : s = 217;
	{8'd104,8'd254} : s = 214;
	{8'd104,8'd255} : s = 373;
	{8'd105,8'd0} : s = 338;
	{8'd105,8'd1} : s = 337;
	{8'd105,8'd2} : s = 454;
	{8'd105,8'd3} : s = 332;
	{8'd105,8'd4} : s = 453;
	{8'd105,8'd5} : s = 451;
	{8'd105,8'd6} : s = 498;
	{8'd105,8'd7} : s = 176;
	{8'd105,8'd8} : s = 330;
	{8'd105,8'd9} : s = 329;
	{8'd105,8'd10} : s = 440;
	{8'd105,8'd11} : s = 326;
	{8'd105,8'd12} : s = 436;
	{8'd105,8'd13} : s = 434;
	{8'd105,8'd14} : s = 497;
	{8'd105,8'd15} : s = 325;
	{8'd105,8'd16} : s = 433;
	{8'd105,8'd17} : s = 428;
	{8'd105,8'd18} : s = 492;
	{8'd105,8'd19} : s = 426;
	{8'd105,8'd20} : s = 490;
	{8'd105,8'd21} : s = 489;
	{8'd105,8'd22} : s = 508;
	{8'd105,8'd23} : s = 2;
	{8'd105,8'd24} : s = 48;
	{8'd105,8'd25} : s = 40;
	{8'd105,8'd26} : s = 168;
	{8'd105,8'd27} : s = 36;
	{8'd105,8'd28} : s = 164;
	{8'd105,8'd29} : s = 162;
	{8'd105,8'd30} : s = 323;
	{8'd105,8'd31} : s = 34;
	{8'd105,8'd32} : s = 161;
	{8'd105,8'd33} : s = 152;
	{8'd105,8'd34} : s = 312;
	{8'd105,8'd35} : s = 148;
	{8'd105,8'd36} : s = 308;
	{8'd105,8'd37} : s = 306;
	{8'd105,8'd38} : s = 425;
	{8'd105,8'd39} : s = 33;
	{8'd105,8'd40} : s = 146;
	{8'd105,8'd41} : s = 145;
	{8'd105,8'd42} : s = 305;
	{8'd105,8'd43} : s = 140;
	{8'd105,8'd44} : s = 300;
	{8'd105,8'd45} : s = 298;
	{8'd105,8'd46} : s = 422;
	{8'd105,8'd47} : s = 138;
	{8'd105,8'd48} : s = 297;
	{8'd105,8'd49} : s = 294;
	{8'd105,8'd50} : s = 421;
	{8'd105,8'd51} : s = 293;
	{8'd105,8'd52} : s = 419;
	{8'd105,8'd53} : s = 412;
	{8'd105,8'd54} : s = 486;
	{8'd105,8'd55} : s = 24;
	{8'd105,8'd56} : s = 137;
	{8'd105,8'd57} : s = 134;
	{8'd105,8'd58} : s = 291;
	{8'd105,8'd59} : s = 133;
	{8'd105,8'd60} : s = 284;
	{8'd105,8'd61} : s = 282;
	{8'd105,8'd62} : s = 410;
	{8'd105,8'd63} : s = 131;
	{8'd105,8'd64} : s = 281;
	{8'd105,8'd65} : s = 278;
	{8'd105,8'd66} : s = 409;
	{8'd105,8'd67} : s = 277;
	{8'd105,8'd68} : s = 406;
	{8'd105,8'd69} : s = 405;
	{8'd105,8'd70} : s = 485;
	{8'd105,8'd71} : s = 112;
	{8'd105,8'd72} : s = 275;
	{8'd105,8'd73} : s = 270;
	{8'd105,8'd74} : s = 403;
	{8'd105,8'd75} : s = 269;
	{8'd105,8'd76} : s = 398;
	{8'd105,8'd77} : s = 397;
	{8'd105,8'd78} : s = 483;
	{8'd105,8'd79} : s = 267;
	{8'd105,8'd80} : s = 395;
	{8'd105,8'd81} : s = 391;
	{8'd105,8'd82} : s = 476;
	{8'd105,8'd83} : s = 376;
	{8'd105,8'd84} : s = 474;
	{8'd105,8'd85} : s = 473;
	{8'd105,8'd86} : s = 506;
	{8'd105,8'd87} : s = 20;
	{8'd105,8'd88} : s = 104;
	{8'd105,8'd89} : s = 100;
	{8'd105,8'd90} : s = 263;
	{8'd105,8'd91} : s = 98;
	{8'd105,8'd92} : s = 240;
	{8'd105,8'd93} : s = 232;
	{8'd105,8'd94} : s = 372;
	{8'd105,8'd95} : s = 97;
	{8'd105,8'd96} : s = 228;
	{8'd105,8'd97} : s = 226;
	{8'd105,8'd98} : s = 370;
	{8'd105,8'd99} : s = 225;
	{8'd105,8'd100} : s = 369;
	{8'd105,8'd101} : s = 364;
	{8'd105,8'd102} : s = 470;
	{8'd105,8'd103} : s = 88;
	{8'd105,8'd104} : s = 216;
	{8'd105,8'd105} : s = 212;
	{8'd105,8'd106} : s = 362;
	{8'd105,8'd107} : s = 210;
	{8'd105,8'd108} : s = 361;
	{8'd105,8'd109} : s = 358;
	{8'd105,8'd110} : s = 469;
	{8'd105,8'd111} : s = 209;
	{8'd105,8'd112} : s = 357;
	{8'd105,8'd113} : s = 355;
	{8'd105,8'd114} : s = 467;
	{8'd105,8'd115} : s = 348;
	{8'd105,8'd116} : s = 462;
	{8'd105,8'd117} : s = 461;
	{8'd105,8'd118} : s = 505;
	{8'd105,8'd119} : s = 84;
	{8'd105,8'd120} : s = 204;
	{8'd105,8'd121} : s = 202;
	{8'd105,8'd122} : s = 346;
	{8'd105,8'd123} : s = 201;
	{8'd105,8'd124} : s = 345;
	{8'd105,8'd125} : s = 342;
	{8'd105,8'd126} : s = 459;
	{8'd105,8'd127} : s = 198;
	{8'd105,8'd128} : s = 341;
	{8'd105,8'd129} : s = 339;
	{8'd105,8'd130} : s = 455;
	{8'd105,8'd131} : s = 334;
	{8'd105,8'd132} : s = 444;
	{8'd105,8'd133} : s = 442;
	{8'd105,8'd134} : s = 502;
	{8'd105,8'd135} : s = 197;
	{8'd105,8'd136} : s = 333;
	{8'd105,8'd137} : s = 331;
	{8'd105,8'd138} : s = 441;
	{8'd105,8'd139} : s = 327;
	{8'd105,8'd140} : s = 438;
	{8'd105,8'd141} : s = 437;
	{8'd105,8'd142} : s = 501;
	{8'd105,8'd143} : s = 316;
	{8'd105,8'd144} : s = 435;
	{8'd105,8'd145} : s = 430;
	{8'd105,8'd146} : s = 499;
	{8'd105,8'd147} : s = 429;
	{8'd105,8'd148} : s = 494;
	{8'd105,8'd149} : s = 493;
	{8'd105,8'd150} : s = 510;
	{8'd105,8'd151} : s = 1;
	{8'd105,8'd152} : s = 18;
	{8'd105,8'd153} : s = 17;
	{8'd105,8'd154} : s = 82;
	{8'd105,8'd155} : s = 12;
	{8'd105,8'd156} : s = 81;
	{8'd105,8'd157} : s = 76;
	{8'd105,8'd158} : s = 195;
	{8'd105,8'd159} : s = 10;
	{8'd105,8'd160} : s = 74;
	{8'd105,8'd161} : s = 73;
	{8'd105,8'd162} : s = 184;
	{8'd105,8'd163} : s = 70;
	{8'd105,8'd164} : s = 180;
	{8'd105,8'd165} : s = 178;
	{8'd105,8'd166} : s = 314;
	{8'd105,8'd167} : s = 9;
	{8'd105,8'd168} : s = 69;
	{8'd105,8'd169} : s = 67;
	{8'd105,8'd170} : s = 177;
	{8'd105,8'd171} : s = 56;
	{8'd105,8'd172} : s = 172;
	{8'd105,8'd173} : s = 170;
	{8'd105,8'd174} : s = 313;
	{8'd105,8'd175} : s = 52;
	{8'd105,8'd176} : s = 169;
	{8'd105,8'd177} : s = 166;
	{8'd105,8'd178} : s = 310;
	{8'd105,8'd179} : s = 165;
	{8'd105,8'd180} : s = 309;
	{8'd105,8'd181} : s = 307;
	{8'd105,8'd182} : s = 427;
	{8'd105,8'd183} : s = 6;
	{8'd105,8'd184} : s = 50;
	{8'd105,8'd185} : s = 49;
	{8'd105,8'd186} : s = 163;
	{8'd105,8'd187} : s = 44;
	{8'd105,8'd188} : s = 156;
	{8'd105,8'd189} : s = 154;
	{8'd105,8'd190} : s = 302;
	{8'd105,8'd191} : s = 42;
	{8'd105,8'd192} : s = 153;
	{8'd105,8'd193} : s = 150;
	{8'd105,8'd194} : s = 301;
	{8'd105,8'd195} : s = 149;
	{8'd105,8'd196} : s = 299;
	{8'd105,8'd197} : s = 295;
	{8'd105,8'd198} : s = 423;
	{8'd105,8'd199} : s = 41;
	{8'd105,8'd200} : s = 147;
	{8'd105,8'd201} : s = 142;
	{8'd105,8'd202} : s = 286;
	{8'd105,8'd203} : s = 141;
	{8'd105,8'd204} : s = 285;
	{8'd105,8'd205} : s = 283;
	{8'd105,8'd206} : s = 414;
	{8'd105,8'd207} : s = 139;
	{8'd105,8'd208} : s = 279;
	{8'd105,8'd209} : s = 271;
	{8'd105,8'd210} : s = 413;
	{8'd105,8'd211} : s = 248;
	{8'd105,8'd212} : s = 411;
	{8'd105,8'd213} : s = 407;
	{8'd105,8'd214} : s = 491;
	{8'd105,8'd215} : s = 5;
	{8'd105,8'd216} : s = 38;
	{8'd105,8'd217} : s = 37;
	{8'd105,8'd218} : s = 135;
	{8'd105,8'd219} : s = 35;
	{8'd105,8'd220} : s = 120;
	{8'd105,8'd221} : s = 116;
	{8'd105,8'd222} : s = 244;
	{8'd105,8'd223} : s = 28;
	{8'd105,8'd224} : s = 114;
	{8'd105,8'd225} : s = 113;
	{8'd105,8'd226} : s = 242;
	{8'd105,8'd227} : s = 108;
	{8'd105,8'd228} : s = 241;
	{8'd105,8'd229} : s = 236;
	{8'd105,8'd230} : s = 399;
	{8'd105,8'd231} : s = 26;
	{8'd105,8'd232} : s = 106;
	{8'd105,8'd233} : s = 105;
	{8'd105,8'd234} : s = 234;
	{8'd105,8'd235} : s = 102;
	{8'd105,8'd236} : s = 233;
	{8'd105,8'd237} : s = 230;
	{8'd105,8'd238} : s = 380;
	{8'd105,8'd239} : s = 101;
	{8'd105,8'd240} : s = 229;
	{8'd105,8'd241} : s = 227;
	{8'd105,8'd242} : s = 378;
	{8'd105,8'd243} : s = 220;
	{8'd105,8'd244} : s = 377;
	{8'd105,8'd245} : s = 374;
	{8'd105,8'd246} : s = 487;
	{8'd105,8'd247} : s = 25;
	{8'd105,8'd248} : s = 99;
	{8'd105,8'd249} : s = 92;
	{8'd105,8'd250} : s = 218;
	{8'd105,8'd251} : s = 90;
	{8'd105,8'd252} : s = 217;
	{8'd105,8'd253} : s = 214;
	{8'd105,8'd254} : s = 373;
	{8'd105,8'd255} : s = 89;
	{8'd106,8'd0} : s = 337;
	{8'd106,8'd1} : s = 454;
	{8'd106,8'd2} : s = 332;
	{8'd106,8'd3} : s = 453;
	{8'd106,8'd4} : s = 451;
	{8'd106,8'd5} : s = 498;
	{8'd106,8'd6} : s = 176;
	{8'd106,8'd7} : s = 330;
	{8'd106,8'd8} : s = 329;
	{8'd106,8'd9} : s = 440;
	{8'd106,8'd10} : s = 326;
	{8'd106,8'd11} : s = 436;
	{8'd106,8'd12} : s = 434;
	{8'd106,8'd13} : s = 497;
	{8'd106,8'd14} : s = 325;
	{8'd106,8'd15} : s = 433;
	{8'd106,8'd16} : s = 428;
	{8'd106,8'd17} : s = 492;
	{8'd106,8'd18} : s = 426;
	{8'd106,8'd19} : s = 490;
	{8'd106,8'd20} : s = 489;
	{8'd106,8'd21} : s = 508;
	{8'd106,8'd22} : s = 2;
	{8'd106,8'd23} : s = 48;
	{8'd106,8'd24} : s = 40;
	{8'd106,8'd25} : s = 168;
	{8'd106,8'd26} : s = 36;
	{8'd106,8'd27} : s = 164;
	{8'd106,8'd28} : s = 162;
	{8'd106,8'd29} : s = 323;
	{8'd106,8'd30} : s = 34;
	{8'd106,8'd31} : s = 161;
	{8'd106,8'd32} : s = 152;
	{8'd106,8'd33} : s = 312;
	{8'd106,8'd34} : s = 148;
	{8'd106,8'd35} : s = 308;
	{8'd106,8'd36} : s = 306;
	{8'd106,8'd37} : s = 425;
	{8'd106,8'd38} : s = 33;
	{8'd106,8'd39} : s = 146;
	{8'd106,8'd40} : s = 145;
	{8'd106,8'd41} : s = 305;
	{8'd106,8'd42} : s = 140;
	{8'd106,8'd43} : s = 300;
	{8'd106,8'd44} : s = 298;
	{8'd106,8'd45} : s = 422;
	{8'd106,8'd46} : s = 138;
	{8'd106,8'd47} : s = 297;
	{8'd106,8'd48} : s = 294;
	{8'd106,8'd49} : s = 421;
	{8'd106,8'd50} : s = 293;
	{8'd106,8'd51} : s = 419;
	{8'd106,8'd52} : s = 412;
	{8'd106,8'd53} : s = 486;
	{8'd106,8'd54} : s = 24;
	{8'd106,8'd55} : s = 137;
	{8'd106,8'd56} : s = 134;
	{8'd106,8'd57} : s = 291;
	{8'd106,8'd58} : s = 133;
	{8'd106,8'd59} : s = 284;
	{8'd106,8'd60} : s = 282;
	{8'd106,8'd61} : s = 410;
	{8'd106,8'd62} : s = 131;
	{8'd106,8'd63} : s = 281;
	{8'd106,8'd64} : s = 278;
	{8'd106,8'd65} : s = 409;
	{8'd106,8'd66} : s = 277;
	{8'd106,8'd67} : s = 406;
	{8'd106,8'd68} : s = 405;
	{8'd106,8'd69} : s = 485;
	{8'd106,8'd70} : s = 112;
	{8'd106,8'd71} : s = 275;
	{8'd106,8'd72} : s = 270;
	{8'd106,8'd73} : s = 403;
	{8'd106,8'd74} : s = 269;
	{8'd106,8'd75} : s = 398;
	{8'd106,8'd76} : s = 397;
	{8'd106,8'd77} : s = 483;
	{8'd106,8'd78} : s = 267;
	{8'd106,8'd79} : s = 395;
	{8'd106,8'd80} : s = 391;
	{8'd106,8'd81} : s = 476;
	{8'd106,8'd82} : s = 376;
	{8'd106,8'd83} : s = 474;
	{8'd106,8'd84} : s = 473;
	{8'd106,8'd85} : s = 506;
	{8'd106,8'd86} : s = 20;
	{8'd106,8'd87} : s = 104;
	{8'd106,8'd88} : s = 100;
	{8'd106,8'd89} : s = 263;
	{8'd106,8'd90} : s = 98;
	{8'd106,8'd91} : s = 240;
	{8'd106,8'd92} : s = 232;
	{8'd106,8'd93} : s = 372;
	{8'd106,8'd94} : s = 97;
	{8'd106,8'd95} : s = 228;
	{8'd106,8'd96} : s = 226;
	{8'd106,8'd97} : s = 370;
	{8'd106,8'd98} : s = 225;
	{8'd106,8'd99} : s = 369;
	{8'd106,8'd100} : s = 364;
	{8'd106,8'd101} : s = 470;
	{8'd106,8'd102} : s = 88;
	{8'd106,8'd103} : s = 216;
	{8'd106,8'd104} : s = 212;
	{8'd106,8'd105} : s = 362;
	{8'd106,8'd106} : s = 210;
	{8'd106,8'd107} : s = 361;
	{8'd106,8'd108} : s = 358;
	{8'd106,8'd109} : s = 469;
	{8'd106,8'd110} : s = 209;
	{8'd106,8'd111} : s = 357;
	{8'd106,8'd112} : s = 355;
	{8'd106,8'd113} : s = 467;
	{8'd106,8'd114} : s = 348;
	{8'd106,8'd115} : s = 462;
	{8'd106,8'd116} : s = 461;
	{8'd106,8'd117} : s = 505;
	{8'd106,8'd118} : s = 84;
	{8'd106,8'd119} : s = 204;
	{8'd106,8'd120} : s = 202;
	{8'd106,8'd121} : s = 346;
	{8'd106,8'd122} : s = 201;
	{8'd106,8'd123} : s = 345;
	{8'd106,8'd124} : s = 342;
	{8'd106,8'd125} : s = 459;
	{8'd106,8'd126} : s = 198;
	{8'd106,8'd127} : s = 341;
	{8'd106,8'd128} : s = 339;
	{8'd106,8'd129} : s = 455;
	{8'd106,8'd130} : s = 334;
	{8'd106,8'd131} : s = 444;
	{8'd106,8'd132} : s = 442;
	{8'd106,8'd133} : s = 502;
	{8'd106,8'd134} : s = 197;
	{8'd106,8'd135} : s = 333;
	{8'd106,8'd136} : s = 331;
	{8'd106,8'd137} : s = 441;
	{8'd106,8'd138} : s = 327;
	{8'd106,8'd139} : s = 438;
	{8'd106,8'd140} : s = 437;
	{8'd106,8'd141} : s = 501;
	{8'd106,8'd142} : s = 316;
	{8'd106,8'd143} : s = 435;
	{8'd106,8'd144} : s = 430;
	{8'd106,8'd145} : s = 499;
	{8'd106,8'd146} : s = 429;
	{8'd106,8'd147} : s = 494;
	{8'd106,8'd148} : s = 493;
	{8'd106,8'd149} : s = 510;
	{8'd106,8'd150} : s = 1;
	{8'd106,8'd151} : s = 18;
	{8'd106,8'd152} : s = 17;
	{8'd106,8'd153} : s = 82;
	{8'd106,8'd154} : s = 12;
	{8'd106,8'd155} : s = 81;
	{8'd106,8'd156} : s = 76;
	{8'd106,8'd157} : s = 195;
	{8'd106,8'd158} : s = 10;
	{8'd106,8'd159} : s = 74;
	{8'd106,8'd160} : s = 73;
	{8'd106,8'd161} : s = 184;
	{8'd106,8'd162} : s = 70;
	{8'd106,8'd163} : s = 180;
	{8'd106,8'd164} : s = 178;
	{8'd106,8'd165} : s = 314;
	{8'd106,8'd166} : s = 9;
	{8'd106,8'd167} : s = 69;
	{8'd106,8'd168} : s = 67;
	{8'd106,8'd169} : s = 177;
	{8'd106,8'd170} : s = 56;
	{8'd106,8'd171} : s = 172;
	{8'd106,8'd172} : s = 170;
	{8'd106,8'd173} : s = 313;
	{8'd106,8'd174} : s = 52;
	{8'd106,8'd175} : s = 169;
	{8'd106,8'd176} : s = 166;
	{8'd106,8'd177} : s = 310;
	{8'd106,8'd178} : s = 165;
	{8'd106,8'd179} : s = 309;
	{8'd106,8'd180} : s = 307;
	{8'd106,8'd181} : s = 427;
	{8'd106,8'd182} : s = 6;
	{8'd106,8'd183} : s = 50;
	{8'd106,8'd184} : s = 49;
	{8'd106,8'd185} : s = 163;
	{8'd106,8'd186} : s = 44;
	{8'd106,8'd187} : s = 156;
	{8'd106,8'd188} : s = 154;
	{8'd106,8'd189} : s = 302;
	{8'd106,8'd190} : s = 42;
	{8'd106,8'd191} : s = 153;
	{8'd106,8'd192} : s = 150;
	{8'd106,8'd193} : s = 301;
	{8'd106,8'd194} : s = 149;
	{8'd106,8'd195} : s = 299;
	{8'd106,8'd196} : s = 295;
	{8'd106,8'd197} : s = 423;
	{8'd106,8'd198} : s = 41;
	{8'd106,8'd199} : s = 147;
	{8'd106,8'd200} : s = 142;
	{8'd106,8'd201} : s = 286;
	{8'd106,8'd202} : s = 141;
	{8'd106,8'd203} : s = 285;
	{8'd106,8'd204} : s = 283;
	{8'd106,8'd205} : s = 414;
	{8'd106,8'd206} : s = 139;
	{8'd106,8'd207} : s = 279;
	{8'd106,8'd208} : s = 271;
	{8'd106,8'd209} : s = 413;
	{8'd106,8'd210} : s = 248;
	{8'd106,8'd211} : s = 411;
	{8'd106,8'd212} : s = 407;
	{8'd106,8'd213} : s = 491;
	{8'd106,8'd214} : s = 5;
	{8'd106,8'd215} : s = 38;
	{8'd106,8'd216} : s = 37;
	{8'd106,8'd217} : s = 135;
	{8'd106,8'd218} : s = 35;
	{8'd106,8'd219} : s = 120;
	{8'd106,8'd220} : s = 116;
	{8'd106,8'd221} : s = 244;
	{8'd106,8'd222} : s = 28;
	{8'd106,8'd223} : s = 114;
	{8'd106,8'd224} : s = 113;
	{8'd106,8'd225} : s = 242;
	{8'd106,8'd226} : s = 108;
	{8'd106,8'd227} : s = 241;
	{8'd106,8'd228} : s = 236;
	{8'd106,8'd229} : s = 399;
	{8'd106,8'd230} : s = 26;
	{8'd106,8'd231} : s = 106;
	{8'd106,8'd232} : s = 105;
	{8'd106,8'd233} : s = 234;
	{8'd106,8'd234} : s = 102;
	{8'd106,8'd235} : s = 233;
	{8'd106,8'd236} : s = 230;
	{8'd106,8'd237} : s = 380;
	{8'd106,8'd238} : s = 101;
	{8'd106,8'd239} : s = 229;
	{8'd106,8'd240} : s = 227;
	{8'd106,8'd241} : s = 378;
	{8'd106,8'd242} : s = 220;
	{8'd106,8'd243} : s = 377;
	{8'd106,8'd244} : s = 374;
	{8'd106,8'd245} : s = 487;
	{8'd106,8'd246} : s = 25;
	{8'd106,8'd247} : s = 99;
	{8'd106,8'd248} : s = 92;
	{8'd106,8'd249} : s = 218;
	{8'd106,8'd250} : s = 90;
	{8'd106,8'd251} : s = 217;
	{8'd106,8'd252} : s = 214;
	{8'd106,8'd253} : s = 373;
	{8'd106,8'd254} : s = 89;
	{8'd106,8'd255} : s = 213;
	{8'd107,8'd0} : s = 454;
	{8'd107,8'd1} : s = 332;
	{8'd107,8'd2} : s = 453;
	{8'd107,8'd3} : s = 451;
	{8'd107,8'd4} : s = 498;
	{8'd107,8'd5} : s = 176;
	{8'd107,8'd6} : s = 330;
	{8'd107,8'd7} : s = 329;
	{8'd107,8'd8} : s = 440;
	{8'd107,8'd9} : s = 326;
	{8'd107,8'd10} : s = 436;
	{8'd107,8'd11} : s = 434;
	{8'd107,8'd12} : s = 497;
	{8'd107,8'd13} : s = 325;
	{8'd107,8'd14} : s = 433;
	{8'd107,8'd15} : s = 428;
	{8'd107,8'd16} : s = 492;
	{8'd107,8'd17} : s = 426;
	{8'd107,8'd18} : s = 490;
	{8'd107,8'd19} : s = 489;
	{8'd107,8'd20} : s = 508;
	{8'd107,8'd21} : s = 2;
	{8'd107,8'd22} : s = 48;
	{8'd107,8'd23} : s = 40;
	{8'd107,8'd24} : s = 168;
	{8'd107,8'd25} : s = 36;
	{8'd107,8'd26} : s = 164;
	{8'd107,8'd27} : s = 162;
	{8'd107,8'd28} : s = 323;
	{8'd107,8'd29} : s = 34;
	{8'd107,8'd30} : s = 161;
	{8'd107,8'd31} : s = 152;
	{8'd107,8'd32} : s = 312;
	{8'd107,8'd33} : s = 148;
	{8'd107,8'd34} : s = 308;
	{8'd107,8'd35} : s = 306;
	{8'd107,8'd36} : s = 425;
	{8'd107,8'd37} : s = 33;
	{8'd107,8'd38} : s = 146;
	{8'd107,8'd39} : s = 145;
	{8'd107,8'd40} : s = 305;
	{8'd107,8'd41} : s = 140;
	{8'd107,8'd42} : s = 300;
	{8'd107,8'd43} : s = 298;
	{8'd107,8'd44} : s = 422;
	{8'd107,8'd45} : s = 138;
	{8'd107,8'd46} : s = 297;
	{8'd107,8'd47} : s = 294;
	{8'd107,8'd48} : s = 421;
	{8'd107,8'd49} : s = 293;
	{8'd107,8'd50} : s = 419;
	{8'd107,8'd51} : s = 412;
	{8'd107,8'd52} : s = 486;
	{8'd107,8'd53} : s = 24;
	{8'd107,8'd54} : s = 137;
	{8'd107,8'd55} : s = 134;
	{8'd107,8'd56} : s = 291;
	{8'd107,8'd57} : s = 133;
	{8'd107,8'd58} : s = 284;
	{8'd107,8'd59} : s = 282;
	{8'd107,8'd60} : s = 410;
	{8'd107,8'd61} : s = 131;
	{8'd107,8'd62} : s = 281;
	{8'd107,8'd63} : s = 278;
	{8'd107,8'd64} : s = 409;
	{8'd107,8'd65} : s = 277;
	{8'd107,8'd66} : s = 406;
	{8'd107,8'd67} : s = 405;
	{8'd107,8'd68} : s = 485;
	{8'd107,8'd69} : s = 112;
	{8'd107,8'd70} : s = 275;
	{8'd107,8'd71} : s = 270;
	{8'd107,8'd72} : s = 403;
	{8'd107,8'd73} : s = 269;
	{8'd107,8'd74} : s = 398;
	{8'd107,8'd75} : s = 397;
	{8'd107,8'd76} : s = 483;
	{8'd107,8'd77} : s = 267;
	{8'd107,8'd78} : s = 395;
	{8'd107,8'd79} : s = 391;
	{8'd107,8'd80} : s = 476;
	{8'd107,8'd81} : s = 376;
	{8'd107,8'd82} : s = 474;
	{8'd107,8'd83} : s = 473;
	{8'd107,8'd84} : s = 506;
	{8'd107,8'd85} : s = 20;
	{8'd107,8'd86} : s = 104;
	{8'd107,8'd87} : s = 100;
	{8'd107,8'd88} : s = 263;
	{8'd107,8'd89} : s = 98;
	{8'd107,8'd90} : s = 240;
	{8'd107,8'd91} : s = 232;
	{8'd107,8'd92} : s = 372;
	{8'd107,8'd93} : s = 97;
	{8'd107,8'd94} : s = 228;
	{8'd107,8'd95} : s = 226;
	{8'd107,8'd96} : s = 370;
	{8'd107,8'd97} : s = 225;
	{8'd107,8'd98} : s = 369;
	{8'd107,8'd99} : s = 364;
	{8'd107,8'd100} : s = 470;
	{8'd107,8'd101} : s = 88;
	{8'd107,8'd102} : s = 216;
	{8'd107,8'd103} : s = 212;
	{8'd107,8'd104} : s = 362;
	{8'd107,8'd105} : s = 210;
	{8'd107,8'd106} : s = 361;
	{8'd107,8'd107} : s = 358;
	{8'd107,8'd108} : s = 469;
	{8'd107,8'd109} : s = 209;
	{8'd107,8'd110} : s = 357;
	{8'd107,8'd111} : s = 355;
	{8'd107,8'd112} : s = 467;
	{8'd107,8'd113} : s = 348;
	{8'd107,8'd114} : s = 462;
	{8'd107,8'd115} : s = 461;
	{8'd107,8'd116} : s = 505;
	{8'd107,8'd117} : s = 84;
	{8'd107,8'd118} : s = 204;
	{8'd107,8'd119} : s = 202;
	{8'd107,8'd120} : s = 346;
	{8'd107,8'd121} : s = 201;
	{8'd107,8'd122} : s = 345;
	{8'd107,8'd123} : s = 342;
	{8'd107,8'd124} : s = 459;
	{8'd107,8'd125} : s = 198;
	{8'd107,8'd126} : s = 341;
	{8'd107,8'd127} : s = 339;
	{8'd107,8'd128} : s = 455;
	{8'd107,8'd129} : s = 334;
	{8'd107,8'd130} : s = 444;
	{8'd107,8'd131} : s = 442;
	{8'd107,8'd132} : s = 502;
	{8'd107,8'd133} : s = 197;
	{8'd107,8'd134} : s = 333;
	{8'd107,8'd135} : s = 331;
	{8'd107,8'd136} : s = 441;
	{8'd107,8'd137} : s = 327;
	{8'd107,8'd138} : s = 438;
	{8'd107,8'd139} : s = 437;
	{8'd107,8'd140} : s = 501;
	{8'd107,8'd141} : s = 316;
	{8'd107,8'd142} : s = 435;
	{8'd107,8'd143} : s = 430;
	{8'd107,8'd144} : s = 499;
	{8'd107,8'd145} : s = 429;
	{8'd107,8'd146} : s = 494;
	{8'd107,8'd147} : s = 493;
	{8'd107,8'd148} : s = 510;
	{8'd107,8'd149} : s = 1;
	{8'd107,8'd150} : s = 18;
	{8'd107,8'd151} : s = 17;
	{8'd107,8'd152} : s = 82;
	{8'd107,8'd153} : s = 12;
	{8'd107,8'd154} : s = 81;
	{8'd107,8'd155} : s = 76;
	{8'd107,8'd156} : s = 195;
	{8'd107,8'd157} : s = 10;
	{8'd107,8'd158} : s = 74;
	{8'd107,8'd159} : s = 73;
	{8'd107,8'd160} : s = 184;
	{8'd107,8'd161} : s = 70;
	{8'd107,8'd162} : s = 180;
	{8'd107,8'd163} : s = 178;
	{8'd107,8'd164} : s = 314;
	{8'd107,8'd165} : s = 9;
	{8'd107,8'd166} : s = 69;
	{8'd107,8'd167} : s = 67;
	{8'd107,8'd168} : s = 177;
	{8'd107,8'd169} : s = 56;
	{8'd107,8'd170} : s = 172;
	{8'd107,8'd171} : s = 170;
	{8'd107,8'd172} : s = 313;
	{8'd107,8'd173} : s = 52;
	{8'd107,8'd174} : s = 169;
	{8'd107,8'd175} : s = 166;
	{8'd107,8'd176} : s = 310;
	{8'd107,8'd177} : s = 165;
	{8'd107,8'd178} : s = 309;
	{8'd107,8'd179} : s = 307;
	{8'd107,8'd180} : s = 427;
	{8'd107,8'd181} : s = 6;
	{8'd107,8'd182} : s = 50;
	{8'd107,8'd183} : s = 49;
	{8'd107,8'd184} : s = 163;
	{8'd107,8'd185} : s = 44;
	{8'd107,8'd186} : s = 156;
	{8'd107,8'd187} : s = 154;
	{8'd107,8'd188} : s = 302;
	{8'd107,8'd189} : s = 42;
	{8'd107,8'd190} : s = 153;
	{8'd107,8'd191} : s = 150;
	{8'd107,8'd192} : s = 301;
	{8'd107,8'd193} : s = 149;
	{8'd107,8'd194} : s = 299;
	{8'd107,8'd195} : s = 295;
	{8'd107,8'd196} : s = 423;
	{8'd107,8'd197} : s = 41;
	{8'd107,8'd198} : s = 147;
	{8'd107,8'd199} : s = 142;
	{8'd107,8'd200} : s = 286;
	{8'd107,8'd201} : s = 141;
	{8'd107,8'd202} : s = 285;
	{8'd107,8'd203} : s = 283;
	{8'd107,8'd204} : s = 414;
	{8'd107,8'd205} : s = 139;
	{8'd107,8'd206} : s = 279;
	{8'd107,8'd207} : s = 271;
	{8'd107,8'd208} : s = 413;
	{8'd107,8'd209} : s = 248;
	{8'd107,8'd210} : s = 411;
	{8'd107,8'd211} : s = 407;
	{8'd107,8'd212} : s = 491;
	{8'd107,8'd213} : s = 5;
	{8'd107,8'd214} : s = 38;
	{8'd107,8'd215} : s = 37;
	{8'd107,8'd216} : s = 135;
	{8'd107,8'd217} : s = 35;
	{8'd107,8'd218} : s = 120;
	{8'd107,8'd219} : s = 116;
	{8'd107,8'd220} : s = 244;
	{8'd107,8'd221} : s = 28;
	{8'd107,8'd222} : s = 114;
	{8'd107,8'd223} : s = 113;
	{8'd107,8'd224} : s = 242;
	{8'd107,8'd225} : s = 108;
	{8'd107,8'd226} : s = 241;
	{8'd107,8'd227} : s = 236;
	{8'd107,8'd228} : s = 399;
	{8'd107,8'd229} : s = 26;
	{8'd107,8'd230} : s = 106;
	{8'd107,8'd231} : s = 105;
	{8'd107,8'd232} : s = 234;
	{8'd107,8'd233} : s = 102;
	{8'd107,8'd234} : s = 233;
	{8'd107,8'd235} : s = 230;
	{8'd107,8'd236} : s = 380;
	{8'd107,8'd237} : s = 101;
	{8'd107,8'd238} : s = 229;
	{8'd107,8'd239} : s = 227;
	{8'd107,8'd240} : s = 378;
	{8'd107,8'd241} : s = 220;
	{8'd107,8'd242} : s = 377;
	{8'd107,8'd243} : s = 374;
	{8'd107,8'd244} : s = 487;
	{8'd107,8'd245} : s = 25;
	{8'd107,8'd246} : s = 99;
	{8'd107,8'd247} : s = 92;
	{8'd107,8'd248} : s = 218;
	{8'd107,8'd249} : s = 90;
	{8'd107,8'd250} : s = 217;
	{8'd107,8'd251} : s = 214;
	{8'd107,8'd252} : s = 373;
	{8'd107,8'd253} : s = 89;
	{8'd107,8'd254} : s = 213;
	{8'd107,8'd255} : s = 211;
	{8'd108,8'd0} : s = 332;
	{8'd108,8'd1} : s = 453;
	{8'd108,8'd2} : s = 451;
	{8'd108,8'd3} : s = 498;
	{8'd108,8'd4} : s = 176;
	{8'd108,8'd5} : s = 330;
	{8'd108,8'd6} : s = 329;
	{8'd108,8'd7} : s = 440;
	{8'd108,8'd8} : s = 326;
	{8'd108,8'd9} : s = 436;
	{8'd108,8'd10} : s = 434;
	{8'd108,8'd11} : s = 497;
	{8'd108,8'd12} : s = 325;
	{8'd108,8'd13} : s = 433;
	{8'd108,8'd14} : s = 428;
	{8'd108,8'd15} : s = 492;
	{8'd108,8'd16} : s = 426;
	{8'd108,8'd17} : s = 490;
	{8'd108,8'd18} : s = 489;
	{8'd108,8'd19} : s = 508;
	{8'd108,8'd20} : s = 2;
	{8'd108,8'd21} : s = 48;
	{8'd108,8'd22} : s = 40;
	{8'd108,8'd23} : s = 168;
	{8'd108,8'd24} : s = 36;
	{8'd108,8'd25} : s = 164;
	{8'd108,8'd26} : s = 162;
	{8'd108,8'd27} : s = 323;
	{8'd108,8'd28} : s = 34;
	{8'd108,8'd29} : s = 161;
	{8'd108,8'd30} : s = 152;
	{8'd108,8'd31} : s = 312;
	{8'd108,8'd32} : s = 148;
	{8'd108,8'd33} : s = 308;
	{8'd108,8'd34} : s = 306;
	{8'd108,8'd35} : s = 425;
	{8'd108,8'd36} : s = 33;
	{8'd108,8'd37} : s = 146;
	{8'd108,8'd38} : s = 145;
	{8'd108,8'd39} : s = 305;
	{8'd108,8'd40} : s = 140;
	{8'd108,8'd41} : s = 300;
	{8'd108,8'd42} : s = 298;
	{8'd108,8'd43} : s = 422;
	{8'd108,8'd44} : s = 138;
	{8'd108,8'd45} : s = 297;
	{8'd108,8'd46} : s = 294;
	{8'd108,8'd47} : s = 421;
	{8'd108,8'd48} : s = 293;
	{8'd108,8'd49} : s = 419;
	{8'd108,8'd50} : s = 412;
	{8'd108,8'd51} : s = 486;
	{8'd108,8'd52} : s = 24;
	{8'd108,8'd53} : s = 137;
	{8'd108,8'd54} : s = 134;
	{8'd108,8'd55} : s = 291;
	{8'd108,8'd56} : s = 133;
	{8'd108,8'd57} : s = 284;
	{8'd108,8'd58} : s = 282;
	{8'd108,8'd59} : s = 410;
	{8'd108,8'd60} : s = 131;
	{8'd108,8'd61} : s = 281;
	{8'd108,8'd62} : s = 278;
	{8'd108,8'd63} : s = 409;
	{8'd108,8'd64} : s = 277;
	{8'd108,8'd65} : s = 406;
	{8'd108,8'd66} : s = 405;
	{8'd108,8'd67} : s = 485;
	{8'd108,8'd68} : s = 112;
	{8'd108,8'd69} : s = 275;
	{8'd108,8'd70} : s = 270;
	{8'd108,8'd71} : s = 403;
	{8'd108,8'd72} : s = 269;
	{8'd108,8'd73} : s = 398;
	{8'd108,8'd74} : s = 397;
	{8'd108,8'd75} : s = 483;
	{8'd108,8'd76} : s = 267;
	{8'd108,8'd77} : s = 395;
	{8'd108,8'd78} : s = 391;
	{8'd108,8'd79} : s = 476;
	{8'd108,8'd80} : s = 376;
	{8'd108,8'd81} : s = 474;
	{8'd108,8'd82} : s = 473;
	{8'd108,8'd83} : s = 506;
	{8'd108,8'd84} : s = 20;
	{8'd108,8'd85} : s = 104;
	{8'd108,8'd86} : s = 100;
	{8'd108,8'd87} : s = 263;
	{8'd108,8'd88} : s = 98;
	{8'd108,8'd89} : s = 240;
	{8'd108,8'd90} : s = 232;
	{8'd108,8'd91} : s = 372;
	{8'd108,8'd92} : s = 97;
	{8'd108,8'd93} : s = 228;
	{8'd108,8'd94} : s = 226;
	{8'd108,8'd95} : s = 370;
	{8'd108,8'd96} : s = 225;
	{8'd108,8'd97} : s = 369;
	{8'd108,8'd98} : s = 364;
	{8'd108,8'd99} : s = 470;
	{8'd108,8'd100} : s = 88;
	{8'd108,8'd101} : s = 216;
	{8'd108,8'd102} : s = 212;
	{8'd108,8'd103} : s = 362;
	{8'd108,8'd104} : s = 210;
	{8'd108,8'd105} : s = 361;
	{8'd108,8'd106} : s = 358;
	{8'd108,8'd107} : s = 469;
	{8'd108,8'd108} : s = 209;
	{8'd108,8'd109} : s = 357;
	{8'd108,8'd110} : s = 355;
	{8'd108,8'd111} : s = 467;
	{8'd108,8'd112} : s = 348;
	{8'd108,8'd113} : s = 462;
	{8'd108,8'd114} : s = 461;
	{8'd108,8'd115} : s = 505;
	{8'd108,8'd116} : s = 84;
	{8'd108,8'd117} : s = 204;
	{8'd108,8'd118} : s = 202;
	{8'd108,8'd119} : s = 346;
	{8'd108,8'd120} : s = 201;
	{8'd108,8'd121} : s = 345;
	{8'd108,8'd122} : s = 342;
	{8'd108,8'd123} : s = 459;
	{8'd108,8'd124} : s = 198;
	{8'd108,8'd125} : s = 341;
	{8'd108,8'd126} : s = 339;
	{8'd108,8'd127} : s = 455;
	{8'd108,8'd128} : s = 334;
	{8'd108,8'd129} : s = 444;
	{8'd108,8'd130} : s = 442;
	{8'd108,8'd131} : s = 502;
	{8'd108,8'd132} : s = 197;
	{8'd108,8'd133} : s = 333;
	{8'd108,8'd134} : s = 331;
	{8'd108,8'd135} : s = 441;
	{8'd108,8'd136} : s = 327;
	{8'd108,8'd137} : s = 438;
	{8'd108,8'd138} : s = 437;
	{8'd108,8'd139} : s = 501;
	{8'd108,8'd140} : s = 316;
	{8'd108,8'd141} : s = 435;
	{8'd108,8'd142} : s = 430;
	{8'd108,8'd143} : s = 499;
	{8'd108,8'd144} : s = 429;
	{8'd108,8'd145} : s = 494;
	{8'd108,8'd146} : s = 493;
	{8'd108,8'd147} : s = 510;
	{8'd108,8'd148} : s = 1;
	{8'd108,8'd149} : s = 18;
	{8'd108,8'd150} : s = 17;
	{8'd108,8'd151} : s = 82;
	{8'd108,8'd152} : s = 12;
	{8'd108,8'd153} : s = 81;
	{8'd108,8'd154} : s = 76;
	{8'd108,8'd155} : s = 195;
	{8'd108,8'd156} : s = 10;
	{8'd108,8'd157} : s = 74;
	{8'd108,8'd158} : s = 73;
	{8'd108,8'd159} : s = 184;
	{8'd108,8'd160} : s = 70;
	{8'd108,8'd161} : s = 180;
	{8'd108,8'd162} : s = 178;
	{8'd108,8'd163} : s = 314;
	{8'd108,8'd164} : s = 9;
	{8'd108,8'd165} : s = 69;
	{8'd108,8'd166} : s = 67;
	{8'd108,8'd167} : s = 177;
	{8'd108,8'd168} : s = 56;
	{8'd108,8'd169} : s = 172;
	{8'd108,8'd170} : s = 170;
	{8'd108,8'd171} : s = 313;
	{8'd108,8'd172} : s = 52;
	{8'd108,8'd173} : s = 169;
	{8'd108,8'd174} : s = 166;
	{8'd108,8'd175} : s = 310;
	{8'd108,8'd176} : s = 165;
	{8'd108,8'd177} : s = 309;
	{8'd108,8'd178} : s = 307;
	{8'd108,8'd179} : s = 427;
	{8'd108,8'd180} : s = 6;
	{8'd108,8'd181} : s = 50;
	{8'd108,8'd182} : s = 49;
	{8'd108,8'd183} : s = 163;
	{8'd108,8'd184} : s = 44;
	{8'd108,8'd185} : s = 156;
	{8'd108,8'd186} : s = 154;
	{8'd108,8'd187} : s = 302;
	{8'd108,8'd188} : s = 42;
	{8'd108,8'd189} : s = 153;
	{8'd108,8'd190} : s = 150;
	{8'd108,8'd191} : s = 301;
	{8'd108,8'd192} : s = 149;
	{8'd108,8'd193} : s = 299;
	{8'd108,8'd194} : s = 295;
	{8'd108,8'd195} : s = 423;
	{8'd108,8'd196} : s = 41;
	{8'd108,8'd197} : s = 147;
	{8'd108,8'd198} : s = 142;
	{8'd108,8'd199} : s = 286;
	{8'd108,8'd200} : s = 141;
	{8'd108,8'd201} : s = 285;
	{8'd108,8'd202} : s = 283;
	{8'd108,8'd203} : s = 414;
	{8'd108,8'd204} : s = 139;
	{8'd108,8'd205} : s = 279;
	{8'd108,8'd206} : s = 271;
	{8'd108,8'd207} : s = 413;
	{8'd108,8'd208} : s = 248;
	{8'd108,8'd209} : s = 411;
	{8'd108,8'd210} : s = 407;
	{8'd108,8'd211} : s = 491;
	{8'd108,8'd212} : s = 5;
	{8'd108,8'd213} : s = 38;
	{8'd108,8'd214} : s = 37;
	{8'd108,8'd215} : s = 135;
	{8'd108,8'd216} : s = 35;
	{8'd108,8'd217} : s = 120;
	{8'd108,8'd218} : s = 116;
	{8'd108,8'd219} : s = 244;
	{8'd108,8'd220} : s = 28;
	{8'd108,8'd221} : s = 114;
	{8'd108,8'd222} : s = 113;
	{8'd108,8'd223} : s = 242;
	{8'd108,8'd224} : s = 108;
	{8'd108,8'd225} : s = 241;
	{8'd108,8'd226} : s = 236;
	{8'd108,8'd227} : s = 399;
	{8'd108,8'd228} : s = 26;
	{8'd108,8'd229} : s = 106;
	{8'd108,8'd230} : s = 105;
	{8'd108,8'd231} : s = 234;
	{8'd108,8'd232} : s = 102;
	{8'd108,8'd233} : s = 233;
	{8'd108,8'd234} : s = 230;
	{8'd108,8'd235} : s = 380;
	{8'd108,8'd236} : s = 101;
	{8'd108,8'd237} : s = 229;
	{8'd108,8'd238} : s = 227;
	{8'd108,8'd239} : s = 378;
	{8'd108,8'd240} : s = 220;
	{8'd108,8'd241} : s = 377;
	{8'd108,8'd242} : s = 374;
	{8'd108,8'd243} : s = 487;
	{8'd108,8'd244} : s = 25;
	{8'd108,8'd245} : s = 99;
	{8'd108,8'd246} : s = 92;
	{8'd108,8'd247} : s = 218;
	{8'd108,8'd248} : s = 90;
	{8'd108,8'd249} : s = 217;
	{8'd108,8'd250} : s = 214;
	{8'd108,8'd251} : s = 373;
	{8'd108,8'd252} : s = 89;
	{8'd108,8'd253} : s = 213;
	{8'd108,8'd254} : s = 211;
	{8'd108,8'd255} : s = 371;
	{8'd109,8'd0} : s = 453;
	{8'd109,8'd1} : s = 451;
	{8'd109,8'd2} : s = 498;
	{8'd109,8'd3} : s = 176;
	{8'd109,8'd4} : s = 330;
	{8'd109,8'd5} : s = 329;
	{8'd109,8'd6} : s = 440;
	{8'd109,8'd7} : s = 326;
	{8'd109,8'd8} : s = 436;
	{8'd109,8'd9} : s = 434;
	{8'd109,8'd10} : s = 497;
	{8'd109,8'd11} : s = 325;
	{8'd109,8'd12} : s = 433;
	{8'd109,8'd13} : s = 428;
	{8'd109,8'd14} : s = 492;
	{8'd109,8'd15} : s = 426;
	{8'd109,8'd16} : s = 490;
	{8'd109,8'd17} : s = 489;
	{8'd109,8'd18} : s = 508;
	{8'd109,8'd19} : s = 2;
	{8'd109,8'd20} : s = 48;
	{8'd109,8'd21} : s = 40;
	{8'd109,8'd22} : s = 168;
	{8'd109,8'd23} : s = 36;
	{8'd109,8'd24} : s = 164;
	{8'd109,8'd25} : s = 162;
	{8'd109,8'd26} : s = 323;
	{8'd109,8'd27} : s = 34;
	{8'd109,8'd28} : s = 161;
	{8'd109,8'd29} : s = 152;
	{8'd109,8'd30} : s = 312;
	{8'd109,8'd31} : s = 148;
	{8'd109,8'd32} : s = 308;
	{8'd109,8'd33} : s = 306;
	{8'd109,8'd34} : s = 425;
	{8'd109,8'd35} : s = 33;
	{8'd109,8'd36} : s = 146;
	{8'd109,8'd37} : s = 145;
	{8'd109,8'd38} : s = 305;
	{8'd109,8'd39} : s = 140;
	{8'd109,8'd40} : s = 300;
	{8'd109,8'd41} : s = 298;
	{8'd109,8'd42} : s = 422;
	{8'd109,8'd43} : s = 138;
	{8'd109,8'd44} : s = 297;
	{8'd109,8'd45} : s = 294;
	{8'd109,8'd46} : s = 421;
	{8'd109,8'd47} : s = 293;
	{8'd109,8'd48} : s = 419;
	{8'd109,8'd49} : s = 412;
	{8'd109,8'd50} : s = 486;
	{8'd109,8'd51} : s = 24;
	{8'd109,8'd52} : s = 137;
	{8'd109,8'd53} : s = 134;
	{8'd109,8'd54} : s = 291;
	{8'd109,8'd55} : s = 133;
	{8'd109,8'd56} : s = 284;
	{8'd109,8'd57} : s = 282;
	{8'd109,8'd58} : s = 410;
	{8'd109,8'd59} : s = 131;
	{8'd109,8'd60} : s = 281;
	{8'd109,8'd61} : s = 278;
	{8'd109,8'd62} : s = 409;
	{8'd109,8'd63} : s = 277;
	{8'd109,8'd64} : s = 406;
	{8'd109,8'd65} : s = 405;
	{8'd109,8'd66} : s = 485;
	{8'd109,8'd67} : s = 112;
	{8'd109,8'd68} : s = 275;
	{8'd109,8'd69} : s = 270;
	{8'd109,8'd70} : s = 403;
	{8'd109,8'd71} : s = 269;
	{8'd109,8'd72} : s = 398;
	{8'd109,8'd73} : s = 397;
	{8'd109,8'd74} : s = 483;
	{8'd109,8'd75} : s = 267;
	{8'd109,8'd76} : s = 395;
	{8'd109,8'd77} : s = 391;
	{8'd109,8'd78} : s = 476;
	{8'd109,8'd79} : s = 376;
	{8'd109,8'd80} : s = 474;
	{8'd109,8'd81} : s = 473;
	{8'd109,8'd82} : s = 506;
	{8'd109,8'd83} : s = 20;
	{8'd109,8'd84} : s = 104;
	{8'd109,8'd85} : s = 100;
	{8'd109,8'd86} : s = 263;
	{8'd109,8'd87} : s = 98;
	{8'd109,8'd88} : s = 240;
	{8'd109,8'd89} : s = 232;
	{8'd109,8'd90} : s = 372;
	{8'd109,8'd91} : s = 97;
	{8'd109,8'd92} : s = 228;
	{8'd109,8'd93} : s = 226;
	{8'd109,8'd94} : s = 370;
	{8'd109,8'd95} : s = 225;
	{8'd109,8'd96} : s = 369;
	{8'd109,8'd97} : s = 364;
	{8'd109,8'd98} : s = 470;
	{8'd109,8'd99} : s = 88;
	{8'd109,8'd100} : s = 216;
	{8'd109,8'd101} : s = 212;
	{8'd109,8'd102} : s = 362;
	{8'd109,8'd103} : s = 210;
	{8'd109,8'd104} : s = 361;
	{8'd109,8'd105} : s = 358;
	{8'd109,8'd106} : s = 469;
	{8'd109,8'd107} : s = 209;
	{8'd109,8'd108} : s = 357;
	{8'd109,8'd109} : s = 355;
	{8'd109,8'd110} : s = 467;
	{8'd109,8'd111} : s = 348;
	{8'd109,8'd112} : s = 462;
	{8'd109,8'd113} : s = 461;
	{8'd109,8'd114} : s = 505;
	{8'd109,8'd115} : s = 84;
	{8'd109,8'd116} : s = 204;
	{8'd109,8'd117} : s = 202;
	{8'd109,8'd118} : s = 346;
	{8'd109,8'd119} : s = 201;
	{8'd109,8'd120} : s = 345;
	{8'd109,8'd121} : s = 342;
	{8'd109,8'd122} : s = 459;
	{8'd109,8'd123} : s = 198;
	{8'd109,8'd124} : s = 341;
	{8'd109,8'd125} : s = 339;
	{8'd109,8'd126} : s = 455;
	{8'd109,8'd127} : s = 334;
	{8'd109,8'd128} : s = 444;
	{8'd109,8'd129} : s = 442;
	{8'd109,8'd130} : s = 502;
	{8'd109,8'd131} : s = 197;
	{8'd109,8'd132} : s = 333;
	{8'd109,8'd133} : s = 331;
	{8'd109,8'd134} : s = 441;
	{8'd109,8'd135} : s = 327;
	{8'd109,8'd136} : s = 438;
	{8'd109,8'd137} : s = 437;
	{8'd109,8'd138} : s = 501;
	{8'd109,8'd139} : s = 316;
	{8'd109,8'd140} : s = 435;
	{8'd109,8'd141} : s = 430;
	{8'd109,8'd142} : s = 499;
	{8'd109,8'd143} : s = 429;
	{8'd109,8'd144} : s = 494;
	{8'd109,8'd145} : s = 493;
	{8'd109,8'd146} : s = 510;
	{8'd109,8'd147} : s = 1;
	{8'd109,8'd148} : s = 18;
	{8'd109,8'd149} : s = 17;
	{8'd109,8'd150} : s = 82;
	{8'd109,8'd151} : s = 12;
	{8'd109,8'd152} : s = 81;
	{8'd109,8'd153} : s = 76;
	{8'd109,8'd154} : s = 195;
	{8'd109,8'd155} : s = 10;
	{8'd109,8'd156} : s = 74;
	{8'd109,8'd157} : s = 73;
	{8'd109,8'd158} : s = 184;
	{8'd109,8'd159} : s = 70;
	{8'd109,8'd160} : s = 180;
	{8'd109,8'd161} : s = 178;
	{8'd109,8'd162} : s = 314;
	{8'd109,8'd163} : s = 9;
	{8'd109,8'd164} : s = 69;
	{8'd109,8'd165} : s = 67;
	{8'd109,8'd166} : s = 177;
	{8'd109,8'd167} : s = 56;
	{8'd109,8'd168} : s = 172;
	{8'd109,8'd169} : s = 170;
	{8'd109,8'd170} : s = 313;
	{8'd109,8'd171} : s = 52;
	{8'd109,8'd172} : s = 169;
	{8'd109,8'd173} : s = 166;
	{8'd109,8'd174} : s = 310;
	{8'd109,8'd175} : s = 165;
	{8'd109,8'd176} : s = 309;
	{8'd109,8'd177} : s = 307;
	{8'd109,8'd178} : s = 427;
	{8'd109,8'd179} : s = 6;
	{8'd109,8'd180} : s = 50;
	{8'd109,8'd181} : s = 49;
	{8'd109,8'd182} : s = 163;
	{8'd109,8'd183} : s = 44;
	{8'd109,8'd184} : s = 156;
	{8'd109,8'd185} : s = 154;
	{8'd109,8'd186} : s = 302;
	{8'd109,8'd187} : s = 42;
	{8'd109,8'd188} : s = 153;
	{8'd109,8'd189} : s = 150;
	{8'd109,8'd190} : s = 301;
	{8'd109,8'd191} : s = 149;
	{8'd109,8'd192} : s = 299;
	{8'd109,8'd193} : s = 295;
	{8'd109,8'd194} : s = 423;
	{8'd109,8'd195} : s = 41;
	{8'd109,8'd196} : s = 147;
	{8'd109,8'd197} : s = 142;
	{8'd109,8'd198} : s = 286;
	{8'd109,8'd199} : s = 141;
	{8'd109,8'd200} : s = 285;
	{8'd109,8'd201} : s = 283;
	{8'd109,8'd202} : s = 414;
	{8'd109,8'd203} : s = 139;
	{8'd109,8'd204} : s = 279;
	{8'd109,8'd205} : s = 271;
	{8'd109,8'd206} : s = 413;
	{8'd109,8'd207} : s = 248;
	{8'd109,8'd208} : s = 411;
	{8'd109,8'd209} : s = 407;
	{8'd109,8'd210} : s = 491;
	{8'd109,8'd211} : s = 5;
	{8'd109,8'd212} : s = 38;
	{8'd109,8'd213} : s = 37;
	{8'd109,8'd214} : s = 135;
	{8'd109,8'd215} : s = 35;
	{8'd109,8'd216} : s = 120;
	{8'd109,8'd217} : s = 116;
	{8'd109,8'd218} : s = 244;
	{8'd109,8'd219} : s = 28;
	{8'd109,8'd220} : s = 114;
	{8'd109,8'd221} : s = 113;
	{8'd109,8'd222} : s = 242;
	{8'd109,8'd223} : s = 108;
	{8'd109,8'd224} : s = 241;
	{8'd109,8'd225} : s = 236;
	{8'd109,8'd226} : s = 399;
	{8'd109,8'd227} : s = 26;
	{8'd109,8'd228} : s = 106;
	{8'd109,8'd229} : s = 105;
	{8'd109,8'd230} : s = 234;
	{8'd109,8'd231} : s = 102;
	{8'd109,8'd232} : s = 233;
	{8'd109,8'd233} : s = 230;
	{8'd109,8'd234} : s = 380;
	{8'd109,8'd235} : s = 101;
	{8'd109,8'd236} : s = 229;
	{8'd109,8'd237} : s = 227;
	{8'd109,8'd238} : s = 378;
	{8'd109,8'd239} : s = 220;
	{8'd109,8'd240} : s = 377;
	{8'd109,8'd241} : s = 374;
	{8'd109,8'd242} : s = 487;
	{8'd109,8'd243} : s = 25;
	{8'd109,8'd244} : s = 99;
	{8'd109,8'd245} : s = 92;
	{8'd109,8'd246} : s = 218;
	{8'd109,8'd247} : s = 90;
	{8'd109,8'd248} : s = 217;
	{8'd109,8'd249} : s = 214;
	{8'd109,8'd250} : s = 373;
	{8'd109,8'd251} : s = 89;
	{8'd109,8'd252} : s = 213;
	{8'd109,8'd253} : s = 211;
	{8'd109,8'd254} : s = 371;
	{8'd109,8'd255} : s = 206;
	{8'd110,8'd0} : s = 451;
	{8'd110,8'd1} : s = 498;
	{8'd110,8'd2} : s = 176;
	{8'd110,8'd3} : s = 330;
	{8'd110,8'd4} : s = 329;
	{8'd110,8'd5} : s = 440;
	{8'd110,8'd6} : s = 326;
	{8'd110,8'd7} : s = 436;
	{8'd110,8'd8} : s = 434;
	{8'd110,8'd9} : s = 497;
	{8'd110,8'd10} : s = 325;
	{8'd110,8'd11} : s = 433;
	{8'd110,8'd12} : s = 428;
	{8'd110,8'd13} : s = 492;
	{8'd110,8'd14} : s = 426;
	{8'd110,8'd15} : s = 490;
	{8'd110,8'd16} : s = 489;
	{8'd110,8'd17} : s = 508;
	{8'd110,8'd18} : s = 2;
	{8'd110,8'd19} : s = 48;
	{8'd110,8'd20} : s = 40;
	{8'd110,8'd21} : s = 168;
	{8'd110,8'd22} : s = 36;
	{8'd110,8'd23} : s = 164;
	{8'd110,8'd24} : s = 162;
	{8'd110,8'd25} : s = 323;
	{8'd110,8'd26} : s = 34;
	{8'd110,8'd27} : s = 161;
	{8'd110,8'd28} : s = 152;
	{8'd110,8'd29} : s = 312;
	{8'd110,8'd30} : s = 148;
	{8'd110,8'd31} : s = 308;
	{8'd110,8'd32} : s = 306;
	{8'd110,8'd33} : s = 425;
	{8'd110,8'd34} : s = 33;
	{8'd110,8'd35} : s = 146;
	{8'd110,8'd36} : s = 145;
	{8'd110,8'd37} : s = 305;
	{8'd110,8'd38} : s = 140;
	{8'd110,8'd39} : s = 300;
	{8'd110,8'd40} : s = 298;
	{8'd110,8'd41} : s = 422;
	{8'd110,8'd42} : s = 138;
	{8'd110,8'd43} : s = 297;
	{8'd110,8'd44} : s = 294;
	{8'd110,8'd45} : s = 421;
	{8'd110,8'd46} : s = 293;
	{8'd110,8'd47} : s = 419;
	{8'd110,8'd48} : s = 412;
	{8'd110,8'd49} : s = 486;
	{8'd110,8'd50} : s = 24;
	{8'd110,8'd51} : s = 137;
	{8'd110,8'd52} : s = 134;
	{8'd110,8'd53} : s = 291;
	{8'd110,8'd54} : s = 133;
	{8'd110,8'd55} : s = 284;
	{8'd110,8'd56} : s = 282;
	{8'd110,8'd57} : s = 410;
	{8'd110,8'd58} : s = 131;
	{8'd110,8'd59} : s = 281;
	{8'd110,8'd60} : s = 278;
	{8'd110,8'd61} : s = 409;
	{8'd110,8'd62} : s = 277;
	{8'd110,8'd63} : s = 406;
	{8'd110,8'd64} : s = 405;
	{8'd110,8'd65} : s = 485;
	{8'd110,8'd66} : s = 112;
	{8'd110,8'd67} : s = 275;
	{8'd110,8'd68} : s = 270;
	{8'd110,8'd69} : s = 403;
	{8'd110,8'd70} : s = 269;
	{8'd110,8'd71} : s = 398;
	{8'd110,8'd72} : s = 397;
	{8'd110,8'd73} : s = 483;
	{8'd110,8'd74} : s = 267;
	{8'd110,8'd75} : s = 395;
	{8'd110,8'd76} : s = 391;
	{8'd110,8'd77} : s = 476;
	{8'd110,8'd78} : s = 376;
	{8'd110,8'd79} : s = 474;
	{8'd110,8'd80} : s = 473;
	{8'd110,8'd81} : s = 506;
	{8'd110,8'd82} : s = 20;
	{8'd110,8'd83} : s = 104;
	{8'd110,8'd84} : s = 100;
	{8'd110,8'd85} : s = 263;
	{8'd110,8'd86} : s = 98;
	{8'd110,8'd87} : s = 240;
	{8'd110,8'd88} : s = 232;
	{8'd110,8'd89} : s = 372;
	{8'd110,8'd90} : s = 97;
	{8'd110,8'd91} : s = 228;
	{8'd110,8'd92} : s = 226;
	{8'd110,8'd93} : s = 370;
	{8'd110,8'd94} : s = 225;
	{8'd110,8'd95} : s = 369;
	{8'd110,8'd96} : s = 364;
	{8'd110,8'd97} : s = 470;
	{8'd110,8'd98} : s = 88;
	{8'd110,8'd99} : s = 216;
	{8'd110,8'd100} : s = 212;
	{8'd110,8'd101} : s = 362;
	{8'd110,8'd102} : s = 210;
	{8'd110,8'd103} : s = 361;
	{8'd110,8'd104} : s = 358;
	{8'd110,8'd105} : s = 469;
	{8'd110,8'd106} : s = 209;
	{8'd110,8'd107} : s = 357;
	{8'd110,8'd108} : s = 355;
	{8'd110,8'd109} : s = 467;
	{8'd110,8'd110} : s = 348;
	{8'd110,8'd111} : s = 462;
	{8'd110,8'd112} : s = 461;
	{8'd110,8'd113} : s = 505;
	{8'd110,8'd114} : s = 84;
	{8'd110,8'd115} : s = 204;
	{8'd110,8'd116} : s = 202;
	{8'd110,8'd117} : s = 346;
	{8'd110,8'd118} : s = 201;
	{8'd110,8'd119} : s = 345;
	{8'd110,8'd120} : s = 342;
	{8'd110,8'd121} : s = 459;
	{8'd110,8'd122} : s = 198;
	{8'd110,8'd123} : s = 341;
	{8'd110,8'd124} : s = 339;
	{8'd110,8'd125} : s = 455;
	{8'd110,8'd126} : s = 334;
	{8'd110,8'd127} : s = 444;
	{8'd110,8'd128} : s = 442;
	{8'd110,8'd129} : s = 502;
	{8'd110,8'd130} : s = 197;
	{8'd110,8'd131} : s = 333;
	{8'd110,8'd132} : s = 331;
	{8'd110,8'd133} : s = 441;
	{8'd110,8'd134} : s = 327;
	{8'd110,8'd135} : s = 438;
	{8'd110,8'd136} : s = 437;
	{8'd110,8'd137} : s = 501;
	{8'd110,8'd138} : s = 316;
	{8'd110,8'd139} : s = 435;
	{8'd110,8'd140} : s = 430;
	{8'd110,8'd141} : s = 499;
	{8'd110,8'd142} : s = 429;
	{8'd110,8'd143} : s = 494;
	{8'd110,8'd144} : s = 493;
	{8'd110,8'd145} : s = 510;
	{8'd110,8'd146} : s = 1;
	{8'd110,8'd147} : s = 18;
	{8'd110,8'd148} : s = 17;
	{8'd110,8'd149} : s = 82;
	{8'd110,8'd150} : s = 12;
	{8'd110,8'd151} : s = 81;
	{8'd110,8'd152} : s = 76;
	{8'd110,8'd153} : s = 195;
	{8'd110,8'd154} : s = 10;
	{8'd110,8'd155} : s = 74;
	{8'd110,8'd156} : s = 73;
	{8'd110,8'd157} : s = 184;
	{8'd110,8'd158} : s = 70;
	{8'd110,8'd159} : s = 180;
	{8'd110,8'd160} : s = 178;
	{8'd110,8'd161} : s = 314;
	{8'd110,8'd162} : s = 9;
	{8'd110,8'd163} : s = 69;
	{8'd110,8'd164} : s = 67;
	{8'd110,8'd165} : s = 177;
	{8'd110,8'd166} : s = 56;
	{8'd110,8'd167} : s = 172;
	{8'd110,8'd168} : s = 170;
	{8'd110,8'd169} : s = 313;
	{8'd110,8'd170} : s = 52;
	{8'd110,8'd171} : s = 169;
	{8'd110,8'd172} : s = 166;
	{8'd110,8'd173} : s = 310;
	{8'd110,8'd174} : s = 165;
	{8'd110,8'd175} : s = 309;
	{8'd110,8'd176} : s = 307;
	{8'd110,8'd177} : s = 427;
	{8'd110,8'd178} : s = 6;
	{8'd110,8'd179} : s = 50;
	{8'd110,8'd180} : s = 49;
	{8'd110,8'd181} : s = 163;
	{8'd110,8'd182} : s = 44;
	{8'd110,8'd183} : s = 156;
	{8'd110,8'd184} : s = 154;
	{8'd110,8'd185} : s = 302;
	{8'd110,8'd186} : s = 42;
	{8'd110,8'd187} : s = 153;
	{8'd110,8'd188} : s = 150;
	{8'd110,8'd189} : s = 301;
	{8'd110,8'd190} : s = 149;
	{8'd110,8'd191} : s = 299;
	{8'd110,8'd192} : s = 295;
	{8'd110,8'd193} : s = 423;
	{8'd110,8'd194} : s = 41;
	{8'd110,8'd195} : s = 147;
	{8'd110,8'd196} : s = 142;
	{8'd110,8'd197} : s = 286;
	{8'd110,8'd198} : s = 141;
	{8'd110,8'd199} : s = 285;
	{8'd110,8'd200} : s = 283;
	{8'd110,8'd201} : s = 414;
	{8'd110,8'd202} : s = 139;
	{8'd110,8'd203} : s = 279;
	{8'd110,8'd204} : s = 271;
	{8'd110,8'd205} : s = 413;
	{8'd110,8'd206} : s = 248;
	{8'd110,8'd207} : s = 411;
	{8'd110,8'd208} : s = 407;
	{8'd110,8'd209} : s = 491;
	{8'd110,8'd210} : s = 5;
	{8'd110,8'd211} : s = 38;
	{8'd110,8'd212} : s = 37;
	{8'd110,8'd213} : s = 135;
	{8'd110,8'd214} : s = 35;
	{8'd110,8'd215} : s = 120;
	{8'd110,8'd216} : s = 116;
	{8'd110,8'd217} : s = 244;
	{8'd110,8'd218} : s = 28;
	{8'd110,8'd219} : s = 114;
	{8'd110,8'd220} : s = 113;
	{8'd110,8'd221} : s = 242;
	{8'd110,8'd222} : s = 108;
	{8'd110,8'd223} : s = 241;
	{8'd110,8'd224} : s = 236;
	{8'd110,8'd225} : s = 399;
	{8'd110,8'd226} : s = 26;
	{8'd110,8'd227} : s = 106;
	{8'd110,8'd228} : s = 105;
	{8'd110,8'd229} : s = 234;
	{8'd110,8'd230} : s = 102;
	{8'd110,8'd231} : s = 233;
	{8'd110,8'd232} : s = 230;
	{8'd110,8'd233} : s = 380;
	{8'd110,8'd234} : s = 101;
	{8'd110,8'd235} : s = 229;
	{8'd110,8'd236} : s = 227;
	{8'd110,8'd237} : s = 378;
	{8'd110,8'd238} : s = 220;
	{8'd110,8'd239} : s = 377;
	{8'd110,8'd240} : s = 374;
	{8'd110,8'd241} : s = 487;
	{8'd110,8'd242} : s = 25;
	{8'd110,8'd243} : s = 99;
	{8'd110,8'd244} : s = 92;
	{8'd110,8'd245} : s = 218;
	{8'd110,8'd246} : s = 90;
	{8'd110,8'd247} : s = 217;
	{8'd110,8'd248} : s = 214;
	{8'd110,8'd249} : s = 373;
	{8'd110,8'd250} : s = 89;
	{8'd110,8'd251} : s = 213;
	{8'd110,8'd252} : s = 211;
	{8'd110,8'd253} : s = 371;
	{8'd110,8'd254} : s = 206;
	{8'd110,8'd255} : s = 366;
	{8'd111,8'd0} : s = 498;
	{8'd111,8'd1} : s = 176;
	{8'd111,8'd2} : s = 330;
	{8'd111,8'd3} : s = 329;
	{8'd111,8'd4} : s = 440;
	{8'd111,8'd5} : s = 326;
	{8'd111,8'd6} : s = 436;
	{8'd111,8'd7} : s = 434;
	{8'd111,8'd8} : s = 497;
	{8'd111,8'd9} : s = 325;
	{8'd111,8'd10} : s = 433;
	{8'd111,8'd11} : s = 428;
	{8'd111,8'd12} : s = 492;
	{8'd111,8'd13} : s = 426;
	{8'd111,8'd14} : s = 490;
	{8'd111,8'd15} : s = 489;
	{8'd111,8'd16} : s = 508;
	{8'd111,8'd17} : s = 2;
	{8'd111,8'd18} : s = 48;
	{8'd111,8'd19} : s = 40;
	{8'd111,8'd20} : s = 168;
	{8'd111,8'd21} : s = 36;
	{8'd111,8'd22} : s = 164;
	{8'd111,8'd23} : s = 162;
	{8'd111,8'd24} : s = 323;
	{8'd111,8'd25} : s = 34;
	{8'd111,8'd26} : s = 161;
	{8'd111,8'd27} : s = 152;
	{8'd111,8'd28} : s = 312;
	{8'd111,8'd29} : s = 148;
	{8'd111,8'd30} : s = 308;
	{8'd111,8'd31} : s = 306;
	{8'd111,8'd32} : s = 425;
	{8'd111,8'd33} : s = 33;
	{8'd111,8'd34} : s = 146;
	{8'd111,8'd35} : s = 145;
	{8'd111,8'd36} : s = 305;
	{8'd111,8'd37} : s = 140;
	{8'd111,8'd38} : s = 300;
	{8'd111,8'd39} : s = 298;
	{8'd111,8'd40} : s = 422;
	{8'd111,8'd41} : s = 138;
	{8'd111,8'd42} : s = 297;
	{8'd111,8'd43} : s = 294;
	{8'd111,8'd44} : s = 421;
	{8'd111,8'd45} : s = 293;
	{8'd111,8'd46} : s = 419;
	{8'd111,8'd47} : s = 412;
	{8'd111,8'd48} : s = 486;
	{8'd111,8'd49} : s = 24;
	{8'd111,8'd50} : s = 137;
	{8'd111,8'd51} : s = 134;
	{8'd111,8'd52} : s = 291;
	{8'd111,8'd53} : s = 133;
	{8'd111,8'd54} : s = 284;
	{8'd111,8'd55} : s = 282;
	{8'd111,8'd56} : s = 410;
	{8'd111,8'd57} : s = 131;
	{8'd111,8'd58} : s = 281;
	{8'd111,8'd59} : s = 278;
	{8'd111,8'd60} : s = 409;
	{8'd111,8'd61} : s = 277;
	{8'd111,8'd62} : s = 406;
	{8'd111,8'd63} : s = 405;
	{8'd111,8'd64} : s = 485;
	{8'd111,8'd65} : s = 112;
	{8'd111,8'd66} : s = 275;
	{8'd111,8'd67} : s = 270;
	{8'd111,8'd68} : s = 403;
	{8'd111,8'd69} : s = 269;
	{8'd111,8'd70} : s = 398;
	{8'd111,8'd71} : s = 397;
	{8'd111,8'd72} : s = 483;
	{8'd111,8'd73} : s = 267;
	{8'd111,8'd74} : s = 395;
	{8'd111,8'd75} : s = 391;
	{8'd111,8'd76} : s = 476;
	{8'd111,8'd77} : s = 376;
	{8'd111,8'd78} : s = 474;
	{8'd111,8'd79} : s = 473;
	{8'd111,8'd80} : s = 506;
	{8'd111,8'd81} : s = 20;
	{8'd111,8'd82} : s = 104;
	{8'd111,8'd83} : s = 100;
	{8'd111,8'd84} : s = 263;
	{8'd111,8'd85} : s = 98;
	{8'd111,8'd86} : s = 240;
	{8'd111,8'd87} : s = 232;
	{8'd111,8'd88} : s = 372;
	{8'd111,8'd89} : s = 97;
	{8'd111,8'd90} : s = 228;
	{8'd111,8'd91} : s = 226;
	{8'd111,8'd92} : s = 370;
	{8'd111,8'd93} : s = 225;
	{8'd111,8'd94} : s = 369;
	{8'd111,8'd95} : s = 364;
	{8'd111,8'd96} : s = 470;
	{8'd111,8'd97} : s = 88;
	{8'd111,8'd98} : s = 216;
	{8'd111,8'd99} : s = 212;
	{8'd111,8'd100} : s = 362;
	{8'd111,8'd101} : s = 210;
	{8'd111,8'd102} : s = 361;
	{8'd111,8'd103} : s = 358;
	{8'd111,8'd104} : s = 469;
	{8'd111,8'd105} : s = 209;
	{8'd111,8'd106} : s = 357;
	{8'd111,8'd107} : s = 355;
	{8'd111,8'd108} : s = 467;
	{8'd111,8'd109} : s = 348;
	{8'd111,8'd110} : s = 462;
	{8'd111,8'd111} : s = 461;
	{8'd111,8'd112} : s = 505;
	{8'd111,8'd113} : s = 84;
	{8'd111,8'd114} : s = 204;
	{8'd111,8'd115} : s = 202;
	{8'd111,8'd116} : s = 346;
	{8'd111,8'd117} : s = 201;
	{8'd111,8'd118} : s = 345;
	{8'd111,8'd119} : s = 342;
	{8'd111,8'd120} : s = 459;
	{8'd111,8'd121} : s = 198;
	{8'd111,8'd122} : s = 341;
	{8'd111,8'd123} : s = 339;
	{8'd111,8'd124} : s = 455;
	{8'd111,8'd125} : s = 334;
	{8'd111,8'd126} : s = 444;
	{8'd111,8'd127} : s = 442;
	{8'd111,8'd128} : s = 502;
	{8'd111,8'd129} : s = 197;
	{8'd111,8'd130} : s = 333;
	{8'd111,8'd131} : s = 331;
	{8'd111,8'd132} : s = 441;
	{8'd111,8'd133} : s = 327;
	{8'd111,8'd134} : s = 438;
	{8'd111,8'd135} : s = 437;
	{8'd111,8'd136} : s = 501;
	{8'd111,8'd137} : s = 316;
	{8'd111,8'd138} : s = 435;
	{8'd111,8'd139} : s = 430;
	{8'd111,8'd140} : s = 499;
	{8'd111,8'd141} : s = 429;
	{8'd111,8'd142} : s = 494;
	{8'd111,8'd143} : s = 493;
	{8'd111,8'd144} : s = 510;
	{8'd111,8'd145} : s = 1;
	{8'd111,8'd146} : s = 18;
	{8'd111,8'd147} : s = 17;
	{8'd111,8'd148} : s = 82;
	{8'd111,8'd149} : s = 12;
	{8'd111,8'd150} : s = 81;
	{8'd111,8'd151} : s = 76;
	{8'd111,8'd152} : s = 195;
	{8'd111,8'd153} : s = 10;
	{8'd111,8'd154} : s = 74;
	{8'd111,8'd155} : s = 73;
	{8'd111,8'd156} : s = 184;
	{8'd111,8'd157} : s = 70;
	{8'd111,8'd158} : s = 180;
	{8'd111,8'd159} : s = 178;
	{8'd111,8'd160} : s = 314;
	{8'd111,8'd161} : s = 9;
	{8'd111,8'd162} : s = 69;
	{8'd111,8'd163} : s = 67;
	{8'd111,8'd164} : s = 177;
	{8'd111,8'd165} : s = 56;
	{8'd111,8'd166} : s = 172;
	{8'd111,8'd167} : s = 170;
	{8'd111,8'd168} : s = 313;
	{8'd111,8'd169} : s = 52;
	{8'd111,8'd170} : s = 169;
	{8'd111,8'd171} : s = 166;
	{8'd111,8'd172} : s = 310;
	{8'd111,8'd173} : s = 165;
	{8'd111,8'd174} : s = 309;
	{8'd111,8'd175} : s = 307;
	{8'd111,8'd176} : s = 427;
	{8'd111,8'd177} : s = 6;
	{8'd111,8'd178} : s = 50;
	{8'd111,8'd179} : s = 49;
	{8'd111,8'd180} : s = 163;
	{8'd111,8'd181} : s = 44;
	{8'd111,8'd182} : s = 156;
	{8'd111,8'd183} : s = 154;
	{8'd111,8'd184} : s = 302;
	{8'd111,8'd185} : s = 42;
	{8'd111,8'd186} : s = 153;
	{8'd111,8'd187} : s = 150;
	{8'd111,8'd188} : s = 301;
	{8'd111,8'd189} : s = 149;
	{8'd111,8'd190} : s = 299;
	{8'd111,8'd191} : s = 295;
	{8'd111,8'd192} : s = 423;
	{8'd111,8'd193} : s = 41;
	{8'd111,8'd194} : s = 147;
	{8'd111,8'd195} : s = 142;
	{8'd111,8'd196} : s = 286;
	{8'd111,8'd197} : s = 141;
	{8'd111,8'd198} : s = 285;
	{8'd111,8'd199} : s = 283;
	{8'd111,8'd200} : s = 414;
	{8'd111,8'd201} : s = 139;
	{8'd111,8'd202} : s = 279;
	{8'd111,8'd203} : s = 271;
	{8'd111,8'd204} : s = 413;
	{8'd111,8'd205} : s = 248;
	{8'd111,8'd206} : s = 411;
	{8'd111,8'd207} : s = 407;
	{8'd111,8'd208} : s = 491;
	{8'd111,8'd209} : s = 5;
	{8'd111,8'd210} : s = 38;
	{8'd111,8'd211} : s = 37;
	{8'd111,8'd212} : s = 135;
	{8'd111,8'd213} : s = 35;
	{8'd111,8'd214} : s = 120;
	{8'd111,8'd215} : s = 116;
	{8'd111,8'd216} : s = 244;
	{8'd111,8'd217} : s = 28;
	{8'd111,8'd218} : s = 114;
	{8'd111,8'd219} : s = 113;
	{8'd111,8'd220} : s = 242;
	{8'd111,8'd221} : s = 108;
	{8'd111,8'd222} : s = 241;
	{8'd111,8'd223} : s = 236;
	{8'd111,8'd224} : s = 399;
	{8'd111,8'd225} : s = 26;
	{8'd111,8'd226} : s = 106;
	{8'd111,8'd227} : s = 105;
	{8'd111,8'd228} : s = 234;
	{8'd111,8'd229} : s = 102;
	{8'd111,8'd230} : s = 233;
	{8'd111,8'd231} : s = 230;
	{8'd111,8'd232} : s = 380;
	{8'd111,8'd233} : s = 101;
	{8'd111,8'd234} : s = 229;
	{8'd111,8'd235} : s = 227;
	{8'd111,8'd236} : s = 378;
	{8'd111,8'd237} : s = 220;
	{8'd111,8'd238} : s = 377;
	{8'd111,8'd239} : s = 374;
	{8'd111,8'd240} : s = 487;
	{8'd111,8'd241} : s = 25;
	{8'd111,8'd242} : s = 99;
	{8'd111,8'd243} : s = 92;
	{8'd111,8'd244} : s = 218;
	{8'd111,8'd245} : s = 90;
	{8'd111,8'd246} : s = 217;
	{8'd111,8'd247} : s = 214;
	{8'd111,8'd248} : s = 373;
	{8'd111,8'd249} : s = 89;
	{8'd111,8'd250} : s = 213;
	{8'd111,8'd251} : s = 211;
	{8'd111,8'd252} : s = 371;
	{8'd111,8'd253} : s = 206;
	{8'd111,8'd254} : s = 366;
	{8'd111,8'd255} : s = 365;
	{8'd112,8'd0} : s = 176;
	{8'd112,8'd1} : s = 330;
	{8'd112,8'd2} : s = 329;
	{8'd112,8'd3} : s = 440;
	{8'd112,8'd4} : s = 326;
	{8'd112,8'd5} : s = 436;
	{8'd112,8'd6} : s = 434;
	{8'd112,8'd7} : s = 497;
	{8'd112,8'd8} : s = 325;
	{8'd112,8'd9} : s = 433;
	{8'd112,8'd10} : s = 428;
	{8'd112,8'd11} : s = 492;
	{8'd112,8'd12} : s = 426;
	{8'd112,8'd13} : s = 490;
	{8'd112,8'd14} : s = 489;
	{8'd112,8'd15} : s = 508;
	{8'd112,8'd16} : s = 2;
	{8'd112,8'd17} : s = 48;
	{8'd112,8'd18} : s = 40;
	{8'd112,8'd19} : s = 168;
	{8'd112,8'd20} : s = 36;
	{8'd112,8'd21} : s = 164;
	{8'd112,8'd22} : s = 162;
	{8'd112,8'd23} : s = 323;
	{8'd112,8'd24} : s = 34;
	{8'd112,8'd25} : s = 161;
	{8'd112,8'd26} : s = 152;
	{8'd112,8'd27} : s = 312;
	{8'd112,8'd28} : s = 148;
	{8'd112,8'd29} : s = 308;
	{8'd112,8'd30} : s = 306;
	{8'd112,8'd31} : s = 425;
	{8'd112,8'd32} : s = 33;
	{8'd112,8'd33} : s = 146;
	{8'd112,8'd34} : s = 145;
	{8'd112,8'd35} : s = 305;
	{8'd112,8'd36} : s = 140;
	{8'd112,8'd37} : s = 300;
	{8'd112,8'd38} : s = 298;
	{8'd112,8'd39} : s = 422;
	{8'd112,8'd40} : s = 138;
	{8'd112,8'd41} : s = 297;
	{8'd112,8'd42} : s = 294;
	{8'd112,8'd43} : s = 421;
	{8'd112,8'd44} : s = 293;
	{8'd112,8'd45} : s = 419;
	{8'd112,8'd46} : s = 412;
	{8'd112,8'd47} : s = 486;
	{8'd112,8'd48} : s = 24;
	{8'd112,8'd49} : s = 137;
	{8'd112,8'd50} : s = 134;
	{8'd112,8'd51} : s = 291;
	{8'd112,8'd52} : s = 133;
	{8'd112,8'd53} : s = 284;
	{8'd112,8'd54} : s = 282;
	{8'd112,8'd55} : s = 410;
	{8'd112,8'd56} : s = 131;
	{8'd112,8'd57} : s = 281;
	{8'd112,8'd58} : s = 278;
	{8'd112,8'd59} : s = 409;
	{8'd112,8'd60} : s = 277;
	{8'd112,8'd61} : s = 406;
	{8'd112,8'd62} : s = 405;
	{8'd112,8'd63} : s = 485;
	{8'd112,8'd64} : s = 112;
	{8'd112,8'd65} : s = 275;
	{8'd112,8'd66} : s = 270;
	{8'd112,8'd67} : s = 403;
	{8'd112,8'd68} : s = 269;
	{8'd112,8'd69} : s = 398;
	{8'd112,8'd70} : s = 397;
	{8'd112,8'd71} : s = 483;
	{8'd112,8'd72} : s = 267;
	{8'd112,8'd73} : s = 395;
	{8'd112,8'd74} : s = 391;
	{8'd112,8'd75} : s = 476;
	{8'd112,8'd76} : s = 376;
	{8'd112,8'd77} : s = 474;
	{8'd112,8'd78} : s = 473;
	{8'd112,8'd79} : s = 506;
	{8'd112,8'd80} : s = 20;
	{8'd112,8'd81} : s = 104;
	{8'd112,8'd82} : s = 100;
	{8'd112,8'd83} : s = 263;
	{8'd112,8'd84} : s = 98;
	{8'd112,8'd85} : s = 240;
	{8'd112,8'd86} : s = 232;
	{8'd112,8'd87} : s = 372;
	{8'd112,8'd88} : s = 97;
	{8'd112,8'd89} : s = 228;
	{8'd112,8'd90} : s = 226;
	{8'd112,8'd91} : s = 370;
	{8'd112,8'd92} : s = 225;
	{8'd112,8'd93} : s = 369;
	{8'd112,8'd94} : s = 364;
	{8'd112,8'd95} : s = 470;
	{8'd112,8'd96} : s = 88;
	{8'd112,8'd97} : s = 216;
	{8'd112,8'd98} : s = 212;
	{8'd112,8'd99} : s = 362;
	{8'd112,8'd100} : s = 210;
	{8'd112,8'd101} : s = 361;
	{8'd112,8'd102} : s = 358;
	{8'd112,8'd103} : s = 469;
	{8'd112,8'd104} : s = 209;
	{8'd112,8'd105} : s = 357;
	{8'd112,8'd106} : s = 355;
	{8'd112,8'd107} : s = 467;
	{8'd112,8'd108} : s = 348;
	{8'd112,8'd109} : s = 462;
	{8'd112,8'd110} : s = 461;
	{8'd112,8'd111} : s = 505;
	{8'd112,8'd112} : s = 84;
	{8'd112,8'd113} : s = 204;
	{8'd112,8'd114} : s = 202;
	{8'd112,8'd115} : s = 346;
	{8'd112,8'd116} : s = 201;
	{8'd112,8'd117} : s = 345;
	{8'd112,8'd118} : s = 342;
	{8'd112,8'd119} : s = 459;
	{8'd112,8'd120} : s = 198;
	{8'd112,8'd121} : s = 341;
	{8'd112,8'd122} : s = 339;
	{8'd112,8'd123} : s = 455;
	{8'd112,8'd124} : s = 334;
	{8'd112,8'd125} : s = 444;
	{8'd112,8'd126} : s = 442;
	{8'd112,8'd127} : s = 502;
	{8'd112,8'd128} : s = 197;
	{8'd112,8'd129} : s = 333;
	{8'd112,8'd130} : s = 331;
	{8'd112,8'd131} : s = 441;
	{8'd112,8'd132} : s = 327;
	{8'd112,8'd133} : s = 438;
	{8'd112,8'd134} : s = 437;
	{8'd112,8'd135} : s = 501;
	{8'd112,8'd136} : s = 316;
	{8'd112,8'd137} : s = 435;
	{8'd112,8'd138} : s = 430;
	{8'd112,8'd139} : s = 499;
	{8'd112,8'd140} : s = 429;
	{8'd112,8'd141} : s = 494;
	{8'd112,8'd142} : s = 493;
	{8'd112,8'd143} : s = 510;
	{8'd112,8'd144} : s = 1;
	{8'd112,8'd145} : s = 18;
	{8'd112,8'd146} : s = 17;
	{8'd112,8'd147} : s = 82;
	{8'd112,8'd148} : s = 12;
	{8'd112,8'd149} : s = 81;
	{8'd112,8'd150} : s = 76;
	{8'd112,8'd151} : s = 195;
	{8'd112,8'd152} : s = 10;
	{8'd112,8'd153} : s = 74;
	{8'd112,8'd154} : s = 73;
	{8'd112,8'd155} : s = 184;
	{8'd112,8'd156} : s = 70;
	{8'd112,8'd157} : s = 180;
	{8'd112,8'd158} : s = 178;
	{8'd112,8'd159} : s = 314;
	{8'd112,8'd160} : s = 9;
	{8'd112,8'd161} : s = 69;
	{8'd112,8'd162} : s = 67;
	{8'd112,8'd163} : s = 177;
	{8'd112,8'd164} : s = 56;
	{8'd112,8'd165} : s = 172;
	{8'd112,8'd166} : s = 170;
	{8'd112,8'd167} : s = 313;
	{8'd112,8'd168} : s = 52;
	{8'd112,8'd169} : s = 169;
	{8'd112,8'd170} : s = 166;
	{8'd112,8'd171} : s = 310;
	{8'd112,8'd172} : s = 165;
	{8'd112,8'd173} : s = 309;
	{8'd112,8'd174} : s = 307;
	{8'd112,8'd175} : s = 427;
	{8'd112,8'd176} : s = 6;
	{8'd112,8'd177} : s = 50;
	{8'd112,8'd178} : s = 49;
	{8'd112,8'd179} : s = 163;
	{8'd112,8'd180} : s = 44;
	{8'd112,8'd181} : s = 156;
	{8'd112,8'd182} : s = 154;
	{8'd112,8'd183} : s = 302;
	{8'd112,8'd184} : s = 42;
	{8'd112,8'd185} : s = 153;
	{8'd112,8'd186} : s = 150;
	{8'd112,8'd187} : s = 301;
	{8'd112,8'd188} : s = 149;
	{8'd112,8'd189} : s = 299;
	{8'd112,8'd190} : s = 295;
	{8'd112,8'd191} : s = 423;
	{8'd112,8'd192} : s = 41;
	{8'd112,8'd193} : s = 147;
	{8'd112,8'd194} : s = 142;
	{8'd112,8'd195} : s = 286;
	{8'd112,8'd196} : s = 141;
	{8'd112,8'd197} : s = 285;
	{8'd112,8'd198} : s = 283;
	{8'd112,8'd199} : s = 414;
	{8'd112,8'd200} : s = 139;
	{8'd112,8'd201} : s = 279;
	{8'd112,8'd202} : s = 271;
	{8'd112,8'd203} : s = 413;
	{8'd112,8'd204} : s = 248;
	{8'd112,8'd205} : s = 411;
	{8'd112,8'd206} : s = 407;
	{8'd112,8'd207} : s = 491;
	{8'd112,8'd208} : s = 5;
	{8'd112,8'd209} : s = 38;
	{8'd112,8'd210} : s = 37;
	{8'd112,8'd211} : s = 135;
	{8'd112,8'd212} : s = 35;
	{8'd112,8'd213} : s = 120;
	{8'd112,8'd214} : s = 116;
	{8'd112,8'd215} : s = 244;
	{8'd112,8'd216} : s = 28;
	{8'd112,8'd217} : s = 114;
	{8'd112,8'd218} : s = 113;
	{8'd112,8'd219} : s = 242;
	{8'd112,8'd220} : s = 108;
	{8'd112,8'd221} : s = 241;
	{8'd112,8'd222} : s = 236;
	{8'd112,8'd223} : s = 399;
	{8'd112,8'd224} : s = 26;
	{8'd112,8'd225} : s = 106;
	{8'd112,8'd226} : s = 105;
	{8'd112,8'd227} : s = 234;
	{8'd112,8'd228} : s = 102;
	{8'd112,8'd229} : s = 233;
	{8'd112,8'd230} : s = 230;
	{8'd112,8'd231} : s = 380;
	{8'd112,8'd232} : s = 101;
	{8'd112,8'd233} : s = 229;
	{8'd112,8'd234} : s = 227;
	{8'd112,8'd235} : s = 378;
	{8'd112,8'd236} : s = 220;
	{8'd112,8'd237} : s = 377;
	{8'd112,8'd238} : s = 374;
	{8'd112,8'd239} : s = 487;
	{8'd112,8'd240} : s = 25;
	{8'd112,8'd241} : s = 99;
	{8'd112,8'd242} : s = 92;
	{8'd112,8'd243} : s = 218;
	{8'd112,8'd244} : s = 90;
	{8'd112,8'd245} : s = 217;
	{8'd112,8'd246} : s = 214;
	{8'd112,8'd247} : s = 373;
	{8'd112,8'd248} : s = 89;
	{8'd112,8'd249} : s = 213;
	{8'd112,8'd250} : s = 211;
	{8'd112,8'd251} : s = 371;
	{8'd112,8'd252} : s = 206;
	{8'd112,8'd253} : s = 366;
	{8'd112,8'd254} : s = 365;
	{8'd112,8'd255} : s = 478;
	{8'd113,8'd0} : s = 330;
	{8'd113,8'd1} : s = 329;
	{8'd113,8'd2} : s = 440;
	{8'd113,8'd3} : s = 326;
	{8'd113,8'd4} : s = 436;
	{8'd113,8'd5} : s = 434;
	{8'd113,8'd6} : s = 497;
	{8'd113,8'd7} : s = 325;
	{8'd113,8'd8} : s = 433;
	{8'd113,8'd9} : s = 428;
	{8'd113,8'd10} : s = 492;
	{8'd113,8'd11} : s = 426;
	{8'd113,8'd12} : s = 490;
	{8'd113,8'd13} : s = 489;
	{8'd113,8'd14} : s = 508;
	{8'd113,8'd15} : s = 2;
	{8'd113,8'd16} : s = 48;
	{8'd113,8'd17} : s = 40;
	{8'd113,8'd18} : s = 168;
	{8'd113,8'd19} : s = 36;
	{8'd113,8'd20} : s = 164;
	{8'd113,8'd21} : s = 162;
	{8'd113,8'd22} : s = 323;
	{8'd113,8'd23} : s = 34;
	{8'd113,8'd24} : s = 161;
	{8'd113,8'd25} : s = 152;
	{8'd113,8'd26} : s = 312;
	{8'd113,8'd27} : s = 148;
	{8'd113,8'd28} : s = 308;
	{8'd113,8'd29} : s = 306;
	{8'd113,8'd30} : s = 425;
	{8'd113,8'd31} : s = 33;
	{8'd113,8'd32} : s = 146;
	{8'd113,8'd33} : s = 145;
	{8'd113,8'd34} : s = 305;
	{8'd113,8'd35} : s = 140;
	{8'd113,8'd36} : s = 300;
	{8'd113,8'd37} : s = 298;
	{8'd113,8'd38} : s = 422;
	{8'd113,8'd39} : s = 138;
	{8'd113,8'd40} : s = 297;
	{8'd113,8'd41} : s = 294;
	{8'd113,8'd42} : s = 421;
	{8'd113,8'd43} : s = 293;
	{8'd113,8'd44} : s = 419;
	{8'd113,8'd45} : s = 412;
	{8'd113,8'd46} : s = 486;
	{8'd113,8'd47} : s = 24;
	{8'd113,8'd48} : s = 137;
	{8'd113,8'd49} : s = 134;
	{8'd113,8'd50} : s = 291;
	{8'd113,8'd51} : s = 133;
	{8'd113,8'd52} : s = 284;
	{8'd113,8'd53} : s = 282;
	{8'd113,8'd54} : s = 410;
	{8'd113,8'd55} : s = 131;
	{8'd113,8'd56} : s = 281;
	{8'd113,8'd57} : s = 278;
	{8'd113,8'd58} : s = 409;
	{8'd113,8'd59} : s = 277;
	{8'd113,8'd60} : s = 406;
	{8'd113,8'd61} : s = 405;
	{8'd113,8'd62} : s = 485;
	{8'd113,8'd63} : s = 112;
	{8'd113,8'd64} : s = 275;
	{8'd113,8'd65} : s = 270;
	{8'd113,8'd66} : s = 403;
	{8'd113,8'd67} : s = 269;
	{8'd113,8'd68} : s = 398;
	{8'd113,8'd69} : s = 397;
	{8'd113,8'd70} : s = 483;
	{8'd113,8'd71} : s = 267;
	{8'd113,8'd72} : s = 395;
	{8'd113,8'd73} : s = 391;
	{8'd113,8'd74} : s = 476;
	{8'd113,8'd75} : s = 376;
	{8'd113,8'd76} : s = 474;
	{8'd113,8'd77} : s = 473;
	{8'd113,8'd78} : s = 506;
	{8'd113,8'd79} : s = 20;
	{8'd113,8'd80} : s = 104;
	{8'd113,8'd81} : s = 100;
	{8'd113,8'd82} : s = 263;
	{8'd113,8'd83} : s = 98;
	{8'd113,8'd84} : s = 240;
	{8'd113,8'd85} : s = 232;
	{8'd113,8'd86} : s = 372;
	{8'd113,8'd87} : s = 97;
	{8'd113,8'd88} : s = 228;
	{8'd113,8'd89} : s = 226;
	{8'd113,8'd90} : s = 370;
	{8'd113,8'd91} : s = 225;
	{8'd113,8'd92} : s = 369;
	{8'd113,8'd93} : s = 364;
	{8'd113,8'd94} : s = 470;
	{8'd113,8'd95} : s = 88;
	{8'd113,8'd96} : s = 216;
	{8'd113,8'd97} : s = 212;
	{8'd113,8'd98} : s = 362;
	{8'd113,8'd99} : s = 210;
	{8'd113,8'd100} : s = 361;
	{8'd113,8'd101} : s = 358;
	{8'd113,8'd102} : s = 469;
	{8'd113,8'd103} : s = 209;
	{8'd113,8'd104} : s = 357;
	{8'd113,8'd105} : s = 355;
	{8'd113,8'd106} : s = 467;
	{8'd113,8'd107} : s = 348;
	{8'd113,8'd108} : s = 462;
	{8'd113,8'd109} : s = 461;
	{8'd113,8'd110} : s = 505;
	{8'd113,8'd111} : s = 84;
	{8'd113,8'd112} : s = 204;
	{8'd113,8'd113} : s = 202;
	{8'd113,8'd114} : s = 346;
	{8'd113,8'd115} : s = 201;
	{8'd113,8'd116} : s = 345;
	{8'd113,8'd117} : s = 342;
	{8'd113,8'd118} : s = 459;
	{8'd113,8'd119} : s = 198;
	{8'd113,8'd120} : s = 341;
	{8'd113,8'd121} : s = 339;
	{8'd113,8'd122} : s = 455;
	{8'd113,8'd123} : s = 334;
	{8'd113,8'd124} : s = 444;
	{8'd113,8'd125} : s = 442;
	{8'd113,8'd126} : s = 502;
	{8'd113,8'd127} : s = 197;
	{8'd113,8'd128} : s = 333;
	{8'd113,8'd129} : s = 331;
	{8'd113,8'd130} : s = 441;
	{8'd113,8'd131} : s = 327;
	{8'd113,8'd132} : s = 438;
	{8'd113,8'd133} : s = 437;
	{8'd113,8'd134} : s = 501;
	{8'd113,8'd135} : s = 316;
	{8'd113,8'd136} : s = 435;
	{8'd113,8'd137} : s = 430;
	{8'd113,8'd138} : s = 499;
	{8'd113,8'd139} : s = 429;
	{8'd113,8'd140} : s = 494;
	{8'd113,8'd141} : s = 493;
	{8'd113,8'd142} : s = 510;
	{8'd113,8'd143} : s = 1;
	{8'd113,8'd144} : s = 18;
	{8'd113,8'd145} : s = 17;
	{8'd113,8'd146} : s = 82;
	{8'd113,8'd147} : s = 12;
	{8'd113,8'd148} : s = 81;
	{8'd113,8'd149} : s = 76;
	{8'd113,8'd150} : s = 195;
	{8'd113,8'd151} : s = 10;
	{8'd113,8'd152} : s = 74;
	{8'd113,8'd153} : s = 73;
	{8'd113,8'd154} : s = 184;
	{8'd113,8'd155} : s = 70;
	{8'd113,8'd156} : s = 180;
	{8'd113,8'd157} : s = 178;
	{8'd113,8'd158} : s = 314;
	{8'd113,8'd159} : s = 9;
	{8'd113,8'd160} : s = 69;
	{8'd113,8'd161} : s = 67;
	{8'd113,8'd162} : s = 177;
	{8'd113,8'd163} : s = 56;
	{8'd113,8'd164} : s = 172;
	{8'd113,8'd165} : s = 170;
	{8'd113,8'd166} : s = 313;
	{8'd113,8'd167} : s = 52;
	{8'd113,8'd168} : s = 169;
	{8'd113,8'd169} : s = 166;
	{8'd113,8'd170} : s = 310;
	{8'd113,8'd171} : s = 165;
	{8'd113,8'd172} : s = 309;
	{8'd113,8'd173} : s = 307;
	{8'd113,8'd174} : s = 427;
	{8'd113,8'd175} : s = 6;
	{8'd113,8'd176} : s = 50;
	{8'd113,8'd177} : s = 49;
	{8'd113,8'd178} : s = 163;
	{8'd113,8'd179} : s = 44;
	{8'd113,8'd180} : s = 156;
	{8'd113,8'd181} : s = 154;
	{8'd113,8'd182} : s = 302;
	{8'd113,8'd183} : s = 42;
	{8'd113,8'd184} : s = 153;
	{8'd113,8'd185} : s = 150;
	{8'd113,8'd186} : s = 301;
	{8'd113,8'd187} : s = 149;
	{8'd113,8'd188} : s = 299;
	{8'd113,8'd189} : s = 295;
	{8'd113,8'd190} : s = 423;
	{8'd113,8'd191} : s = 41;
	{8'd113,8'd192} : s = 147;
	{8'd113,8'd193} : s = 142;
	{8'd113,8'd194} : s = 286;
	{8'd113,8'd195} : s = 141;
	{8'd113,8'd196} : s = 285;
	{8'd113,8'd197} : s = 283;
	{8'd113,8'd198} : s = 414;
	{8'd113,8'd199} : s = 139;
	{8'd113,8'd200} : s = 279;
	{8'd113,8'd201} : s = 271;
	{8'd113,8'd202} : s = 413;
	{8'd113,8'd203} : s = 248;
	{8'd113,8'd204} : s = 411;
	{8'd113,8'd205} : s = 407;
	{8'd113,8'd206} : s = 491;
	{8'd113,8'd207} : s = 5;
	{8'd113,8'd208} : s = 38;
	{8'd113,8'd209} : s = 37;
	{8'd113,8'd210} : s = 135;
	{8'd113,8'd211} : s = 35;
	{8'd113,8'd212} : s = 120;
	{8'd113,8'd213} : s = 116;
	{8'd113,8'd214} : s = 244;
	{8'd113,8'd215} : s = 28;
	{8'd113,8'd216} : s = 114;
	{8'd113,8'd217} : s = 113;
	{8'd113,8'd218} : s = 242;
	{8'd113,8'd219} : s = 108;
	{8'd113,8'd220} : s = 241;
	{8'd113,8'd221} : s = 236;
	{8'd113,8'd222} : s = 399;
	{8'd113,8'd223} : s = 26;
	{8'd113,8'd224} : s = 106;
	{8'd113,8'd225} : s = 105;
	{8'd113,8'd226} : s = 234;
	{8'd113,8'd227} : s = 102;
	{8'd113,8'd228} : s = 233;
	{8'd113,8'd229} : s = 230;
	{8'd113,8'd230} : s = 380;
	{8'd113,8'd231} : s = 101;
	{8'd113,8'd232} : s = 229;
	{8'd113,8'd233} : s = 227;
	{8'd113,8'd234} : s = 378;
	{8'd113,8'd235} : s = 220;
	{8'd113,8'd236} : s = 377;
	{8'd113,8'd237} : s = 374;
	{8'd113,8'd238} : s = 487;
	{8'd113,8'd239} : s = 25;
	{8'd113,8'd240} : s = 99;
	{8'd113,8'd241} : s = 92;
	{8'd113,8'd242} : s = 218;
	{8'd113,8'd243} : s = 90;
	{8'd113,8'd244} : s = 217;
	{8'd113,8'd245} : s = 214;
	{8'd113,8'd246} : s = 373;
	{8'd113,8'd247} : s = 89;
	{8'd113,8'd248} : s = 213;
	{8'd113,8'd249} : s = 211;
	{8'd113,8'd250} : s = 371;
	{8'd113,8'd251} : s = 206;
	{8'd113,8'd252} : s = 366;
	{8'd113,8'd253} : s = 365;
	{8'd113,8'd254} : s = 478;
	{8'd113,8'd255} : s = 86;
	{8'd114,8'd0} : s = 329;
	{8'd114,8'd1} : s = 440;
	{8'd114,8'd2} : s = 326;
	{8'd114,8'd3} : s = 436;
	{8'd114,8'd4} : s = 434;
	{8'd114,8'd5} : s = 497;
	{8'd114,8'd6} : s = 325;
	{8'd114,8'd7} : s = 433;
	{8'd114,8'd8} : s = 428;
	{8'd114,8'd9} : s = 492;
	{8'd114,8'd10} : s = 426;
	{8'd114,8'd11} : s = 490;
	{8'd114,8'd12} : s = 489;
	{8'd114,8'd13} : s = 508;
	{8'd114,8'd14} : s = 2;
	{8'd114,8'd15} : s = 48;
	{8'd114,8'd16} : s = 40;
	{8'd114,8'd17} : s = 168;
	{8'd114,8'd18} : s = 36;
	{8'd114,8'd19} : s = 164;
	{8'd114,8'd20} : s = 162;
	{8'd114,8'd21} : s = 323;
	{8'd114,8'd22} : s = 34;
	{8'd114,8'd23} : s = 161;
	{8'd114,8'd24} : s = 152;
	{8'd114,8'd25} : s = 312;
	{8'd114,8'd26} : s = 148;
	{8'd114,8'd27} : s = 308;
	{8'd114,8'd28} : s = 306;
	{8'd114,8'd29} : s = 425;
	{8'd114,8'd30} : s = 33;
	{8'd114,8'd31} : s = 146;
	{8'd114,8'd32} : s = 145;
	{8'd114,8'd33} : s = 305;
	{8'd114,8'd34} : s = 140;
	{8'd114,8'd35} : s = 300;
	{8'd114,8'd36} : s = 298;
	{8'd114,8'd37} : s = 422;
	{8'd114,8'd38} : s = 138;
	{8'd114,8'd39} : s = 297;
	{8'd114,8'd40} : s = 294;
	{8'd114,8'd41} : s = 421;
	{8'd114,8'd42} : s = 293;
	{8'd114,8'd43} : s = 419;
	{8'd114,8'd44} : s = 412;
	{8'd114,8'd45} : s = 486;
	{8'd114,8'd46} : s = 24;
	{8'd114,8'd47} : s = 137;
	{8'd114,8'd48} : s = 134;
	{8'd114,8'd49} : s = 291;
	{8'd114,8'd50} : s = 133;
	{8'd114,8'd51} : s = 284;
	{8'd114,8'd52} : s = 282;
	{8'd114,8'd53} : s = 410;
	{8'd114,8'd54} : s = 131;
	{8'd114,8'd55} : s = 281;
	{8'd114,8'd56} : s = 278;
	{8'd114,8'd57} : s = 409;
	{8'd114,8'd58} : s = 277;
	{8'd114,8'd59} : s = 406;
	{8'd114,8'd60} : s = 405;
	{8'd114,8'd61} : s = 485;
	{8'd114,8'd62} : s = 112;
	{8'd114,8'd63} : s = 275;
	{8'd114,8'd64} : s = 270;
	{8'd114,8'd65} : s = 403;
	{8'd114,8'd66} : s = 269;
	{8'd114,8'd67} : s = 398;
	{8'd114,8'd68} : s = 397;
	{8'd114,8'd69} : s = 483;
	{8'd114,8'd70} : s = 267;
	{8'd114,8'd71} : s = 395;
	{8'd114,8'd72} : s = 391;
	{8'd114,8'd73} : s = 476;
	{8'd114,8'd74} : s = 376;
	{8'd114,8'd75} : s = 474;
	{8'd114,8'd76} : s = 473;
	{8'd114,8'd77} : s = 506;
	{8'd114,8'd78} : s = 20;
	{8'd114,8'd79} : s = 104;
	{8'd114,8'd80} : s = 100;
	{8'd114,8'd81} : s = 263;
	{8'd114,8'd82} : s = 98;
	{8'd114,8'd83} : s = 240;
	{8'd114,8'd84} : s = 232;
	{8'd114,8'd85} : s = 372;
	{8'd114,8'd86} : s = 97;
	{8'd114,8'd87} : s = 228;
	{8'd114,8'd88} : s = 226;
	{8'd114,8'd89} : s = 370;
	{8'd114,8'd90} : s = 225;
	{8'd114,8'd91} : s = 369;
	{8'd114,8'd92} : s = 364;
	{8'd114,8'd93} : s = 470;
	{8'd114,8'd94} : s = 88;
	{8'd114,8'd95} : s = 216;
	{8'd114,8'd96} : s = 212;
	{8'd114,8'd97} : s = 362;
	{8'd114,8'd98} : s = 210;
	{8'd114,8'd99} : s = 361;
	{8'd114,8'd100} : s = 358;
	{8'd114,8'd101} : s = 469;
	{8'd114,8'd102} : s = 209;
	{8'd114,8'd103} : s = 357;
	{8'd114,8'd104} : s = 355;
	{8'd114,8'd105} : s = 467;
	{8'd114,8'd106} : s = 348;
	{8'd114,8'd107} : s = 462;
	{8'd114,8'd108} : s = 461;
	{8'd114,8'd109} : s = 505;
	{8'd114,8'd110} : s = 84;
	{8'd114,8'd111} : s = 204;
	{8'd114,8'd112} : s = 202;
	{8'd114,8'd113} : s = 346;
	{8'd114,8'd114} : s = 201;
	{8'd114,8'd115} : s = 345;
	{8'd114,8'd116} : s = 342;
	{8'd114,8'd117} : s = 459;
	{8'd114,8'd118} : s = 198;
	{8'd114,8'd119} : s = 341;
	{8'd114,8'd120} : s = 339;
	{8'd114,8'd121} : s = 455;
	{8'd114,8'd122} : s = 334;
	{8'd114,8'd123} : s = 444;
	{8'd114,8'd124} : s = 442;
	{8'd114,8'd125} : s = 502;
	{8'd114,8'd126} : s = 197;
	{8'd114,8'd127} : s = 333;
	{8'd114,8'd128} : s = 331;
	{8'd114,8'd129} : s = 441;
	{8'd114,8'd130} : s = 327;
	{8'd114,8'd131} : s = 438;
	{8'd114,8'd132} : s = 437;
	{8'd114,8'd133} : s = 501;
	{8'd114,8'd134} : s = 316;
	{8'd114,8'd135} : s = 435;
	{8'd114,8'd136} : s = 430;
	{8'd114,8'd137} : s = 499;
	{8'd114,8'd138} : s = 429;
	{8'd114,8'd139} : s = 494;
	{8'd114,8'd140} : s = 493;
	{8'd114,8'd141} : s = 510;
	{8'd114,8'd142} : s = 1;
	{8'd114,8'd143} : s = 18;
	{8'd114,8'd144} : s = 17;
	{8'd114,8'd145} : s = 82;
	{8'd114,8'd146} : s = 12;
	{8'd114,8'd147} : s = 81;
	{8'd114,8'd148} : s = 76;
	{8'd114,8'd149} : s = 195;
	{8'd114,8'd150} : s = 10;
	{8'd114,8'd151} : s = 74;
	{8'd114,8'd152} : s = 73;
	{8'd114,8'd153} : s = 184;
	{8'd114,8'd154} : s = 70;
	{8'd114,8'd155} : s = 180;
	{8'd114,8'd156} : s = 178;
	{8'd114,8'd157} : s = 314;
	{8'd114,8'd158} : s = 9;
	{8'd114,8'd159} : s = 69;
	{8'd114,8'd160} : s = 67;
	{8'd114,8'd161} : s = 177;
	{8'd114,8'd162} : s = 56;
	{8'd114,8'd163} : s = 172;
	{8'd114,8'd164} : s = 170;
	{8'd114,8'd165} : s = 313;
	{8'd114,8'd166} : s = 52;
	{8'd114,8'd167} : s = 169;
	{8'd114,8'd168} : s = 166;
	{8'd114,8'd169} : s = 310;
	{8'd114,8'd170} : s = 165;
	{8'd114,8'd171} : s = 309;
	{8'd114,8'd172} : s = 307;
	{8'd114,8'd173} : s = 427;
	{8'd114,8'd174} : s = 6;
	{8'd114,8'd175} : s = 50;
	{8'd114,8'd176} : s = 49;
	{8'd114,8'd177} : s = 163;
	{8'd114,8'd178} : s = 44;
	{8'd114,8'd179} : s = 156;
	{8'd114,8'd180} : s = 154;
	{8'd114,8'd181} : s = 302;
	{8'd114,8'd182} : s = 42;
	{8'd114,8'd183} : s = 153;
	{8'd114,8'd184} : s = 150;
	{8'd114,8'd185} : s = 301;
	{8'd114,8'd186} : s = 149;
	{8'd114,8'd187} : s = 299;
	{8'd114,8'd188} : s = 295;
	{8'd114,8'd189} : s = 423;
	{8'd114,8'd190} : s = 41;
	{8'd114,8'd191} : s = 147;
	{8'd114,8'd192} : s = 142;
	{8'd114,8'd193} : s = 286;
	{8'd114,8'd194} : s = 141;
	{8'd114,8'd195} : s = 285;
	{8'd114,8'd196} : s = 283;
	{8'd114,8'd197} : s = 414;
	{8'd114,8'd198} : s = 139;
	{8'd114,8'd199} : s = 279;
	{8'd114,8'd200} : s = 271;
	{8'd114,8'd201} : s = 413;
	{8'd114,8'd202} : s = 248;
	{8'd114,8'd203} : s = 411;
	{8'd114,8'd204} : s = 407;
	{8'd114,8'd205} : s = 491;
	{8'd114,8'd206} : s = 5;
	{8'd114,8'd207} : s = 38;
	{8'd114,8'd208} : s = 37;
	{8'd114,8'd209} : s = 135;
	{8'd114,8'd210} : s = 35;
	{8'd114,8'd211} : s = 120;
	{8'd114,8'd212} : s = 116;
	{8'd114,8'd213} : s = 244;
	{8'd114,8'd214} : s = 28;
	{8'd114,8'd215} : s = 114;
	{8'd114,8'd216} : s = 113;
	{8'd114,8'd217} : s = 242;
	{8'd114,8'd218} : s = 108;
	{8'd114,8'd219} : s = 241;
	{8'd114,8'd220} : s = 236;
	{8'd114,8'd221} : s = 399;
	{8'd114,8'd222} : s = 26;
	{8'd114,8'd223} : s = 106;
	{8'd114,8'd224} : s = 105;
	{8'd114,8'd225} : s = 234;
	{8'd114,8'd226} : s = 102;
	{8'd114,8'd227} : s = 233;
	{8'd114,8'd228} : s = 230;
	{8'd114,8'd229} : s = 380;
	{8'd114,8'd230} : s = 101;
	{8'd114,8'd231} : s = 229;
	{8'd114,8'd232} : s = 227;
	{8'd114,8'd233} : s = 378;
	{8'd114,8'd234} : s = 220;
	{8'd114,8'd235} : s = 377;
	{8'd114,8'd236} : s = 374;
	{8'd114,8'd237} : s = 487;
	{8'd114,8'd238} : s = 25;
	{8'd114,8'd239} : s = 99;
	{8'd114,8'd240} : s = 92;
	{8'd114,8'd241} : s = 218;
	{8'd114,8'd242} : s = 90;
	{8'd114,8'd243} : s = 217;
	{8'd114,8'd244} : s = 214;
	{8'd114,8'd245} : s = 373;
	{8'd114,8'd246} : s = 89;
	{8'd114,8'd247} : s = 213;
	{8'd114,8'd248} : s = 211;
	{8'd114,8'd249} : s = 371;
	{8'd114,8'd250} : s = 206;
	{8'd114,8'd251} : s = 366;
	{8'd114,8'd252} : s = 365;
	{8'd114,8'd253} : s = 478;
	{8'd114,8'd254} : s = 86;
	{8'd114,8'd255} : s = 205;
	{8'd115,8'd0} : s = 440;
	{8'd115,8'd1} : s = 326;
	{8'd115,8'd2} : s = 436;
	{8'd115,8'd3} : s = 434;
	{8'd115,8'd4} : s = 497;
	{8'd115,8'd5} : s = 325;
	{8'd115,8'd6} : s = 433;
	{8'd115,8'd7} : s = 428;
	{8'd115,8'd8} : s = 492;
	{8'd115,8'd9} : s = 426;
	{8'd115,8'd10} : s = 490;
	{8'd115,8'd11} : s = 489;
	{8'd115,8'd12} : s = 508;
	{8'd115,8'd13} : s = 2;
	{8'd115,8'd14} : s = 48;
	{8'd115,8'd15} : s = 40;
	{8'd115,8'd16} : s = 168;
	{8'd115,8'd17} : s = 36;
	{8'd115,8'd18} : s = 164;
	{8'd115,8'd19} : s = 162;
	{8'd115,8'd20} : s = 323;
	{8'd115,8'd21} : s = 34;
	{8'd115,8'd22} : s = 161;
	{8'd115,8'd23} : s = 152;
	{8'd115,8'd24} : s = 312;
	{8'd115,8'd25} : s = 148;
	{8'd115,8'd26} : s = 308;
	{8'd115,8'd27} : s = 306;
	{8'd115,8'd28} : s = 425;
	{8'd115,8'd29} : s = 33;
	{8'd115,8'd30} : s = 146;
	{8'd115,8'd31} : s = 145;
	{8'd115,8'd32} : s = 305;
	{8'd115,8'd33} : s = 140;
	{8'd115,8'd34} : s = 300;
	{8'd115,8'd35} : s = 298;
	{8'd115,8'd36} : s = 422;
	{8'd115,8'd37} : s = 138;
	{8'd115,8'd38} : s = 297;
	{8'd115,8'd39} : s = 294;
	{8'd115,8'd40} : s = 421;
	{8'd115,8'd41} : s = 293;
	{8'd115,8'd42} : s = 419;
	{8'd115,8'd43} : s = 412;
	{8'd115,8'd44} : s = 486;
	{8'd115,8'd45} : s = 24;
	{8'd115,8'd46} : s = 137;
	{8'd115,8'd47} : s = 134;
	{8'd115,8'd48} : s = 291;
	{8'd115,8'd49} : s = 133;
	{8'd115,8'd50} : s = 284;
	{8'd115,8'd51} : s = 282;
	{8'd115,8'd52} : s = 410;
	{8'd115,8'd53} : s = 131;
	{8'd115,8'd54} : s = 281;
	{8'd115,8'd55} : s = 278;
	{8'd115,8'd56} : s = 409;
	{8'd115,8'd57} : s = 277;
	{8'd115,8'd58} : s = 406;
	{8'd115,8'd59} : s = 405;
	{8'd115,8'd60} : s = 485;
	{8'd115,8'd61} : s = 112;
	{8'd115,8'd62} : s = 275;
	{8'd115,8'd63} : s = 270;
	{8'd115,8'd64} : s = 403;
	{8'd115,8'd65} : s = 269;
	{8'd115,8'd66} : s = 398;
	{8'd115,8'd67} : s = 397;
	{8'd115,8'd68} : s = 483;
	{8'd115,8'd69} : s = 267;
	{8'd115,8'd70} : s = 395;
	{8'd115,8'd71} : s = 391;
	{8'd115,8'd72} : s = 476;
	{8'd115,8'd73} : s = 376;
	{8'd115,8'd74} : s = 474;
	{8'd115,8'd75} : s = 473;
	{8'd115,8'd76} : s = 506;
	{8'd115,8'd77} : s = 20;
	{8'd115,8'd78} : s = 104;
	{8'd115,8'd79} : s = 100;
	{8'd115,8'd80} : s = 263;
	{8'd115,8'd81} : s = 98;
	{8'd115,8'd82} : s = 240;
	{8'd115,8'd83} : s = 232;
	{8'd115,8'd84} : s = 372;
	{8'd115,8'd85} : s = 97;
	{8'd115,8'd86} : s = 228;
	{8'd115,8'd87} : s = 226;
	{8'd115,8'd88} : s = 370;
	{8'd115,8'd89} : s = 225;
	{8'd115,8'd90} : s = 369;
	{8'd115,8'd91} : s = 364;
	{8'd115,8'd92} : s = 470;
	{8'd115,8'd93} : s = 88;
	{8'd115,8'd94} : s = 216;
	{8'd115,8'd95} : s = 212;
	{8'd115,8'd96} : s = 362;
	{8'd115,8'd97} : s = 210;
	{8'd115,8'd98} : s = 361;
	{8'd115,8'd99} : s = 358;
	{8'd115,8'd100} : s = 469;
	{8'd115,8'd101} : s = 209;
	{8'd115,8'd102} : s = 357;
	{8'd115,8'd103} : s = 355;
	{8'd115,8'd104} : s = 467;
	{8'd115,8'd105} : s = 348;
	{8'd115,8'd106} : s = 462;
	{8'd115,8'd107} : s = 461;
	{8'd115,8'd108} : s = 505;
	{8'd115,8'd109} : s = 84;
	{8'd115,8'd110} : s = 204;
	{8'd115,8'd111} : s = 202;
	{8'd115,8'd112} : s = 346;
	{8'd115,8'd113} : s = 201;
	{8'd115,8'd114} : s = 345;
	{8'd115,8'd115} : s = 342;
	{8'd115,8'd116} : s = 459;
	{8'd115,8'd117} : s = 198;
	{8'd115,8'd118} : s = 341;
	{8'd115,8'd119} : s = 339;
	{8'd115,8'd120} : s = 455;
	{8'd115,8'd121} : s = 334;
	{8'd115,8'd122} : s = 444;
	{8'd115,8'd123} : s = 442;
	{8'd115,8'd124} : s = 502;
	{8'd115,8'd125} : s = 197;
	{8'd115,8'd126} : s = 333;
	{8'd115,8'd127} : s = 331;
	{8'd115,8'd128} : s = 441;
	{8'd115,8'd129} : s = 327;
	{8'd115,8'd130} : s = 438;
	{8'd115,8'd131} : s = 437;
	{8'd115,8'd132} : s = 501;
	{8'd115,8'd133} : s = 316;
	{8'd115,8'd134} : s = 435;
	{8'd115,8'd135} : s = 430;
	{8'd115,8'd136} : s = 499;
	{8'd115,8'd137} : s = 429;
	{8'd115,8'd138} : s = 494;
	{8'd115,8'd139} : s = 493;
	{8'd115,8'd140} : s = 510;
	{8'd115,8'd141} : s = 1;
	{8'd115,8'd142} : s = 18;
	{8'd115,8'd143} : s = 17;
	{8'd115,8'd144} : s = 82;
	{8'd115,8'd145} : s = 12;
	{8'd115,8'd146} : s = 81;
	{8'd115,8'd147} : s = 76;
	{8'd115,8'd148} : s = 195;
	{8'd115,8'd149} : s = 10;
	{8'd115,8'd150} : s = 74;
	{8'd115,8'd151} : s = 73;
	{8'd115,8'd152} : s = 184;
	{8'd115,8'd153} : s = 70;
	{8'd115,8'd154} : s = 180;
	{8'd115,8'd155} : s = 178;
	{8'd115,8'd156} : s = 314;
	{8'd115,8'd157} : s = 9;
	{8'd115,8'd158} : s = 69;
	{8'd115,8'd159} : s = 67;
	{8'd115,8'd160} : s = 177;
	{8'd115,8'd161} : s = 56;
	{8'd115,8'd162} : s = 172;
	{8'd115,8'd163} : s = 170;
	{8'd115,8'd164} : s = 313;
	{8'd115,8'd165} : s = 52;
	{8'd115,8'd166} : s = 169;
	{8'd115,8'd167} : s = 166;
	{8'd115,8'd168} : s = 310;
	{8'd115,8'd169} : s = 165;
	{8'd115,8'd170} : s = 309;
	{8'd115,8'd171} : s = 307;
	{8'd115,8'd172} : s = 427;
	{8'd115,8'd173} : s = 6;
	{8'd115,8'd174} : s = 50;
	{8'd115,8'd175} : s = 49;
	{8'd115,8'd176} : s = 163;
	{8'd115,8'd177} : s = 44;
	{8'd115,8'd178} : s = 156;
	{8'd115,8'd179} : s = 154;
	{8'd115,8'd180} : s = 302;
	{8'd115,8'd181} : s = 42;
	{8'd115,8'd182} : s = 153;
	{8'd115,8'd183} : s = 150;
	{8'd115,8'd184} : s = 301;
	{8'd115,8'd185} : s = 149;
	{8'd115,8'd186} : s = 299;
	{8'd115,8'd187} : s = 295;
	{8'd115,8'd188} : s = 423;
	{8'd115,8'd189} : s = 41;
	{8'd115,8'd190} : s = 147;
	{8'd115,8'd191} : s = 142;
	{8'd115,8'd192} : s = 286;
	{8'd115,8'd193} : s = 141;
	{8'd115,8'd194} : s = 285;
	{8'd115,8'd195} : s = 283;
	{8'd115,8'd196} : s = 414;
	{8'd115,8'd197} : s = 139;
	{8'd115,8'd198} : s = 279;
	{8'd115,8'd199} : s = 271;
	{8'd115,8'd200} : s = 413;
	{8'd115,8'd201} : s = 248;
	{8'd115,8'd202} : s = 411;
	{8'd115,8'd203} : s = 407;
	{8'd115,8'd204} : s = 491;
	{8'd115,8'd205} : s = 5;
	{8'd115,8'd206} : s = 38;
	{8'd115,8'd207} : s = 37;
	{8'd115,8'd208} : s = 135;
	{8'd115,8'd209} : s = 35;
	{8'd115,8'd210} : s = 120;
	{8'd115,8'd211} : s = 116;
	{8'd115,8'd212} : s = 244;
	{8'd115,8'd213} : s = 28;
	{8'd115,8'd214} : s = 114;
	{8'd115,8'd215} : s = 113;
	{8'd115,8'd216} : s = 242;
	{8'd115,8'd217} : s = 108;
	{8'd115,8'd218} : s = 241;
	{8'd115,8'd219} : s = 236;
	{8'd115,8'd220} : s = 399;
	{8'd115,8'd221} : s = 26;
	{8'd115,8'd222} : s = 106;
	{8'd115,8'd223} : s = 105;
	{8'd115,8'd224} : s = 234;
	{8'd115,8'd225} : s = 102;
	{8'd115,8'd226} : s = 233;
	{8'd115,8'd227} : s = 230;
	{8'd115,8'd228} : s = 380;
	{8'd115,8'd229} : s = 101;
	{8'd115,8'd230} : s = 229;
	{8'd115,8'd231} : s = 227;
	{8'd115,8'd232} : s = 378;
	{8'd115,8'd233} : s = 220;
	{8'd115,8'd234} : s = 377;
	{8'd115,8'd235} : s = 374;
	{8'd115,8'd236} : s = 487;
	{8'd115,8'd237} : s = 25;
	{8'd115,8'd238} : s = 99;
	{8'd115,8'd239} : s = 92;
	{8'd115,8'd240} : s = 218;
	{8'd115,8'd241} : s = 90;
	{8'd115,8'd242} : s = 217;
	{8'd115,8'd243} : s = 214;
	{8'd115,8'd244} : s = 373;
	{8'd115,8'd245} : s = 89;
	{8'd115,8'd246} : s = 213;
	{8'd115,8'd247} : s = 211;
	{8'd115,8'd248} : s = 371;
	{8'd115,8'd249} : s = 206;
	{8'd115,8'd250} : s = 366;
	{8'd115,8'd251} : s = 365;
	{8'd115,8'd252} : s = 478;
	{8'd115,8'd253} : s = 86;
	{8'd115,8'd254} : s = 205;
	{8'd115,8'd255} : s = 203;
	{8'd116,8'd0} : s = 326;
	{8'd116,8'd1} : s = 436;
	{8'd116,8'd2} : s = 434;
	{8'd116,8'd3} : s = 497;
	{8'd116,8'd4} : s = 325;
	{8'd116,8'd5} : s = 433;
	{8'd116,8'd6} : s = 428;
	{8'd116,8'd7} : s = 492;
	{8'd116,8'd8} : s = 426;
	{8'd116,8'd9} : s = 490;
	{8'd116,8'd10} : s = 489;
	{8'd116,8'd11} : s = 508;
	{8'd116,8'd12} : s = 2;
	{8'd116,8'd13} : s = 48;
	{8'd116,8'd14} : s = 40;
	{8'd116,8'd15} : s = 168;
	{8'd116,8'd16} : s = 36;
	{8'd116,8'd17} : s = 164;
	{8'd116,8'd18} : s = 162;
	{8'd116,8'd19} : s = 323;
	{8'd116,8'd20} : s = 34;
	{8'd116,8'd21} : s = 161;
	{8'd116,8'd22} : s = 152;
	{8'd116,8'd23} : s = 312;
	{8'd116,8'd24} : s = 148;
	{8'd116,8'd25} : s = 308;
	{8'd116,8'd26} : s = 306;
	{8'd116,8'd27} : s = 425;
	{8'd116,8'd28} : s = 33;
	{8'd116,8'd29} : s = 146;
	{8'd116,8'd30} : s = 145;
	{8'd116,8'd31} : s = 305;
	{8'd116,8'd32} : s = 140;
	{8'd116,8'd33} : s = 300;
	{8'd116,8'd34} : s = 298;
	{8'd116,8'd35} : s = 422;
	{8'd116,8'd36} : s = 138;
	{8'd116,8'd37} : s = 297;
	{8'd116,8'd38} : s = 294;
	{8'd116,8'd39} : s = 421;
	{8'd116,8'd40} : s = 293;
	{8'd116,8'd41} : s = 419;
	{8'd116,8'd42} : s = 412;
	{8'd116,8'd43} : s = 486;
	{8'd116,8'd44} : s = 24;
	{8'd116,8'd45} : s = 137;
	{8'd116,8'd46} : s = 134;
	{8'd116,8'd47} : s = 291;
	{8'd116,8'd48} : s = 133;
	{8'd116,8'd49} : s = 284;
	{8'd116,8'd50} : s = 282;
	{8'd116,8'd51} : s = 410;
	{8'd116,8'd52} : s = 131;
	{8'd116,8'd53} : s = 281;
	{8'd116,8'd54} : s = 278;
	{8'd116,8'd55} : s = 409;
	{8'd116,8'd56} : s = 277;
	{8'd116,8'd57} : s = 406;
	{8'd116,8'd58} : s = 405;
	{8'd116,8'd59} : s = 485;
	{8'd116,8'd60} : s = 112;
	{8'd116,8'd61} : s = 275;
	{8'd116,8'd62} : s = 270;
	{8'd116,8'd63} : s = 403;
	{8'd116,8'd64} : s = 269;
	{8'd116,8'd65} : s = 398;
	{8'd116,8'd66} : s = 397;
	{8'd116,8'd67} : s = 483;
	{8'd116,8'd68} : s = 267;
	{8'd116,8'd69} : s = 395;
	{8'd116,8'd70} : s = 391;
	{8'd116,8'd71} : s = 476;
	{8'd116,8'd72} : s = 376;
	{8'd116,8'd73} : s = 474;
	{8'd116,8'd74} : s = 473;
	{8'd116,8'd75} : s = 506;
	{8'd116,8'd76} : s = 20;
	{8'd116,8'd77} : s = 104;
	{8'd116,8'd78} : s = 100;
	{8'd116,8'd79} : s = 263;
	{8'd116,8'd80} : s = 98;
	{8'd116,8'd81} : s = 240;
	{8'd116,8'd82} : s = 232;
	{8'd116,8'd83} : s = 372;
	{8'd116,8'd84} : s = 97;
	{8'd116,8'd85} : s = 228;
	{8'd116,8'd86} : s = 226;
	{8'd116,8'd87} : s = 370;
	{8'd116,8'd88} : s = 225;
	{8'd116,8'd89} : s = 369;
	{8'd116,8'd90} : s = 364;
	{8'd116,8'd91} : s = 470;
	{8'd116,8'd92} : s = 88;
	{8'd116,8'd93} : s = 216;
	{8'd116,8'd94} : s = 212;
	{8'd116,8'd95} : s = 362;
	{8'd116,8'd96} : s = 210;
	{8'd116,8'd97} : s = 361;
	{8'd116,8'd98} : s = 358;
	{8'd116,8'd99} : s = 469;
	{8'd116,8'd100} : s = 209;
	{8'd116,8'd101} : s = 357;
	{8'd116,8'd102} : s = 355;
	{8'd116,8'd103} : s = 467;
	{8'd116,8'd104} : s = 348;
	{8'd116,8'd105} : s = 462;
	{8'd116,8'd106} : s = 461;
	{8'd116,8'd107} : s = 505;
	{8'd116,8'd108} : s = 84;
	{8'd116,8'd109} : s = 204;
	{8'd116,8'd110} : s = 202;
	{8'd116,8'd111} : s = 346;
	{8'd116,8'd112} : s = 201;
	{8'd116,8'd113} : s = 345;
	{8'd116,8'd114} : s = 342;
	{8'd116,8'd115} : s = 459;
	{8'd116,8'd116} : s = 198;
	{8'd116,8'd117} : s = 341;
	{8'd116,8'd118} : s = 339;
	{8'd116,8'd119} : s = 455;
	{8'd116,8'd120} : s = 334;
	{8'd116,8'd121} : s = 444;
	{8'd116,8'd122} : s = 442;
	{8'd116,8'd123} : s = 502;
	{8'd116,8'd124} : s = 197;
	{8'd116,8'd125} : s = 333;
	{8'd116,8'd126} : s = 331;
	{8'd116,8'd127} : s = 441;
	{8'd116,8'd128} : s = 327;
	{8'd116,8'd129} : s = 438;
	{8'd116,8'd130} : s = 437;
	{8'd116,8'd131} : s = 501;
	{8'd116,8'd132} : s = 316;
	{8'd116,8'd133} : s = 435;
	{8'd116,8'd134} : s = 430;
	{8'd116,8'd135} : s = 499;
	{8'd116,8'd136} : s = 429;
	{8'd116,8'd137} : s = 494;
	{8'd116,8'd138} : s = 493;
	{8'd116,8'd139} : s = 510;
	{8'd116,8'd140} : s = 1;
	{8'd116,8'd141} : s = 18;
	{8'd116,8'd142} : s = 17;
	{8'd116,8'd143} : s = 82;
	{8'd116,8'd144} : s = 12;
	{8'd116,8'd145} : s = 81;
	{8'd116,8'd146} : s = 76;
	{8'd116,8'd147} : s = 195;
	{8'd116,8'd148} : s = 10;
	{8'd116,8'd149} : s = 74;
	{8'd116,8'd150} : s = 73;
	{8'd116,8'd151} : s = 184;
	{8'd116,8'd152} : s = 70;
	{8'd116,8'd153} : s = 180;
	{8'd116,8'd154} : s = 178;
	{8'd116,8'd155} : s = 314;
	{8'd116,8'd156} : s = 9;
	{8'd116,8'd157} : s = 69;
	{8'd116,8'd158} : s = 67;
	{8'd116,8'd159} : s = 177;
	{8'd116,8'd160} : s = 56;
	{8'd116,8'd161} : s = 172;
	{8'd116,8'd162} : s = 170;
	{8'd116,8'd163} : s = 313;
	{8'd116,8'd164} : s = 52;
	{8'd116,8'd165} : s = 169;
	{8'd116,8'd166} : s = 166;
	{8'd116,8'd167} : s = 310;
	{8'd116,8'd168} : s = 165;
	{8'd116,8'd169} : s = 309;
	{8'd116,8'd170} : s = 307;
	{8'd116,8'd171} : s = 427;
	{8'd116,8'd172} : s = 6;
	{8'd116,8'd173} : s = 50;
	{8'd116,8'd174} : s = 49;
	{8'd116,8'd175} : s = 163;
	{8'd116,8'd176} : s = 44;
	{8'd116,8'd177} : s = 156;
	{8'd116,8'd178} : s = 154;
	{8'd116,8'd179} : s = 302;
	{8'd116,8'd180} : s = 42;
	{8'd116,8'd181} : s = 153;
	{8'd116,8'd182} : s = 150;
	{8'd116,8'd183} : s = 301;
	{8'd116,8'd184} : s = 149;
	{8'd116,8'd185} : s = 299;
	{8'd116,8'd186} : s = 295;
	{8'd116,8'd187} : s = 423;
	{8'd116,8'd188} : s = 41;
	{8'd116,8'd189} : s = 147;
	{8'd116,8'd190} : s = 142;
	{8'd116,8'd191} : s = 286;
	{8'd116,8'd192} : s = 141;
	{8'd116,8'd193} : s = 285;
	{8'd116,8'd194} : s = 283;
	{8'd116,8'd195} : s = 414;
	{8'd116,8'd196} : s = 139;
	{8'd116,8'd197} : s = 279;
	{8'd116,8'd198} : s = 271;
	{8'd116,8'd199} : s = 413;
	{8'd116,8'd200} : s = 248;
	{8'd116,8'd201} : s = 411;
	{8'd116,8'd202} : s = 407;
	{8'd116,8'd203} : s = 491;
	{8'd116,8'd204} : s = 5;
	{8'd116,8'd205} : s = 38;
	{8'd116,8'd206} : s = 37;
	{8'd116,8'd207} : s = 135;
	{8'd116,8'd208} : s = 35;
	{8'd116,8'd209} : s = 120;
	{8'd116,8'd210} : s = 116;
	{8'd116,8'd211} : s = 244;
	{8'd116,8'd212} : s = 28;
	{8'd116,8'd213} : s = 114;
	{8'd116,8'd214} : s = 113;
	{8'd116,8'd215} : s = 242;
	{8'd116,8'd216} : s = 108;
	{8'd116,8'd217} : s = 241;
	{8'd116,8'd218} : s = 236;
	{8'd116,8'd219} : s = 399;
	{8'd116,8'd220} : s = 26;
	{8'd116,8'd221} : s = 106;
	{8'd116,8'd222} : s = 105;
	{8'd116,8'd223} : s = 234;
	{8'd116,8'd224} : s = 102;
	{8'd116,8'd225} : s = 233;
	{8'd116,8'd226} : s = 230;
	{8'd116,8'd227} : s = 380;
	{8'd116,8'd228} : s = 101;
	{8'd116,8'd229} : s = 229;
	{8'd116,8'd230} : s = 227;
	{8'd116,8'd231} : s = 378;
	{8'd116,8'd232} : s = 220;
	{8'd116,8'd233} : s = 377;
	{8'd116,8'd234} : s = 374;
	{8'd116,8'd235} : s = 487;
	{8'd116,8'd236} : s = 25;
	{8'd116,8'd237} : s = 99;
	{8'd116,8'd238} : s = 92;
	{8'd116,8'd239} : s = 218;
	{8'd116,8'd240} : s = 90;
	{8'd116,8'd241} : s = 217;
	{8'd116,8'd242} : s = 214;
	{8'd116,8'd243} : s = 373;
	{8'd116,8'd244} : s = 89;
	{8'd116,8'd245} : s = 213;
	{8'd116,8'd246} : s = 211;
	{8'd116,8'd247} : s = 371;
	{8'd116,8'd248} : s = 206;
	{8'd116,8'd249} : s = 366;
	{8'd116,8'd250} : s = 365;
	{8'd116,8'd251} : s = 478;
	{8'd116,8'd252} : s = 86;
	{8'd116,8'd253} : s = 205;
	{8'd116,8'd254} : s = 203;
	{8'd116,8'd255} : s = 363;
	{8'd117,8'd0} : s = 436;
	{8'd117,8'd1} : s = 434;
	{8'd117,8'd2} : s = 497;
	{8'd117,8'd3} : s = 325;
	{8'd117,8'd4} : s = 433;
	{8'd117,8'd5} : s = 428;
	{8'd117,8'd6} : s = 492;
	{8'd117,8'd7} : s = 426;
	{8'd117,8'd8} : s = 490;
	{8'd117,8'd9} : s = 489;
	{8'd117,8'd10} : s = 508;
	{8'd117,8'd11} : s = 2;
	{8'd117,8'd12} : s = 48;
	{8'd117,8'd13} : s = 40;
	{8'd117,8'd14} : s = 168;
	{8'd117,8'd15} : s = 36;
	{8'd117,8'd16} : s = 164;
	{8'd117,8'd17} : s = 162;
	{8'd117,8'd18} : s = 323;
	{8'd117,8'd19} : s = 34;
	{8'd117,8'd20} : s = 161;
	{8'd117,8'd21} : s = 152;
	{8'd117,8'd22} : s = 312;
	{8'd117,8'd23} : s = 148;
	{8'd117,8'd24} : s = 308;
	{8'd117,8'd25} : s = 306;
	{8'd117,8'd26} : s = 425;
	{8'd117,8'd27} : s = 33;
	{8'd117,8'd28} : s = 146;
	{8'd117,8'd29} : s = 145;
	{8'd117,8'd30} : s = 305;
	{8'd117,8'd31} : s = 140;
	{8'd117,8'd32} : s = 300;
	{8'd117,8'd33} : s = 298;
	{8'd117,8'd34} : s = 422;
	{8'd117,8'd35} : s = 138;
	{8'd117,8'd36} : s = 297;
	{8'd117,8'd37} : s = 294;
	{8'd117,8'd38} : s = 421;
	{8'd117,8'd39} : s = 293;
	{8'd117,8'd40} : s = 419;
	{8'd117,8'd41} : s = 412;
	{8'd117,8'd42} : s = 486;
	{8'd117,8'd43} : s = 24;
	{8'd117,8'd44} : s = 137;
	{8'd117,8'd45} : s = 134;
	{8'd117,8'd46} : s = 291;
	{8'd117,8'd47} : s = 133;
	{8'd117,8'd48} : s = 284;
	{8'd117,8'd49} : s = 282;
	{8'd117,8'd50} : s = 410;
	{8'd117,8'd51} : s = 131;
	{8'd117,8'd52} : s = 281;
	{8'd117,8'd53} : s = 278;
	{8'd117,8'd54} : s = 409;
	{8'd117,8'd55} : s = 277;
	{8'd117,8'd56} : s = 406;
	{8'd117,8'd57} : s = 405;
	{8'd117,8'd58} : s = 485;
	{8'd117,8'd59} : s = 112;
	{8'd117,8'd60} : s = 275;
	{8'd117,8'd61} : s = 270;
	{8'd117,8'd62} : s = 403;
	{8'd117,8'd63} : s = 269;
	{8'd117,8'd64} : s = 398;
	{8'd117,8'd65} : s = 397;
	{8'd117,8'd66} : s = 483;
	{8'd117,8'd67} : s = 267;
	{8'd117,8'd68} : s = 395;
	{8'd117,8'd69} : s = 391;
	{8'd117,8'd70} : s = 476;
	{8'd117,8'd71} : s = 376;
	{8'd117,8'd72} : s = 474;
	{8'd117,8'd73} : s = 473;
	{8'd117,8'd74} : s = 506;
	{8'd117,8'd75} : s = 20;
	{8'd117,8'd76} : s = 104;
	{8'd117,8'd77} : s = 100;
	{8'd117,8'd78} : s = 263;
	{8'd117,8'd79} : s = 98;
	{8'd117,8'd80} : s = 240;
	{8'd117,8'd81} : s = 232;
	{8'd117,8'd82} : s = 372;
	{8'd117,8'd83} : s = 97;
	{8'd117,8'd84} : s = 228;
	{8'd117,8'd85} : s = 226;
	{8'd117,8'd86} : s = 370;
	{8'd117,8'd87} : s = 225;
	{8'd117,8'd88} : s = 369;
	{8'd117,8'd89} : s = 364;
	{8'd117,8'd90} : s = 470;
	{8'd117,8'd91} : s = 88;
	{8'd117,8'd92} : s = 216;
	{8'd117,8'd93} : s = 212;
	{8'd117,8'd94} : s = 362;
	{8'd117,8'd95} : s = 210;
	{8'd117,8'd96} : s = 361;
	{8'd117,8'd97} : s = 358;
	{8'd117,8'd98} : s = 469;
	{8'd117,8'd99} : s = 209;
	{8'd117,8'd100} : s = 357;
	{8'd117,8'd101} : s = 355;
	{8'd117,8'd102} : s = 467;
	{8'd117,8'd103} : s = 348;
	{8'd117,8'd104} : s = 462;
	{8'd117,8'd105} : s = 461;
	{8'd117,8'd106} : s = 505;
	{8'd117,8'd107} : s = 84;
	{8'd117,8'd108} : s = 204;
	{8'd117,8'd109} : s = 202;
	{8'd117,8'd110} : s = 346;
	{8'd117,8'd111} : s = 201;
	{8'd117,8'd112} : s = 345;
	{8'd117,8'd113} : s = 342;
	{8'd117,8'd114} : s = 459;
	{8'd117,8'd115} : s = 198;
	{8'd117,8'd116} : s = 341;
	{8'd117,8'd117} : s = 339;
	{8'd117,8'd118} : s = 455;
	{8'd117,8'd119} : s = 334;
	{8'd117,8'd120} : s = 444;
	{8'd117,8'd121} : s = 442;
	{8'd117,8'd122} : s = 502;
	{8'd117,8'd123} : s = 197;
	{8'd117,8'd124} : s = 333;
	{8'd117,8'd125} : s = 331;
	{8'd117,8'd126} : s = 441;
	{8'd117,8'd127} : s = 327;
	{8'd117,8'd128} : s = 438;
	{8'd117,8'd129} : s = 437;
	{8'd117,8'd130} : s = 501;
	{8'd117,8'd131} : s = 316;
	{8'd117,8'd132} : s = 435;
	{8'd117,8'd133} : s = 430;
	{8'd117,8'd134} : s = 499;
	{8'd117,8'd135} : s = 429;
	{8'd117,8'd136} : s = 494;
	{8'd117,8'd137} : s = 493;
	{8'd117,8'd138} : s = 510;
	{8'd117,8'd139} : s = 1;
	{8'd117,8'd140} : s = 18;
	{8'd117,8'd141} : s = 17;
	{8'd117,8'd142} : s = 82;
	{8'd117,8'd143} : s = 12;
	{8'd117,8'd144} : s = 81;
	{8'd117,8'd145} : s = 76;
	{8'd117,8'd146} : s = 195;
	{8'd117,8'd147} : s = 10;
	{8'd117,8'd148} : s = 74;
	{8'd117,8'd149} : s = 73;
	{8'd117,8'd150} : s = 184;
	{8'd117,8'd151} : s = 70;
	{8'd117,8'd152} : s = 180;
	{8'd117,8'd153} : s = 178;
	{8'd117,8'd154} : s = 314;
	{8'd117,8'd155} : s = 9;
	{8'd117,8'd156} : s = 69;
	{8'd117,8'd157} : s = 67;
	{8'd117,8'd158} : s = 177;
	{8'd117,8'd159} : s = 56;
	{8'd117,8'd160} : s = 172;
	{8'd117,8'd161} : s = 170;
	{8'd117,8'd162} : s = 313;
	{8'd117,8'd163} : s = 52;
	{8'd117,8'd164} : s = 169;
	{8'd117,8'd165} : s = 166;
	{8'd117,8'd166} : s = 310;
	{8'd117,8'd167} : s = 165;
	{8'd117,8'd168} : s = 309;
	{8'd117,8'd169} : s = 307;
	{8'd117,8'd170} : s = 427;
	{8'd117,8'd171} : s = 6;
	{8'd117,8'd172} : s = 50;
	{8'd117,8'd173} : s = 49;
	{8'd117,8'd174} : s = 163;
	{8'd117,8'd175} : s = 44;
	{8'd117,8'd176} : s = 156;
	{8'd117,8'd177} : s = 154;
	{8'd117,8'd178} : s = 302;
	{8'd117,8'd179} : s = 42;
	{8'd117,8'd180} : s = 153;
	{8'd117,8'd181} : s = 150;
	{8'd117,8'd182} : s = 301;
	{8'd117,8'd183} : s = 149;
	{8'd117,8'd184} : s = 299;
	{8'd117,8'd185} : s = 295;
	{8'd117,8'd186} : s = 423;
	{8'd117,8'd187} : s = 41;
	{8'd117,8'd188} : s = 147;
	{8'd117,8'd189} : s = 142;
	{8'd117,8'd190} : s = 286;
	{8'd117,8'd191} : s = 141;
	{8'd117,8'd192} : s = 285;
	{8'd117,8'd193} : s = 283;
	{8'd117,8'd194} : s = 414;
	{8'd117,8'd195} : s = 139;
	{8'd117,8'd196} : s = 279;
	{8'd117,8'd197} : s = 271;
	{8'd117,8'd198} : s = 413;
	{8'd117,8'd199} : s = 248;
	{8'd117,8'd200} : s = 411;
	{8'd117,8'd201} : s = 407;
	{8'd117,8'd202} : s = 491;
	{8'd117,8'd203} : s = 5;
	{8'd117,8'd204} : s = 38;
	{8'd117,8'd205} : s = 37;
	{8'd117,8'd206} : s = 135;
	{8'd117,8'd207} : s = 35;
	{8'd117,8'd208} : s = 120;
	{8'd117,8'd209} : s = 116;
	{8'd117,8'd210} : s = 244;
	{8'd117,8'd211} : s = 28;
	{8'd117,8'd212} : s = 114;
	{8'd117,8'd213} : s = 113;
	{8'd117,8'd214} : s = 242;
	{8'd117,8'd215} : s = 108;
	{8'd117,8'd216} : s = 241;
	{8'd117,8'd217} : s = 236;
	{8'd117,8'd218} : s = 399;
	{8'd117,8'd219} : s = 26;
	{8'd117,8'd220} : s = 106;
	{8'd117,8'd221} : s = 105;
	{8'd117,8'd222} : s = 234;
	{8'd117,8'd223} : s = 102;
	{8'd117,8'd224} : s = 233;
	{8'd117,8'd225} : s = 230;
	{8'd117,8'd226} : s = 380;
	{8'd117,8'd227} : s = 101;
	{8'd117,8'd228} : s = 229;
	{8'd117,8'd229} : s = 227;
	{8'd117,8'd230} : s = 378;
	{8'd117,8'd231} : s = 220;
	{8'd117,8'd232} : s = 377;
	{8'd117,8'd233} : s = 374;
	{8'd117,8'd234} : s = 487;
	{8'd117,8'd235} : s = 25;
	{8'd117,8'd236} : s = 99;
	{8'd117,8'd237} : s = 92;
	{8'd117,8'd238} : s = 218;
	{8'd117,8'd239} : s = 90;
	{8'd117,8'd240} : s = 217;
	{8'd117,8'd241} : s = 214;
	{8'd117,8'd242} : s = 373;
	{8'd117,8'd243} : s = 89;
	{8'd117,8'd244} : s = 213;
	{8'd117,8'd245} : s = 211;
	{8'd117,8'd246} : s = 371;
	{8'd117,8'd247} : s = 206;
	{8'd117,8'd248} : s = 366;
	{8'd117,8'd249} : s = 365;
	{8'd117,8'd250} : s = 478;
	{8'd117,8'd251} : s = 86;
	{8'd117,8'd252} : s = 205;
	{8'd117,8'd253} : s = 203;
	{8'd117,8'd254} : s = 363;
	{8'd117,8'd255} : s = 199;
	{8'd118,8'd0} : s = 434;
	{8'd118,8'd1} : s = 497;
	{8'd118,8'd2} : s = 325;
	{8'd118,8'd3} : s = 433;
	{8'd118,8'd4} : s = 428;
	{8'd118,8'd5} : s = 492;
	{8'd118,8'd6} : s = 426;
	{8'd118,8'd7} : s = 490;
	{8'd118,8'd8} : s = 489;
	{8'd118,8'd9} : s = 508;
	{8'd118,8'd10} : s = 2;
	{8'd118,8'd11} : s = 48;
	{8'd118,8'd12} : s = 40;
	{8'd118,8'd13} : s = 168;
	{8'd118,8'd14} : s = 36;
	{8'd118,8'd15} : s = 164;
	{8'd118,8'd16} : s = 162;
	{8'd118,8'd17} : s = 323;
	{8'd118,8'd18} : s = 34;
	{8'd118,8'd19} : s = 161;
	{8'd118,8'd20} : s = 152;
	{8'd118,8'd21} : s = 312;
	{8'd118,8'd22} : s = 148;
	{8'd118,8'd23} : s = 308;
	{8'd118,8'd24} : s = 306;
	{8'd118,8'd25} : s = 425;
	{8'd118,8'd26} : s = 33;
	{8'd118,8'd27} : s = 146;
	{8'd118,8'd28} : s = 145;
	{8'd118,8'd29} : s = 305;
	{8'd118,8'd30} : s = 140;
	{8'd118,8'd31} : s = 300;
	{8'd118,8'd32} : s = 298;
	{8'd118,8'd33} : s = 422;
	{8'd118,8'd34} : s = 138;
	{8'd118,8'd35} : s = 297;
	{8'd118,8'd36} : s = 294;
	{8'd118,8'd37} : s = 421;
	{8'd118,8'd38} : s = 293;
	{8'd118,8'd39} : s = 419;
	{8'd118,8'd40} : s = 412;
	{8'd118,8'd41} : s = 486;
	{8'd118,8'd42} : s = 24;
	{8'd118,8'd43} : s = 137;
	{8'd118,8'd44} : s = 134;
	{8'd118,8'd45} : s = 291;
	{8'd118,8'd46} : s = 133;
	{8'd118,8'd47} : s = 284;
	{8'd118,8'd48} : s = 282;
	{8'd118,8'd49} : s = 410;
	{8'd118,8'd50} : s = 131;
	{8'd118,8'd51} : s = 281;
	{8'd118,8'd52} : s = 278;
	{8'd118,8'd53} : s = 409;
	{8'd118,8'd54} : s = 277;
	{8'd118,8'd55} : s = 406;
	{8'd118,8'd56} : s = 405;
	{8'd118,8'd57} : s = 485;
	{8'd118,8'd58} : s = 112;
	{8'd118,8'd59} : s = 275;
	{8'd118,8'd60} : s = 270;
	{8'd118,8'd61} : s = 403;
	{8'd118,8'd62} : s = 269;
	{8'd118,8'd63} : s = 398;
	{8'd118,8'd64} : s = 397;
	{8'd118,8'd65} : s = 483;
	{8'd118,8'd66} : s = 267;
	{8'd118,8'd67} : s = 395;
	{8'd118,8'd68} : s = 391;
	{8'd118,8'd69} : s = 476;
	{8'd118,8'd70} : s = 376;
	{8'd118,8'd71} : s = 474;
	{8'd118,8'd72} : s = 473;
	{8'd118,8'd73} : s = 506;
	{8'd118,8'd74} : s = 20;
	{8'd118,8'd75} : s = 104;
	{8'd118,8'd76} : s = 100;
	{8'd118,8'd77} : s = 263;
	{8'd118,8'd78} : s = 98;
	{8'd118,8'd79} : s = 240;
	{8'd118,8'd80} : s = 232;
	{8'd118,8'd81} : s = 372;
	{8'd118,8'd82} : s = 97;
	{8'd118,8'd83} : s = 228;
	{8'd118,8'd84} : s = 226;
	{8'd118,8'd85} : s = 370;
	{8'd118,8'd86} : s = 225;
	{8'd118,8'd87} : s = 369;
	{8'd118,8'd88} : s = 364;
	{8'd118,8'd89} : s = 470;
	{8'd118,8'd90} : s = 88;
	{8'd118,8'd91} : s = 216;
	{8'd118,8'd92} : s = 212;
	{8'd118,8'd93} : s = 362;
	{8'd118,8'd94} : s = 210;
	{8'd118,8'd95} : s = 361;
	{8'd118,8'd96} : s = 358;
	{8'd118,8'd97} : s = 469;
	{8'd118,8'd98} : s = 209;
	{8'd118,8'd99} : s = 357;
	{8'd118,8'd100} : s = 355;
	{8'd118,8'd101} : s = 467;
	{8'd118,8'd102} : s = 348;
	{8'd118,8'd103} : s = 462;
	{8'd118,8'd104} : s = 461;
	{8'd118,8'd105} : s = 505;
	{8'd118,8'd106} : s = 84;
	{8'd118,8'd107} : s = 204;
	{8'd118,8'd108} : s = 202;
	{8'd118,8'd109} : s = 346;
	{8'd118,8'd110} : s = 201;
	{8'd118,8'd111} : s = 345;
	{8'd118,8'd112} : s = 342;
	{8'd118,8'd113} : s = 459;
	{8'd118,8'd114} : s = 198;
	{8'd118,8'd115} : s = 341;
	{8'd118,8'd116} : s = 339;
	{8'd118,8'd117} : s = 455;
	{8'd118,8'd118} : s = 334;
	{8'd118,8'd119} : s = 444;
	{8'd118,8'd120} : s = 442;
	{8'd118,8'd121} : s = 502;
	{8'd118,8'd122} : s = 197;
	{8'd118,8'd123} : s = 333;
	{8'd118,8'd124} : s = 331;
	{8'd118,8'd125} : s = 441;
	{8'd118,8'd126} : s = 327;
	{8'd118,8'd127} : s = 438;
	{8'd118,8'd128} : s = 437;
	{8'd118,8'd129} : s = 501;
	{8'd118,8'd130} : s = 316;
	{8'd118,8'd131} : s = 435;
	{8'd118,8'd132} : s = 430;
	{8'd118,8'd133} : s = 499;
	{8'd118,8'd134} : s = 429;
	{8'd118,8'd135} : s = 494;
	{8'd118,8'd136} : s = 493;
	{8'd118,8'd137} : s = 510;
	{8'd118,8'd138} : s = 1;
	{8'd118,8'd139} : s = 18;
	{8'd118,8'd140} : s = 17;
	{8'd118,8'd141} : s = 82;
	{8'd118,8'd142} : s = 12;
	{8'd118,8'd143} : s = 81;
	{8'd118,8'd144} : s = 76;
	{8'd118,8'd145} : s = 195;
	{8'd118,8'd146} : s = 10;
	{8'd118,8'd147} : s = 74;
	{8'd118,8'd148} : s = 73;
	{8'd118,8'd149} : s = 184;
	{8'd118,8'd150} : s = 70;
	{8'd118,8'd151} : s = 180;
	{8'd118,8'd152} : s = 178;
	{8'd118,8'd153} : s = 314;
	{8'd118,8'd154} : s = 9;
	{8'd118,8'd155} : s = 69;
	{8'd118,8'd156} : s = 67;
	{8'd118,8'd157} : s = 177;
	{8'd118,8'd158} : s = 56;
	{8'd118,8'd159} : s = 172;
	{8'd118,8'd160} : s = 170;
	{8'd118,8'd161} : s = 313;
	{8'd118,8'd162} : s = 52;
	{8'd118,8'd163} : s = 169;
	{8'd118,8'd164} : s = 166;
	{8'd118,8'd165} : s = 310;
	{8'd118,8'd166} : s = 165;
	{8'd118,8'd167} : s = 309;
	{8'd118,8'd168} : s = 307;
	{8'd118,8'd169} : s = 427;
	{8'd118,8'd170} : s = 6;
	{8'd118,8'd171} : s = 50;
	{8'd118,8'd172} : s = 49;
	{8'd118,8'd173} : s = 163;
	{8'd118,8'd174} : s = 44;
	{8'd118,8'd175} : s = 156;
	{8'd118,8'd176} : s = 154;
	{8'd118,8'd177} : s = 302;
	{8'd118,8'd178} : s = 42;
	{8'd118,8'd179} : s = 153;
	{8'd118,8'd180} : s = 150;
	{8'd118,8'd181} : s = 301;
	{8'd118,8'd182} : s = 149;
	{8'd118,8'd183} : s = 299;
	{8'd118,8'd184} : s = 295;
	{8'd118,8'd185} : s = 423;
	{8'd118,8'd186} : s = 41;
	{8'd118,8'd187} : s = 147;
	{8'd118,8'd188} : s = 142;
	{8'd118,8'd189} : s = 286;
	{8'd118,8'd190} : s = 141;
	{8'd118,8'd191} : s = 285;
	{8'd118,8'd192} : s = 283;
	{8'd118,8'd193} : s = 414;
	{8'd118,8'd194} : s = 139;
	{8'd118,8'd195} : s = 279;
	{8'd118,8'd196} : s = 271;
	{8'd118,8'd197} : s = 413;
	{8'd118,8'd198} : s = 248;
	{8'd118,8'd199} : s = 411;
	{8'd118,8'd200} : s = 407;
	{8'd118,8'd201} : s = 491;
	{8'd118,8'd202} : s = 5;
	{8'd118,8'd203} : s = 38;
	{8'd118,8'd204} : s = 37;
	{8'd118,8'd205} : s = 135;
	{8'd118,8'd206} : s = 35;
	{8'd118,8'd207} : s = 120;
	{8'd118,8'd208} : s = 116;
	{8'd118,8'd209} : s = 244;
	{8'd118,8'd210} : s = 28;
	{8'd118,8'd211} : s = 114;
	{8'd118,8'd212} : s = 113;
	{8'd118,8'd213} : s = 242;
	{8'd118,8'd214} : s = 108;
	{8'd118,8'd215} : s = 241;
	{8'd118,8'd216} : s = 236;
	{8'd118,8'd217} : s = 399;
	{8'd118,8'd218} : s = 26;
	{8'd118,8'd219} : s = 106;
	{8'd118,8'd220} : s = 105;
	{8'd118,8'd221} : s = 234;
	{8'd118,8'd222} : s = 102;
	{8'd118,8'd223} : s = 233;
	{8'd118,8'd224} : s = 230;
	{8'd118,8'd225} : s = 380;
	{8'd118,8'd226} : s = 101;
	{8'd118,8'd227} : s = 229;
	{8'd118,8'd228} : s = 227;
	{8'd118,8'd229} : s = 378;
	{8'd118,8'd230} : s = 220;
	{8'd118,8'd231} : s = 377;
	{8'd118,8'd232} : s = 374;
	{8'd118,8'd233} : s = 487;
	{8'd118,8'd234} : s = 25;
	{8'd118,8'd235} : s = 99;
	{8'd118,8'd236} : s = 92;
	{8'd118,8'd237} : s = 218;
	{8'd118,8'd238} : s = 90;
	{8'd118,8'd239} : s = 217;
	{8'd118,8'd240} : s = 214;
	{8'd118,8'd241} : s = 373;
	{8'd118,8'd242} : s = 89;
	{8'd118,8'd243} : s = 213;
	{8'd118,8'd244} : s = 211;
	{8'd118,8'd245} : s = 371;
	{8'd118,8'd246} : s = 206;
	{8'd118,8'd247} : s = 366;
	{8'd118,8'd248} : s = 365;
	{8'd118,8'd249} : s = 478;
	{8'd118,8'd250} : s = 86;
	{8'd118,8'd251} : s = 205;
	{8'd118,8'd252} : s = 203;
	{8'd118,8'd253} : s = 363;
	{8'd118,8'd254} : s = 199;
	{8'd118,8'd255} : s = 359;
	{8'd119,8'd0} : s = 497;
	{8'd119,8'd1} : s = 325;
	{8'd119,8'd2} : s = 433;
	{8'd119,8'd3} : s = 428;
	{8'd119,8'd4} : s = 492;
	{8'd119,8'd5} : s = 426;
	{8'd119,8'd6} : s = 490;
	{8'd119,8'd7} : s = 489;
	{8'd119,8'd8} : s = 508;
	{8'd119,8'd9} : s = 2;
	{8'd119,8'd10} : s = 48;
	{8'd119,8'd11} : s = 40;
	{8'd119,8'd12} : s = 168;
	{8'd119,8'd13} : s = 36;
	{8'd119,8'd14} : s = 164;
	{8'd119,8'd15} : s = 162;
	{8'd119,8'd16} : s = 323;
	{8'd119,8'd17} : s = 34;
	{8'd119,8'd18} : s = 161;
	{8'd119,8'd19} : s = 152;
	{8'd119,8'd20} : s = 312;
	{8'd119,8'd21} : s = 148;
	{8'd119,8'd22} : s = 308;
	{8'd119,8'd23} : s = 306;
	{8'd119,8'd24} : s = 425;
	{8'd119,8'd25} : s = 33;
	{8'd119,8'd26} : s = 146;
	{8'd119,8'd27} : s = 145;
	{8'd119,8'd28} : s = 305;
	{8'd119,8'd29} : s = 140;
	{8'd119,8'd30} : s = 300;
	{8'd119,8'd31} : s = 298;
	{8'd119,8'd32} : s = 422;
	{8'd119,8'd33} : s = 138;
	{8'd119,8'd34} : s = 297;
	{8'd119,8'd35} : s = 294;
	{8'd119,8'd36} : s = 421;
	{8'd119,8'd37} : s = 293;
	{8'd119,8'd38} : s = 419;
	{8'd119,8'd39} : s = 412;
	{8'd119,8'd40} : s = 486;
	{8'd119,8'd41} : s = 24;
	{8'd119,8'd42} : s = 137;
	{8'd119,8'd43} : s = 134;
	{8'd119,8'd44} : s = 291;
	{8'd119,8'd45} : s = 133;
	{8'd119,8'd46} : s = 284;
	{8'd119,8'd47} : s = 282;
	{8'd119,8'd48} : s = 410;
	{8'd119,8'd49} : s = 131;
	{8'd119,8'd50} : s = 281;
	{8'd119,8'd51} : s = 278;
	{8'd119,8'd52} : s = 409;
	{8'd119,8'd53} : s = 277;
	{8'd119,8'd54} : s = 406;
	{8'd119,8'd55} : s = 405;
	{8'd119,8'd56} : s = 485;
	{8'd119,8'd57} : s = 112;
	{8'd119,8'd58} : s = 275;
	{8'd119,8'd59} : s = 270;
	{8'd119,8'd60} : s = 403;
	{8'd119,8'd61} : s = 269;
	{8'd119,8'd62} : s = 398;
	{8'd119,8'd63} : s = 397;
	{8'd119,8'd64} : s = 483;
	{8'd119,8'd65} : s = 267;
	{8'd119,8'd66} : s = 395;
	{8'd119,8'd67} : s = 391;
	{8'd119,8'd68} : s = 476;
	{8'd119,8'd69} : s = 376;
	{8'd119,8'd70} : s = 474;
	{8'd119,8'd71} : s = 473;
	{8'd119,8'd72} : s = 506;
	{8'd119,8'd73} : s = 20;
	{8'd119,8'd74} : s = 104;
	{8'd119,8'd75} : s = 100;
	{8'd119,8'd76} : s = 263;
	{8'd119,8'd77} : s = 98;
	{8'd119,8'd78} : s = 240;
	{8'd119,8'd79} : s = 232;
	{8'd119,8'd80} : s = 372;
	{8'd119,8'd81} : s = 97;
	{8'd119,8'd82} : s = 228;
	{8'd119,8'd83} : s = 226;
	{8'd119,8'd84} : s = 370;
	{8'd119,8'd85} : s = 225;
	{8'd119,8'd86} : s = 369;
	{8'd119,8'd87} : s = 364;
	{8'd119,8'd88} : s = 470;
	{8'd119,8'd89} : s = 88;
	{8'd119,8'd90} : s = 216;
	{8'd119,8'd91} : s = 212;
	{8'd119,8'd92} : s = 362;
	{8'd119,8'd93} : s = 210;
	{8'd119,8'd94} : s = 361;
	{8'd119,8'd95} : s = 358;
	{8'd119,8'd96} : s = 469;
	{8'd119,8'd97} : s = 209;
	{8'd119,8'd98} : s = 357;
	{8'd119,8'd99} : s = 355;
	{8'd119,8'd100} : s = 467;
	{8'd119,8'd101} : s = 348;
	{8'd119,8'd102} : s = 462;
	{8'd119,8'd103} : s = 461;
	{8'd119,8'd104} : s = 505;
	{8'd119,8'd105} : s = 84;
	{8'd119,8'd106} : s = 204;
	{8'd119,8'd107} : s = 202;
	{8'd119,8'd108} : s = 346;
	{8'd119,8'd109} : s = 201;
	{8'd119,8'd110} : s = 345;
	{8'd119,8'd111} : s = 342;
	{8'd119,8'd112} : s = 459;
	{8'd119,8'd113} : s = 198;
	{8'd119,8'd114} : s = 341;
	{8'd119,8'd115} : s = 339;
	{8'd119,8'd116} : s = 455;
	{8'd119,8'd117} : s = 334;
	{8'd119,8'd118} : s = 444;
	{8'd119,8'd119} : s = 442;
	{8'd119,8'd120} : s = 502;
	{8'd119,8'd121} : s = 197;
	{8'd119,8'd122} : s = 333;
	{8'd119,8'd123} : s = 331;
	{8'd119,8'd124} : s = 441;
	{8'd119,8'd125} : s = 327;
	{8'd119,8'd126} : s = 438;
	{8'd119,8'd127} : s = 437;
	{8'd119,8'd128} : s = 501;
	{8'd119,8'd129} : s = 316;
	{8'd119,8'd130} : s = 435;
	{8'd119,8'd131} : s = 430;
	{8'd119,8'd132} : s = 499;
	{8'd119,8'd133} : s = 429;
	{8'd119,8'd134} : s = 494;
	{8'd119,8'd135} : s = 493;
	{8'd119,8'd136} : s = 510;
	{8'd119,8'd137} : s = 1;
	{8'd119,8'd138} : s = 18;
	{8'd119,8'd139} : s = 17;
	{8'd119,8'd140} : s = 82;
	{8'd119,8'd141} : s = 12;
	{8'd119,8'd142} : s = 81;
	{8'd119,8'd143} : s = 76;
	{8'd119,8'd144} : s = 195;
	{8'd119,8'd145} : s = 10;
	{8'd119,8'd146} : s = 74;
	{8'd119,8'd147} : s = 73;
	{8'd119,8'd148} : s = 184;
	{8'd119,8'd149} : s = 70;
	{8'd119,8'd150} : s = 180;
	{8'd119,8'd151} : s = 178;
	{8'd119,8'd152} : s = 314;
	{8'd119,8'd153} : s = 9;
	{8'd119,8'd154} : s = 69;
	{8'd119,8'd155} : s = 67;
	{8'd119,8'd156} : s = 177;
	{8'd119,8'd157} : s = 56;
	{8'd119,8'd158} : s = 172;
	{8'd119,8'd159} : s = 170;
	{8'd119,8'd160} : s = 313;
	{8'd119,8'd161} : s = 52;
	{8'd119,8'd162} : s = 169;
	{8'd119,8'd163} : s = 166;
	{8'd119,8'd164} : s = 310;
	{8'd119,8'd165} : s = 165;
	{8'd119,8'd166} : s = 309;
	{8'd119,8'd167} : s = 307;
	{8'd119,8'd168} : s = 427;
	{8'd119,8'd169} : s = 6;
	{8'd119,8'd170} : s = 50;
	{8'd119,8'd171} : s = 49;
	{8'd119,8'd172} : s = 163;
	{8'd119,8'd173} : s = 44;
	{8'd119,8'd174} : s = 156;
	{8'd119,8'd175} : s = 154;
	{8'd119,8'd176} : s = 302;
	{8'd119,8'd177} : s = 42;
	{8'd119,8'd178} : s = 153;
	{8'd119,8'd179} : s = 150;
	{8'd119,8'd180} : s = 301;
	{8'd119,8'd181} : s = 149;
	{8'd119,8'd182} : s = 299;
	{8'd119,8'd183} : s = 295;
	{8'd119,8'd184} : s = 423;
	{8'd119,8'd185} : s = 41;
	{8'd119,8'd186} : s = 147;
	{8'd119,8'd187} : s = 142;
	{8'd119,8'd188} : s = 286;
	{8'd119,8'd189} : s = 141;
	{8'd119,8'd190} : s = 285;
	{8'd119,8'd191} : s = 283;
	{8'd119,8'd192} : s = 414;
	{8'd119,8'd193} : s = 139;
	{8'd119,8'd194} : s = 279;
	{8'd119,8'd195} : s = 271;
	{8'd119,8'd196} : s = 413;
	{8'd119,8'd197} : s = 248;
	{8'd119,8'd198} : s = 411;
	{8'd119,8'd199} : s = 407;
	{8'd119,8'd200} : s = 491;
	{8'd119,8'd201} : s = 5;
	{8'd119,8'd202} : s = 38;
	{8'd119,8'd203} : s = 37;
	{8'd119,8'd204} : s = 135;
	{8'd119,8'd205} : s = 35;
	{8'd119,8'd206} : s = 120;
	{8'd119,8'd207} : s = 116;
	{8'd119,8'd208} : s = 244;
	{8'd119,8'd209} : s = 28;
	{8'd119,8'd210} : s = 114;
	{8'd119,8'd211} : s = 113;
	{8'd119,8'd212} : s = 242;
	{8'd119,8'd213} : s = 108;
	{8'd119,8'd214} : s = 241;
	{8'd119,8'd215} : s = 236;
	{8'd119,8'd216} : s = 399;
	{8'd119,8'd217} : s = 26;
	{8'd119,8'd218} : s = 106;
	{8'd119,8'd219} : s = 105;
	{8'd119,8'd220} : s = 234;
	{8'd119,8'd221} : s = 102;
	{8'd119,8'd222} : s = 233;
	{8'd119,8'd223} : s = 230;
	{8'd119,8'd224} : s = 380;
	{8'd119,8'd225} : s = 101;
	{8'd119,8'd226} : s = 229;
	{8'd119,8'd227} : s = 227;
	{8'd119,8'd228} : s = 378;
	{8'd119,8'd229} : s = 220;
	{8'd119,8'd230} : s = 377;
	{8'd119,8'd231} : s = 374;
	{8'd119,8'd232} : s = 487;
	{8'd119,8'd233} : s = 25;
	{8'd119,8'd234} : s = 99;
	{8'd119,8'd235} : s = 92;
	{8'd119,8'd236} : s = 218;
	{8'd119,8'd237} : s = 90;
	{8'd119,8'd238} : s = 217;
	{8'd119,8'd239} : s = 214;
	{8'd119,8'd240} : s = 373;
	{8'd119,8'd241} : s = 89;
	{8'd119,8'd242} : s = 213;
	{8'd119,8'd243} : s = 211;
	{8'd119,8'd244} : s = 371;
	{8'd119,8'd245} : s = 206;
	{8'd119,8'd246} : s = 366;
	{8'd119,8'd247} : s = 365;
	{8'd119,8'd248} : s = 478;
	{8'd119,8'd249} : s = 86;
	{8'd119,8'd250} : s = 205;
	{8'd119,8'd251} : s = 203;
	{8'd119,8'd252} : s = 363;
	{8'd119,8'd253} : s = 199;
	{8'd119,8'd254} : s = 359;
	{8'd119,8'd255} : s = 350;
	{8'd120,8'd0} : s = 325;
	{8'd120,8'd1} : s = 433;
	{8'd120,8'd2} : s = 428;
	{8'd120,8'd3} : s = 492;
	{8'd120,8'd4} : s = 426;
	{8'd120,8'd5} : s = 490;
	{8'd120,8'd6} : s = 489;
	{8'd120,8'd7} : s = 508;
	{8'd120,8'd8} : s = 2;
	{8'd120,8'd9} : s = 48;
	{8'd120,8'd10} : s = 40;
	{8'd120,8'd11} : s = 168;
	{8'd120,8'd12} : s = 36;
	{8'd120,8'd13} : s = 164;
	{8'd120,8'd14} : s = 162;
	{8'd120,8'd15} : s = 323;
	{8'd120,8'd16} : s = 34;
	{8'd120,8'd17} : s = 161;
	{8'd120,8'd18} : s = 152;
	{8'd120,8'd19} : s = 312;
	{8'd120,8'd20} : s = 148;
	{8'd120,8'd21} : s = 308;
	{8'd120,8'd22} : s = 306;
	{8'd120,8'd23} : s = 425;
	{8'd120,8'd24} : s = 33;
	{8'd120,8'd25} : s = 146;
	{8'd120,8'd26} : s = 145;
	{8'd120,8'd27} : s = 305;
	{8'd120,8'd28} : s = 140;
	{8'd120,8'd29} : s = 300;
	{8'd120,8'd30} : s = 298;
	{8'd120,8'd31} : s = 422;
	{8'd120,8'd32} : s = 138;
	{8'd120,8'd33} : s = 297;
	{8'd120,8'd34} : s = 294;
	{8'd120,8'd35} : s = 421;
	{8'd120,8'd36} : s = 293;
	{8'd120,8'd37} : s = 419;
	{8'd120,8'd38} : s = 412;
	{8'd120,8'd39} : s = 486;
	{8'd120,8'd40} : s = 24;
	{8'd120,8'd41} : s = 137;
	{8'd120,8'd42} : s = 134;
	{8'd120,8'd43} : s = 291;
	{8'd120,8'd44} : s = 133;
	{8'd120,8'd45} : s = 284;
	{8'd120,8'd46} : s = 282;
	{8'd120,8'd47} : s = 410;
	{8'd120,8'd48} : s = 131;
	{8'd120,8'd49} : s = 281;
	{8'd120,8'd50} : s = 278;
	{8'd120,8'd51} : s = 409;
	{8'd120,8'd52} : s = 277;
	{8'd120,8'd53} : s = 406;
	{8'd120,8'd54} : s = 405;
	{8'd120,8'd55} : s = 485;
	{8'd120,8'd56} : s = 112;
	{8'd120,8'd57} : s = 275;
	{8'd120,8'd58} : s = 270;
	{8'd120,8'd59} : s = 403;
	{8'd120,8'd60} : s = 269;
	{8'd120,8'd61} : s = 398;
	{8'd120,8'd62} : s = 397;
	{8'd120,8'd63} : s = 483;
	{8'd120,8'd64} : s = 267;
	{8'd120,8'd65} : s = 395;
	{8'd120,8'd66} : s = 391;
	{8'd120,8'd67} : s = 476;
	{8'd120,8'd68} : s = 376;
	{8'd120,8'd69} : s = 474;
	{8'd120,8'd70} : s = 473;
	{8'd120,8'd71} : s = 506;
	{8'd120,8'd72} : s = 20;
	{8'd120,8'd73} : s = 104;
	{8'd120,8'd74} : s = 100;
	{8'd120,8'd75} : s = 263;
	{8'd120,8'd76} : s = 98;
	{8'd120,8'd77} : s = 240;
	{8'd120,8'd78} : s = 232;
	{8'd120,8'd79} : s = 372;
	{8'd120,8'd80} : s = 97;
	{8'd120,8'd81} : s = 228;
	{8'd120,8'd82} : s = 226;
	{8'd120,8'd83} : s = 370;
	{8'd120,8'd84} : s = 225;
	{8'd120,8'd85} : s = 369;
	{8'd120,8'd86} : s = 364;
	{8'd120,8'd87} : s = 470;
	{8'd120,8'd88} : s = 88;
	{8'd120,8'd89} : s = 216;
	{8'd120,8'd90} : s = 212;
	{8'd120,8'd91} : s = 362;
	{8'd120,8'd92} : s = 210;
	{8'd120,8'd93} : s = 361;
	{8'd120,8'd94} : s = 358;
	{8'd120,8'd95} : s = 469;
	{8'd120,8'd96} : s = 209;
	{8'd120,8'd97} : s = 357;
	{8'd120,8'd98} : s = 355;
	{8'd120,8'd99} : s = 467;
	{8'd120,8'd100} : s = 348;
	{8'd120,8'd101} : s = 462;
	{8'd120,8'd102} : s = 461;
	{8'd120,8'd103} : s = 505;
	{8'd120,8'd104} : s = 84;
	{8'd120,8'd105} : s = 204;
	{8'd120,8'd106} : s = 202;
	{8'd120,8'd107} : s = 346;
	{8'd120,8'd108} : s = 201;
	{8'd120,8'd109} : s = 345;
	{8'd120,8'd110} : s = 342;
	{8'd120,8'd111} : s = 459;
	{8'd120,8'd112} : s = 198;
	{8'd120,8'd113} : s = 341;
	{8'd120,8'd114} : s = 339;
	{8'd120,8'd115} : s = 455;
	{8'd120,8'd116} : s = 334;
	{8'd120,8'd117} : s = 444;
	{8'd120,8'd118} : s = 442;
	{8'd120,8'd119} : s = 502;
	{8'd120,8'd120} : s = 197;
	{8'd120,8'd121} : s = 333;
	{8'd120,8'd122} : s = 331;
	{8'd120,8'd123} : s = 441;
	{8'd120,8'd124} : s = 327;
	{8'd120,8'd125} : s = 438;
	{8'd120,8'd126} : s = 437;
	{8'd120,8'd127} : s = 501;
	{8'd120,8'd128} : s = 316;
	{8'd120,8'd129} : s = 435;
	{8'd120,8'd130} : s = 430;
	{8'd120,8'd131} : s = 499;
	{8'd120,8'd132} : s = 429;
	{8'd120,8'd133} : s = 494;
	{8'd120,8'd134} : s = 493;
	{8'd120,8'd135} : s = 510;
	{8'd120,8'd136} : s = 1;
	{8'd120,8'd137} : s = 18;
	{8'd120,8'd138} : s = 17;
	{8'd120,8'd139} : s = 82;
	{8'd120,8'd140} : s = 12;
	{8'd120,8'd141} : s = 81;
	{8'd120,8'd142} : s = 76;
	{8'd120,8'd143} : s = 195;
	{8'd120,8'd144} : s = 10;
	{8'd120,8'd145} : s = 74;
	{8'd120,8'd146} : s = 73;
	{8'd120,8'd147} : s = 184;
	{8'd120,8'd148} : s = 70;
	{8'd120,8'd149} : s = 180;
	{8'd120,8'd150} : s = 178;
	{8'd120,8'd151} : s = 314;
	{8'd120,8'd152} : s = 9;
	{8'd120,8'd153} : s = 69;
	{8'd120,8'd154} : s = 67;
	{8'd120,8'd155} : s = 177;
	{8'd120,8'd156} : s = 56;
	{8'd120,8'd157} : s = 172;
	{8'd120,8'd158} : s = 170;
	{8'd120,8'd159} : s = 313;
	{8'd120,8'd160} : s = 52;
	{8'd120,8'd161} : s = 169;
	{8'd120,8'd162} : s = 166;
	{8'd120,8'd163} : s = 310;
	{8'd120,8'd164} : s = 165;
	{8'd120,8'd165} : s = 309;
	{8'd120,8'd166} : s = 307;
	{8'd120,8'd167} : s = 427;
	{8'd120,8'd168} : s = 6;
	{8'd120,8'd169} : s = 50;
	{8'd120,8'd170} : s = 49;
	{8'd120,8'd171} : s = 163;
	{8'd120,8'd172} : s = 44;
	{8'd120,8'd173} : s = 156;
	{8'd120,8'd174} : s = 154;
	{8'd120,8'd175} : s = 302;
	{8'd120,8'd176} : s = 42;
	{8'd120,8'd177} : s = 153;
	{8'd120,8'd178} : s = 150;
	{8'd120,8'd179} : s = 301;
	{8'd120,8'd180} : s = 149;
	{8'd120,8'd181} : s = 299;
	{8'd120,8'd182} : s = 295;
	{8'd120,8'd183} : s = 423;
	{8'd120,8'd184} : s = 41;
	{8'd120,8'd185} : s = 147;
	{8'd120,8'd186} : s = 142;
	{8'd120,8'd187} : s = 286;
	{8'd120,8'd188} : s = 141;
	{8'd120,8'd189} : s = 285;
	{8'd120,8'd190} : s = 283;
	{8'd120,8'd191} : s = 414;
	{8'd120,8'd192} : s = 139;
	{8'd120,8'd193} : s = 279;
	{8'd120,8'd194} : s = 271;
	{8'd120,8'd195} : s = 413;
	{8'd120,8'd196} : s = 248;
	{8'd120,8'd197} : s = 411;
	{8'd120,8'd198} : s = 407;
	{8'd120,8'd199} : s = 491;
	{8'd120,8'd200} : s = 5;
	{8'd120,8'd201} : s = 38;
	{8'd120,8'd202} : s = 37;
	{8'd120,8'd203} : s = 135;
	{8'd120,8'd204} : s = 35;
	{8'd120,8'd205} : s = 120;
	{8'd120,8'd206} : s = 116;
	{8'd120,8'd207} : s = 244;
	{8'd120,8'd208} : s = 28;
	{8'd120,8'd209} : s = 114;
	{8'd120,8'd210} : s = 113;
	{8'd120,8'd211} : s = 242;
	{8'd120,8'd212} : s = 108;
	{8'd120,8'd213} : s = 241;
	{8'd120,8'd214} : s = 236;
	{8'd120,8'd215} : s = 399;
	{8'd120,8'd216} : s = 26;
	{8'd120,8'd217} : s = 106;
	{8'd120,8'd218} : s = 105;
	{8'd120,8'd219} : s = 234;
	{8'd120,8'd220} : s = 102;
	{8'd120,8'd221} : s = 233;
	{8'd120,8'd222} : s = 230;
	{8'd120,8'd223} : s = 380;
	{8'd120,8'd224} : s = 101;
	{8'd120,8'd225} : s = 229;
	{8'd120,8'd226} : s = 227;
	{8'd120,8'd227} : s = 378;
	{8'd120,8'd228} : s = 220;
	{8'd120,8'd229} : s = 377;
	{8'd120,8'd230} : s = 374;
	{8'd120,8'd231} : s = 487;
	{8'd120,8'd232} : s = 25;
	{8'd120,8'd233} : s = 99;
	{8'd120,8'd234} : s = 92;
	{8'd120,8'd235} : s = 218;
	{8'd120,8'd236} : s = 90;
	{8'd120,8'd237} : s = 217;
	{8'd120,8'd238} : s = 214;
	{8'd120,8'd239} : s = 373;
	{8'd120,8'd240} : s = 89;
	{8'd120,8'd241} : s = 213;
	{8'd120,8'd242} : s = 211;
	{8'd120,8'd243} : s = 371;
	{8'd120,8'd244} : s = 206;
	{8'd120,8'd245} : s = 366;
	{8'd120,8'd246} : s = 365;
	{8'd120,8'd247} : s = 478;
	{8'd120,8'd248} : s = 86;
	{8'd120,8'd249} : s = 205;
	{8'd120,8'd250} : s = 203;
	{8'd120,8'd251} : s = 363;
	{8'd120,8'd252} : s = 199;
	{8'd120,8'd253} : s = 359;
	{8'd120,8'd254} : s = 350;
	{8'd120,8'd255} : s = 477;
	{8'd121,8'd0} : s = 433;
	{8'd121,8'd1} : s = 428;
	{8'd121,8'd2} : s = 492;
	{8'd121,8'd3} : s = 426;
	{8'd121,8'd4} : s = 490;
	{8'd121,8'd5} : s = 489;
	{8'd121,8'd6} : s = 508;
	{8'd121,8'd7} : s = 2;
	{8'd121,8'd8} : s = 48;
	{8'd121,8'd9} : s = 40;
	{8'd121,8'd10} : s = 168;
	{8'd121,8'd11} : s = 36;
	{8'd121,8'd12} : s = 164;
	{8'd121,8'd13} : s = 162;
	{8'd121,8'd14} : s = 323;
	{8'd121,8'd15} : s = 34;
	{8'd121,8'd16} : s = 161;
	{8'd121,8'd17} : s = 152;
	{8'd121,8'd18} : s = 312;
	{8'd121,8'd19} : s = 148;
	{8'd121,8'd20} : s = 308;
	{8'd121,8'd21} : s = 306;
	{8'd121,8'd22} : s = 425;
	{8'd121,8'd23} : s = 33;
	{8'd121,8'd24} : s = 146;
	{8'd121,8'd25} : s = 145;
	{8'd121,8'd26} : s = 305;
	{8'd121,8'd27} : s = 140;
	{8'd121,8'd28} : s = 300;
	{8'd121,8'd29} : s = 298;
	{8'd121,8'd30} : s = 422;
	{8'd121,8'd31} : s = 138;
	{8'd121,8'd32} : s = 297;
	{8'd121,8'd33} : s = 294;
	{8'd121,8'd34} : s = 421;
	{8'd121,8'd35} : s = 293;
	{8'd121,8'd36} : s = 419;
	{8'd121,8'd37} : s = 412;
	{8'd121,8'd38} : s = 486;
	{8'd121,8'd39} : s = 24;
	{8'd121,8'd40} : s = 137;
	{8'd121,8'd41} : s = 134;
	{8'd121,8'd42} : s = 291;
	{8'd121,8'd43} : s = 133;
	{8'd121,8'd44} : s = 284;
	{8'd121,8'd45} : s = 282;
	{8'd121,8'd46} : s = 410;
	{8'd121,8'd47} : s = 131;
	{8'd121,8'd48} : s = 281;
	{8'd121,8'd49} : s = 278;
	{8'd121,8'd50} : s = 409;
	{8'd121,8'd51} : s = 277;
	{8'd121,8'd52} : s = 406;
	{8'd121,8'd53} : s = 405;
	{8'd121,8'd54} : s = 485;
	{8'd121,8'd55} : s = 112;
	{8'd121,8'd56} : s = 275;
	{8'd121,8'd57} : s = 270;
	{8'd121,8'd58} : s = 403;
	{8'd121,8'd59} : s = 269;
	{8'd121,8'd60} : s = 398;
	{8'd121,8'd61} : s = 397;
	{8'd121,8'd62} : s = 483;
	{8'd121,8'd63} : s = 267;
	{8'd121,8'd64} : s = 395;
	{8'd121,8'd65} : s = 391;
	{8'd121,8'd66} : s = 476;
	{8'd121,8'd67} : s = 376;
	{8'd121,8'd68} : s = 474;
	{8'd121,8'd69} : s = 473;
	{8'd121,8'd70} : s = 506;
	{8'd121,8'd71} : s = 20;
	{8'd121,8'd72} : s = 104;
	{8'd121,8'd73} : s = 100;
	{8'd121,8'd74} : s = 263;
	{8'd121,8'd75} : s = 98;
	{8'd121,8'd76} : s = 240;
	{8'd121,8'd77} : s = 232;
	{8'd121,8'd78} : s = 372;
	{8'd121,8'd79} : s = 97;
	{8'd121,8'd80} : s = 228;
	{8'd121,8'd81} : s = 226;
	{8'd121,8'd82} : s = 370;
	{8'd121,8'd83} : s = 225;
	{8'd121,8'd84} : s = 369;
	{8'd121,8'd85} : s = 364;
	{8'd121,8'd86} : s = 470;
	{8'd121,8'd87} : s = 88;
	{8'd121,8'd88} : s = 216;
	{8'd121,8'd89} : s = 212;
	{8'd121,8'd90} : s = 362;
	{8'd121,8'd91} : s = 210;
	{8'd121,8'd92} : s = 361;
	{8'd121,8'd93} : s = 358;
	{8'd121,8'd94} : s = 469;
	{8'd121,8'd95} : s = 209;
	{8'd121,8'd96} : s = 357;
	{8'd121,8'd97} : s = 355;
	{8'd121,8'd98} : s = 467;
	{8'd121,8'd99} : s = 348;
	{8'd121,8'd100} : s = 462;
	{8'd121,8'd101} : s = 461;
	{8'd121,8'd102} : s = 505;
	{8'd121,8'd103} : s = 84;
	{8'd121,8'd104} : s = 204;
	{8'd121,8'd105} : s = 202;
	{8'd121,8'd106} : s = 346;
	{8'd121,8'd107} : s = 201;
	{8'd121,8'd108} : s = 345;
	{8'd121,8'd109} : s = 342;
	{8'd121,8'd110} : s = 459;
	{8'd121,8'd111} : s = 198;
	{8'd121,8'd112} : s = 341;
	{8'd121,8'd113} : s = 339;
	{8'd121,8'd114} : s = 455;
	{8'd121,8'd115} : s = 334;
	{8'd121,8'd116} : s = 444;
	{8'd121,8'd117} : s = 442;
	{8'd121,8'd118} : s = 502;
	{8'd121,8'd119} : s = 197;
	{8'd121,8'd120} : s = 333;
	{8'd121,8'd121} : s = 331;
	{8'd121,8'd122} : s = 441;
	{8'd121,8'd123} : s = 327;
	{8'd121,8'd124} : s = 438;
	{8'd121,8'd125} : s = 437;
	{8'd121,8'd126} : s = 501;
	{8'd121,8'd127} : s = 316;
	{8'd121,8'd128} : s = 435;
	{8'd121,8'd129} : s = 430;
	{8'd121,8'd130} : s = 499;
	{8'd121,8'd131} : s = 429;
	{8'd121,8'd132} : s = 494;
	{8'd121,8'd133} : s = 493;
	{8'd121,8'd134} : s = 510;
	{8'd121,8'd135} : s = 1;
	{8'd121,8'd136} : s = 18;
	{8'd121,8'd137} : s = 17;
	{8'd121,8'd138} : s = 82;
	{8'd121,8'd139} : s = 12;
	{8'd121,8'd140} : s = 81;
	{8'd121,8'd141} : s = 76;
	{8'd121,8'd142} : s = 195;
	{8'd121,8'd143} : s = 10;
	{8'd121,8'd144} : s = 74;
	{8'd121,8'd145} : s = 73;
	{8'd121,8'd146} : s = 184;
	{8'd121,8'd147} : s = 70;
	{8'd121,8'd148} : s = 180;
	{8'd121,8'd149} : s = 178;
	{8'd121,8'd150} : s = 314;
	{8'd121,8'd151} : s = 9;
	{8'd121,8'd152} : s = 69;
	{8'd121,8'd153} : s = 67;
	{8'd121,8'd154} : s = 177;
	{8'd121,8'd155} : s = 56;
	{8'd121,8'd156} : s = 172;
	{8'd121,8'd157} : s = 170;
	{8'd121,8'd158} : s = 313;
	{8'd121,8'd159} : s = 52;
	{8'd121,8'd160} : s = 169;
	{8'd121,8'd161} : s = 166;
	{8'd121,8'd162} : s = 310;
	{8'd121,8'd163} : s = 165;
	{8'd121,8'd164} : s = 309;
	{8'd121,8'd165} : s = 307;
	{8'd121,8'd166} : s = 427;
	{8'd121,8'd167} : s = 6;
	{8'd121,8'd168} : s = 50;
	{8'd121,8'd169} : s = 49;
	{8'd121,8'd170} : s = 163;
	{8'd121,8'd171} : s = 44;
	{8'd121,8'd172} : s = 156;
	{8'd121,8'd173} : s = 154;
	{8'd121,8'd174} : s = 302;
	{8'd121,8'd175} : s = 42;
	{8'd121,8'd176} : s = 153;
	{8'd121,8'd177} : s = 150;
	{8'd121,8'd178} : s = 301;
	{8'd121,8'd179} : s = 149;
	{8'd121,8'd180} : s = 299;
	{8'd121,8'd181} : s = 295;
	{8'd121,8'd182} : s = 423;
	{8'd121,8'd183} : s = 41;
	{8'd121,8'd184} : s = 147;
	{8'd121,8'd185} : s = 142;
	{8'd121,8'd186} : s = 286;
	{8'd121,8'd187} : s = 141;
	{8'd121,8'd188} : s = 285;
	{8'd121,8'd189} : s = 283;
	{8'd121,8'd190} : s = 414;
	{8'd121,8'd191} : s = 139;
	{8'd121,8'd192} : s = 279;
	{8'd121,8'd193} : s = 271;
	{8'd121,8'd194} : s = 413;
	{8'd121,8'd195} : s = 248;
	{8'd121,8'd196} : s = 411;
	{8'd121,8'd197} : s = 407;
	{8'd121,8'd198} : s = 491;
	{8'd121,8'd199} : s = 5;
	{8'd121,8'd200} : s = 38;
	{8'd121,8'd201} : s = 37;
	{8'd121,8'd202} : s = 135;
	{8'd121,8'd203} : s = 35;
	{8'd121,8'd204} : s = 120;
	{8'd121,8'd205} : s = 116;
	{8'd121,8'd206} : s = 244;
	{8'd121,8'd207} : s = 28;
	{8'd121,8'd208} : s = 114;
	{8'd121,8'd209} : s = 113;
	{8'd121,8'd210} : s = 242;
	{8'd121,8'd211} : s = 108;
	{8'd121,8'd212} : s = 241;
	{8'd121,8'd213} : s = 236;
	{8'd121,8'd214} : s = 399;
	{8'd121,8'd215} : s = 26;
	{8'd121,8'd216} : s = 106;
	{8'd121,8'd217} : s = 105;
	{8'd121,8'd218} : s = 234;
	{8'd121,8'd219} : s = 102;
	{8'd121,8'd220} : s = 233;
	{8'd121,8'd221} : s = 230;
	{8'd121,8'd222} : s = 380;
	{8'd121,8'd223} : s = 101;
	{8'd121,8'd224} : s = 229;
	{8'd121,8'd225} : s = 227;
	{8'd121,8'd226} : s = 378;
	{8'd121,8'd227} : s = 220;
	{8'd121,8'd228} : s = 377;
	{8'd121,8'd229} : s = 374;
	{8'd121,8'd230} : s = 487;
	{8'd121,8'd231} : s = 25;
	{8'd121,8'd232} : s = 99;
	{8'd121,8'd233} : s = 92;
	{8'd121,8'd234} : s = 218;
	{8'd121,8'd235} : s = 90;
	{8'd121,8'd236} : s = 217;
	{8'd121,8'd237} : s = 214;
	{8'd121,8'd238} : s = 373;
	{8'd121,8'd239} : s = 89;
	{8'd121,8'd240} : s = 213;
	{8'd121,8'd241} : s = 211;
	{8'd121,8'd242} : s = 371;
	{8'd121,8'd243} : s = 206;
	{8'd121,8'd244} : s = 366;
	{8'd121,8'd245} : s = 365;
	{8'd121,8'd246} : s = 478;
	{8'd121,8'd247} : s = 86;
	{8'd121,8'd248} : s = 205;
	{8'd121,8'd249} : s = 203;
	{8'd121,8'd250} : s = 363;
	{8'd121,8'd251} : s = 199;
	{8'd121,8'd252} : s = 359;
	{8'd121,8'd253} : s = 350;
	{8'd121,8'd254} : s = 477;
	{8'd121,8'd255} : s = 188;
	{8'd122,8'd0} : s = 428;
	{8'd122,8'd1} : s = 492;
	{8'd122,8'd2} : s = 426;
	{8'd122,8'd3} : s = 490;
	{8'd122,8'd4} : s = 489;
	{8'd122,8'd5} : s = 508;
	{8'd122,8'd6} : s = 2;
	{8'd122,8'd7} : s = 48;
	{8'd122,8'd8} : s = 40;
	{8'd122,8'd9} : s = 168;
	{8'd122,8'd10} : s = 36;
	{8'd122,8'd11} : s = 164;
	{8'd122,8'd12} : s = 162;
	{8'd122,8'd13} : s = 323;
	{8'd122,8'd14} : s = 34;
	{8'd122,8'd15} : s = 161;
	{8'd122,8'd16} : s = 152;
	{8'd122,8'd17} : s = 312;
	{8'd122,8'd18} : s = 148;
	{8'd122,8'd19} : s = 308;
	{8'd122,8'd20} : s = 306;
	{8'd122,8'd21} : s = 425;
	{8'd122,8'd22} : s = 33;
	{8'd122,8'd23} : s = 146;
	{8'd122,8'd24} : s = 145;
	{8'd122,8'd25} : s = 305;
	{8'd122,8'd26} : s = 140;
	{8'd122,8'd27} : s = 300;
	{8'd122,8'd28} : s = 298;
	{8'd122,8'd29} : s = 422;
	{8'd122,8'd30} : s = 138;
	{8'd122,8'd31} : s = 297;
	{8'd122,8'd32} : s = 294;
	{8'd122,8'd33} : s = 421;
	{8'd122,8'd34} : s = 293;
	{8'd122,8'd35} : s = 419;
	{8'd122,8'd36} : s = 412;
	{8'd122,8'd37} : s = 486;
	{8'd122,8'd38} : s = 24;
	{8'd122,8'd39} : s = 137;
	{8'd122,8'd40} : s = 134;
	{8'd122,8'd41} : s = 291;
	{8'd122,8'd42} : s = 133;
	{8'd122,8'd43} : s = 284;
	{8'd122,8'd44} : s = 282;
	{8'd122,8'd45} : s = 410;
	{8'd122,8'd46} : s = 131;
	{8'd122,8'd47} : s = 281;
	{8'd122,8'd48} : s = 278;
	{8'd122,8'd49} : s = 409;
	{8'd122,8'd50} : s = 277;
	{8'd122,8'd51} : s = 406;
	{8'd122,8'd52} : s = 405;
	{8'd122,8'd53} : s = 485;
	{8'd122,8'd54} : s = 112;
	{8'd122,8'd55} : s = 275;
	{8'd122,8'd56} : s = 270;
	{8'd122,8'd57} : s = 403;
	{8'd122,8'd58} : s = 269;
	{8'd122,8'd59} : s = 398;
	{8'd122,8'd60} : s = 397;
	{8'd122,8'd61} : s = 483;
	{8'd122,8'd62} : s = 267;
	{8'd122,8'd63} : s = 395;
	{8'd122,8'd64} : s = 391;
	{8'd122,8'd65} : s = 476;
	{8'd122,8'd66} : s = 376;
	{8'd122,8'd67} : s = 474;
	{8'd122,8'd68} : s = 473;
	{8'd122,8'd69} : s = 506;
	{8'd122,8'd70} : s = 20;
	{8'd122,8'd71} : s = 104;
	{8'd122,8'd72} : s = 100;
	{8'd122,8'd73} : s = 263;
	{8'd122,8'd74} : s = 98;
	{8'd122,8'd75} : s = 240;
	{8'd122,8'd76} : s = 232;
	{8'd122,8'd77} : s = 372;
	{8'd122,8'd78} : s = 97;
	{8'd122,8'd79} : s = 228;
	{8'd122,8'd80} : s = 226;
	{8'd122,8'd81} : s = 370;
	{8'd122,8'd82} : s = 225;
	{8'd122,8'd83} : s = 369;
	{8'd122,8'd84} : s = 364;
	{8'd122,8'd85} : s = 470;
	{8'd122,8'd86} : s = 88;
	{8'd122,8'd87} : s = 216;
	{8'd122,8'd88} : s = 212;
	{8'd122,8'd89} : s = 362;
	{8'd122,8'd90} : s = 210;
	{8'd122,8'd91} : s = 361;
	{8'd122,8'd92} : s = 358;
	{8'd122,8'd93} : s = 469;
	{8'd122,8'd94} : s = 209;
	{8'd122,8'd95} : s = 357;
	{8'd122,8'd96} : s = 355;
	{8'd122,8'd97} : s = 467;
	{8'd122,8'd98} : s = 348;
	{8'd122,8'd99} : s = 462;
	{8'd122,8'd100} : s = 461;
	{8'd122,8'd101} : s = 505;
	{8'd122,8'd102} : s = 84;
	{8'd122,8'd103} : s = 204;
	{8'd122,8'd104} : s = 202;
	{8'd122,8'd105} : s = 346;
	{8'd122,8'd106} : s = 201;
	{8'd122,8'd107} : s = 345;
	{8'd122,8'd108} : s = 342;
	{8'd122,8'd109} : s = 459;
	{8'd122,8'd110} : s = 198;
	{8'd122,8'd111} : s = 341;
	{8'd122,8'd112} : s = 339;
	{8'd122,8'd113} : s = 455;
	{8'd122,8'd114} : s = 334;
	{8'd122,8'd115} : s = 444;
	{8'd122,8'd116} : s = 442;
	{8'd122,8'd117} : s = 502;
	{8'd122,8'd118} : s = 197;
	{8'd122,8'd119} : s = 333;
	{8'd122,8'd120} : s = 331;
	{8'd122,8'd121} : s = 441;
	{8'd122,8'd122} : s = 327;
	{8'd122,8'd123} : s = 438;
	{8'd122,8'd124} : s = 437;
	{8'd122,8'd125} : s = 501;
	{8'd122,8'd126} : s = 316;
	{8'd122,8'd127} : s = 435;
	{8'd122,8'd128} : s = 430;
	{8'd122,8'd129} : s = 499;
	{8'd122,8'd130} : s = 429;
	{8'd122,8'd131} : s = 494;
	{8'd122,8'd132} : s = 493;
	{8'd122,8'd133} : s = 510;
	{8'd122,8'd134} : s = 1;
	{8'd122,8'd135} : s = 18;
	{8'd122,8'd136} : s = 17;
	{8'd122,8'd137} : s = 82;
	{8'd122,8'd138} : s = 12;
	{8'd122,8'd139} : s = 81;
	{8'd122,8'd140} : s = 76;
	{8'd122,8'd141} : s = 195;
	{8'd122,8'd142} : s = 10;
	{8'd122,8'd143} : s = 74;
	{8'd122,8'd144} : s = 73;
	{8'd122,8'd145} : s = 184;
	{8'd122,8'd146} : s = 70;
	{8'd122,8'd147} : s = 180;
	{8'd122,8'd148} : s = 178;
	{8'd122,8'd149} : s = 314;
	{8'd122,8'd150} : s = 9;
	{8'd122,8'd151} : s = 69;
	{8'd122,8'd152} : s = 67;
	{8'd122,8'd153} : s = 177;
	{8'd122,8'd154} : s = 56;
	{8'd122,8'd155} : s = 172;
	{8'd122,8'd156} : s = 170;
	{8'd122,8'd157} : s = 313;
	{8'd122,8'd158} : s = 52;
	{8'd122,8'd159} : s = 169;
	{8'd122,8'd160} : s = 166;
	{8'd122,8'd161} : s = 310;
	{8'd122,8'd162} : s = 165;
	{8'd122,8'd163} : s = 309;
	{8'd122,8'd164} : s = 307;
	{8'd122,8'd165} : s = 427;
	{8'd122,8'd166} : s = 6;
	{8'd122,8'd167} : s = 50;
	{8'd122,8'd168} : s = 49;
	{8'd122,8'd169} : s = 163;
	{8'd122,8'd170} : s = 44;
	{8'd122,8'd171} : s = 156;
	{8'd122,8'd172} : s = 154;
	{8'd122,8'd173} : s = 302;
	{8'd122,8'd174} : s = 42;
	{8'd122,8'd175} : s = 153;
	{8'd122,8'd176} : s = 150;
	{8'd122,8'd177} : s = 301;
	{8'd122,8'd178} : s = 149;
	{8'd122,8'd179} : s = 299;
	{8'd122,8'd180} : s = 295;
	{8'd122,8'd181} : s = 423;
	{8'd122,8'd182} : s = 41;
	{8'd122,8'd183} : s = 147;
	{8'd122,8'd184} : s = 142;
	{8'd122,8'd185} : s = 286;
	{8'd122,8'd186} : s = 141;
	{8'd122,8'd187} : s = 285;
	{8'd122,8'd188} : s = 283;
	{8'd122,8'd189} : s = 414;
	{8'd122,8'd190} : s = 139;
	{8'd122,8'd191} : s = 279;
	{8'd122,8'd192} : s = 271;
	{8'd122,8'd193} : s = 413;
	{8'd122,8'd194} : s = 248;
	{8'd122,8'd195} : s = 411;
	{8'd122,8'd196} : s = 407;
	{8'd122,8'd197} : s = 491;
	{8'd122,8'd198} : s = 5;
	{8'd122,8'd199} : s = 38;
	{8'd122,8'd200} : s = 37;
	{8'd122,8'd201} : s = 135;
	{8'd122,8'd202} : s = 35;
	{8'd122,8'd203} : s = 120;
	{8'd122,8'd204} : s = 116;
	{8'd122,8'd205} : s = 244;
	{8'd122,8'd206} : s = 28;
	{8'd122,8'd207} : s = 114;
	{8'd122,8'd208} : s = 113;
	{8'd122,8'd209} : s = 242;
	{8'd122,8'd210} : s = 108;
	{8'd122,8'd211} : s = 241;
	{8'd122,8'd212} : s = 236;
	{8'd122,8'd213} : s = 399;
	{8'd122,8'd214} : s = 26;
	{8'd122,8'd215} : s = 106;
	{8'd122,8'd216} : s = 105;
	{8'd122,8'd217} : s = 234;
	{8'd122,8'd218} : s = 102;
	{8'd122,8'd219} : s = 233;
	{8'd122,8'd220} : s = 230;
	{8'd122,8'd221} : s = 380;
	{8'd122,8'd222} : s = 101;
	{8'd122,8'd223} : s = 229;
	{8'd122,8'd224} : s = 227;
	{8'd122,8'd225} : s = 378;
	{8'd122,8'd226} : s = 220;
	{8'd122,8'd227} : s = 377;
	{8'd122,8'd228} : s = 374;
	{8'd122,8'd229} : s = 487;
	{8'd122,8'd230} : s = 25;
	{8'd122,8'd231} : s = 99;
	{8'd122,8'd232} : s = 92;
	{8'd122,8'd233} : s = 218;
	{8'd122,8'd234} : s = 90;
	{8'd122,8'd235} : s = 217;
	{8'd122,8'd236} : s = 214;
	{8'd122,8'd237} : s = 373;
	{8'd122,8'd238} : s = 89;
	{8'd122,8'd239} : s = 213;
	{8'd122,8'd240} : s = 211;
	{8'd122,8'd241} : s = 371;
	{8'd122,8'd242} : s = 206;
	{8'd122,8'd243} : s = 366;
	{8'd122,8'd244} : s = 365;
	{8'd122,8'd245} : s = 478;
	{8'd122,8'd246} : s = 86;
	{8'd122,8'd247} : s = 205;
	{8'd122,8'd248} : s = 203;
	{8'd122,8'd249} : s = 363;
	{8'd122,8'd250} : s = 199;
	{8'd122,8'd251} : s = 359;
	{8'd122,8'd252} : s = 350;
	{8'd122,8'd253} : s = 477;
	{8'd122,8'd254} : s = 188;
	{8'd122,8'd255} : s = 349;
	{8'd123,8'd0} : s = 492;
	{8'd123,8'd1} : s = 426;
	{8'd123,8'd2} : s = 490;
	{8'd123,8'd3} : s = 489;
	{8'd123,8'd4} : s = 508;
	{8'd123,8'd5} : s = 2;
	{8'd123,8'd6} : s = 48;
	{8'd123,8'd7} : s = 40;
	{8'd123,8'd8} : s = 168;
	{8'd123,8'd9} : s = 36;
	{8'd123,8'd10} : s = 164;
	{8'd123,8'd11} : s = 162;
	{8'd123,8'd12} : s = 323;
	{8'd123,8'd13} : s = 34;
	{8'd123,8'd14} : s = 161;
	{8'd123,8'd15} : s = 152;
	{8'd123,8'd16} : s = 312;
	{8'd123,8'd17} : s = 148;
	{8'd123,8'd18} : s = 308;
	{8'd123,8'd19} : s = 306;
	{8'd123,8'd20} : s = 425;
	{8'd123,8'd21} : s = 33;
	{8'd123,8'd22} : s = 146;
	{8'd123,8'd23} : s = 145;
	{8'd123,8'd24} : s = 305;
	{8'd123,8'd25} : s = 140;
	{8'd123,8'd26} : s = 300;
	{8'd123,8'd27} : s = 298;
	{8'd123,8'd28} : s = 422;
	{8'd123,8'd29} : s = 138;
	{8'd123,8'd30} : s = 297;
	{8'd123,8'd31} : s = 294;
	{8'd123,8'd32} : s = 421;
	{8'd123,8'd33} : s = 293;
	{8'd123,8'd34} : s = 419;
	{8'd123,8'd35} : s = 412;
	{8'd123,8'd36} : s = 486;
	{8'd123,8'd37} : s = 24;
	{8'd123,8'd38} : s = 137;
	{8'd123,8'd39} : s = 134;
	{8'd123,8'd40} : s = 291;
	{8'd123,8'd41} : s = 133;
	{8'd123,8'd42} : s = 284;
	{8'd123,8'd43} : s = 282;
	{8'd123,8'd44} : s = 410;
	{8'd123,8'd45} : s = 131;
	{8'd123,8'd46} : s = 281;
	{8'd123,8'd47} : s = 278;
	{8'd123,8'd48} : s = 409;
	{8'd123,8'd49} : s = 277;
	{8'd123,8'd50} : s = 406;
	{8'd123,8'd51} : s = 405;
	{8'd123,8'd52} : s = 485;
	{8'd123,8'd53} : s = 112;
	{8'd123,8'd54} : s = 275;
	{8'd123,8'd55} : s = 270;
	{8'd123,8'd56} : s = 403;
	{8'd123,8'd57} : s = 269;
	{8'd123,8'd58} : s = 398;
	{8'd123,8'd59} : s = 397;
	{8'd123,8'd60} : s = 483;
	{8'd123,8'd61} : s = 267;
	{8'd123,8'd62} : s = 395;
	{8'd123,8'd63} : s = 391;
	{8'd123,8'd64} : s = 476;
	{8'd123,8'd65} : s = 376;
	{8'd123,8'd66} : s = 474;
	{8'd123,8'd67} : s = 473;
	{8'd123,8'd68} : s = 506;
	{8'd123,8'd69} : s = 20;
	{8'd123,8'd70} : s = 104;
	{8'd123,8'd71} : s = 100;
	{8'd123,8'd72} : s = 263;
	{8'd123,8'd73} : s = 98;
	{8'd123,8'd74} : s = 240;
	{8'd123,8'd75} : s = 232;
	{8'd123,8'd76} : s = 372;
	{8'd123,8'd77} : s = 97;
	{8'd123,8'd78} : s = 228;
	{8'd123,8'd79} : s = 226;
	{8'd123,8'd80} : s = 370;
	{8'd123,8'd81} : s = 225;
	{8'd123,8'd82} : s = 369;
	{8'd123,8'd83} : s = 364;
	{8'd123,8'd84} : s = 470;
	{8'd123,8'd85} : s = 88;
	{8'd123,8'd86} : s = 216;
	{8'd123,8'd87} : s = 212;
	{8'd123,8'd88} : s = 362;
	{8'd123,8'd89} : s = 210;
	{8'd123,8'd90} : s = 361;
	{8'd123,8'd91} : s = 358;
	{8'd123,8'd92} : s = 469;
	{8'd123,8'd93} : s = 209;
	{8'd123,8'd94} : s = 357;
	{8'd123,8'd95} : s = 355;
	{8'd123,8'd96} : s = 467;
	{8'd123,8'd97} : s = 348;
	{8'd123,8'd98} : s = 462;
	{8'd123,8'd99} : s = 461;
	{8'd123,8'd100} : s = 505;
	{8'd123,8'd101} : s = 84;
	{8'd123,8'd102} : s = 204;
	{8'd123,8'd103} : s = 202;
	{8'd123,8'd104} : s = 346;
	{8'd123,8'd105} : s = 201;
	{8'd123,8'd106} : s = 345;
	{8'd123,8'd107} : s = 342;
	{8'd123,8'd108} : s = 459;
	{8'd123,8'd109} : s = 198;
	{8'd123,8'd110} : s = 341;
	{8'd123,8'd111} : s = 339;
	{8'd123,8'd112} : s = 455;
	{8'd123,8'd113} : s = 334;
	{8'd123,8'd114} : s = 444;
	{8'd123,8'd115} : s = 442;
	{8'd123,8'd116} : s = 502;
	{8'd123,8'd117} : s = 197;
	{8'd123,8'd118} : s = 333;
	{8'd123,8'd119} : s = 331;
	{8'd123,8'd120} : s = 441;
	{8'd123,8'd121} : s = 327;
	{8'd123,8'd122} : s = 438;
	{8'd123,8'd123} : s = 437;
	{8'd123,8'd124} : s = 501;
	{8'd123,8'd125} : s = 316;
	{8'd123,8'd126} : s = 435;
	{8'd123,8'd127} : s = 430;
	{8'd123,8'd128} : s = 499;
	{8'd123,8'd129} : s = 429;
	{8'd123,8'd130} : s = 494;
	{8'd123,8'd131} : s = 493;
	{8'd123,8'd132} : s = 510;
	{8'd123,8'd133} : s = 1;
	{8'd123,8'd134} : s = 18;
	{8'd123,8'd135} : s = 17;
	{8'd123,8'd136} : s = 82;
	{8'd123,8'd137} : s = 12;
	{8'd123,8'd138} : s = 81;
	{8'd123,8'd139} : s = 76;
	{8'd123,8'd140} : s = 195;
	{8'd123,8'd141} : s = 10;
	{8'd123,8'd142} : s = 74;
	{8'd123,8'd143} : s = 73;
	{8'd123,8'd144} : s = 184;
	{8'd123,8'd145} : s = 70;
	{8'd123,8'd146} : s = 180;
	{8'd123,8'd147} : s = 178;
	{8'd123,8'd148} : s = 314;
	{8'd123,8'd149} : s = 9;
	{8'd123,8'd150} : s = 69;
	{8'd123,8'd151} : s = 67;
	{8'd123,8'd152} : s = 177;
	{8'd123,8'd153} : s = 56;
	{8'd123,8'd154} : s = 172;
	{8'd123,8'd155} : s = 170;
	{8'd123,8'd156} : s = 313;
	{8'd123,8'd157} : s = 52;
	{8'd123,8'd158} : s = 169;
	{8'd123,8'd159} : s = 166;
	{8'd123,8'd160} : s = 310;
	{8'd123,8'd161} : s = 165;
	{8'd123,8'd162} : s = 309;
	{8'd123,8'd163} : s = 307;
	{8'd123,8'd164} : s = 427;
	{8'd123,8'd165} : s = 6;
	{8'd123,8'd166} : s = 50;
	{8'd123,8'd167} : s = 49;
	{8'd123,8'd168} : s = 163;
	{8'd123,8'd169} : s = 44;
	{8'd123,8'd170} : s = 156;
	{8'd123,8'd171} : s = 154;
	{8'd123,8'd172} : s = 302;
	{8'd123,8'd173} : s = 42;
	{8'd123,8'd174} : s = 153;
	{8'd123,8'd175} : s = 150;
	{8'd123,8'd176} : s = 301;
	{8'd123,8'd177} : s = 149;
	{8'd123,8'd178} : s = 299;
	{8'd123,8'd179} : s = 295;
	{8'd123,8'd180} : s = 423;
	{8'd123,8'd181} : s = 41;
	{8'd123,8'd182} : s = 147;
	{8'd123,8'd183} : s = 142;
	{8'd123,8'd184} : s = 286;
	{8'd123,8'd185} : s = 141;
	{8'd123,8'd186} : s = 285;
	{8'd123,8'd187} : s = 283;
	{8'd123,8'd188} : s = 414;
	{8'd123,8'd189} : s = 139;
	{8'd123,8'd190} : s = 279;
	{8'd123,8'd191} : s = 271;
	{8'd123,8'd192} : s = 413;
	{8'd123,8'd193} : s = 248;
	{8'd123,8'd194} : s = 411;
	{8'd123,8'd195} : s = 407;
	{8'd123,8'd196} : s = 491;
	{8'd123,8'd197} : s = 5;
	{8'd123,8'd198} : s = 38;
	{8'd123,8'd199} : s = 37;
	{8'd123,8'd200} : s = 135;
	{8'd123,8'd201} : s = 35;
	{8'd123,8'd202} : s = 120;
	{8'd123,8'd203} : s = 116;
	{8'd123,8'd204} : s = 244;
	{8'd123,8'd205} : s = 28;
	{8'd123,8'd206} : s = 114;
	{8'd123,8'd207} : s = 113;
	{8'd123,8'd208} : s = 242;
	{8'd123,8'd209} : s = 108;
	{8'd123,8'd210} : s = 241;
	{8'd123,8'd211} : s = 236;
	{8'd123,8'd212} : s = 399;
	{8'd123,8'd213} : s = 26;
	{8'd123,8'd214} : s = 106;
	{8'd123,8'd215} : s = 105;
	{8'd123,8'd216} : s = 234;
	{8'd123,8'd217} : s = 102;
	{8'd123,8'd218} : s = 233;
	{8'd123,8'd219} : s = 230;
	{8'd123,8'd220} : s = 380;
	{8'd123,8'd221} : s = 101;
	{8'd123,8'd222} : s = 229;
	{8'd123,8'd223} : s = 227;
	{8'd123,8'd224} : s = 378;
	{8'd123,8'd225} : s = 220;
	{8'd123,8'd226} : s = 377;
	{8'd123,8'd227} : s = 374;
	{8'd123,8'd228} : s = 487;
	{8'd123,8'd229} : s = 25;
	{8'd123,8'd230} : s = 99;
	{8'd123,8'd231} : s = 92;
	{8'd123,8'd232} : s = 218;
	{8'd123,8'd233} : s = 90;
	{8'd123,8'd234} : s = 217;
	{8'd123,8'd235} : s = 214;
	{8'd123,8'd236} : s = 373;
	{8'd123,8'd237} : s = 89;
	{8'd123,8'd238} : s = 213;
	{8'd123,8'd239} : s = 211;
	{8'd123,8'd240} : s = 371;
	{8'd123,8'd241} : s = 206;
	{8'd123,8'd242} : s = 366;
	{8'd123,8'd243} : s = 365;
	{8'd123,8'd244} : s = 478;
	{8'd123,8'd245} : s = 86;
	{8'd123,8'd246} : s = 205;
	{8'd123,8'd247} : s = 203;
	{8'd123,8'd248} : s = 363;
	{8'd123,8'd249} : s = 199;
	{8'd123,8'd250} : s = 359;
	{8'd123,8'd251} : s = 350;
	{8'd123,8'd252} : s = 477;
	{8'd123,8'd253} : s = 188;
	{8'd123,8'd254} : s = 349;
	{8'd123,8'd255} : s = 347;
	{8'd124,8'd0} : s = 426;
	{8'd124,8'd1} : s = 490;
	{8'd124,8'd2} : s = 489;
	{8'd124,8'd3} : s = 508;
	{8'd124,8'd4} : s = 2;
	{8'd124,8'd5} : s = 48;
	{8'd124,8'd6} : s = 40;
	{8'd124,8'd7} : s = 168;
	{8'd124,8'd8} : s = 36;
	{8'd124,8'd9} : s = 164;
	{8'd124,8'd10} : s = 162;
	{8'd124,8'd11} : s = 323;
	{8'd124,8'd12} : s = 34;
	{8'd124,8'd13} : s = 161;
	{8'd124,8'd14} : s = 152;
	{8'd124,8'd15} : s = 312;
	{8'd124,8'd16} : s = 148;
	{8'd124,8'd17} : s = 308;
	{8'd124,8'd18} : s = 306;
	{8'd124,8'd19} : s = 425;
	{8'd124,8'd20} : s = 33;
	{8'd124,8'd21} : s = 146;
	{8'd124,8'd22} : s = 145;
	{8'd124,8'd23} : s = 305;
	{8'd124,8'd24} : s = 140;
	{8'd124,8'd25} : s = 300;
	{8'd124,8'd26} : s = 298;
	{8'd124,8'd27} : s = 422;
	{8'd124,8'd28} : s = 138;
	{8'd124,8'd29} : s = 297;
	{8'd124,8'd30} : s = 294;
	{8'd124,8'd31} : s = 421;
	{8'd124,8'd32} : s = 293;
	{8'd124,8'd33} : s = 419;
	{8'd124,8'd34} : s = 412;
	{8'd124,8'd35} : s = 486;
	{8'd124,8'd36} : s = 24;
	{8'd124,8'd37} : s = 137;
	{8'd124,8'd38} : s = 134;
	{8'd124,8'd39} : s = 291;
	{8'd124,8'd40} : s = 133;
	{8'd124,8'd41} : s = 284;
	{8'd124,8'd42} : s = 282;
	{8'd124,8'd43} : s = 410;
	{8'd124,8'd44} : s = 131;
	{8'd124,8'd45} : s = 281;
	{8'd124,8'd46} : s = 278;
	{8'd124,8'd47} : s = 409;
	{8'd124,8'd48} : s = 277;
	{8'd124,8'd49} : s = 406;
	{8'd124,8'd50} : s = 405;
	{8'd124,8'd51} : s = 485;
	{8'd124,8'd52} : s = 112;
	{8'd124,8'd53} : s = 275;
	{8'd124,8'd54} : s = 270;
	{8'd124,8'd55} : s = 403;
	{8'd124,8'd56} : s = 269;
	{8'd124,8'd57} : s = 398;
	{8'd124,8'd58} : s = 397;
	{8'd124,8'd59} : s = 483;
	{8'd124,8'd60} : s = 267;
	{8'd124,8'd61} : s = 395;
	{8'd124,8'd62} : s = 391;
	{8'd124,8'd63} : s = 476;
	{8'd124,8'd64} : s = 376;
	{8'd124,8'd65} : s = 474;
	{8'd124,8'd66} : s = 473;
	{8'd124,8'd67} : s = 506;
	{8'd124,8'd68} : s = 20;
	{8'd124,8'd69} : s = 104;
	{8'd124,8'd70} : s = 100;
	{8'd124,8'd71} : s = 263;
	{8'd124,8'd72} : s = 98;
	{8'd124,8'd73} : s = 240;
	{8'd124,8'd74} : s = 232;
	{8'd124,8'd75} : s = 372;
	{8'd124,8'd76} : s = 97;
	{8'd124,8'd77} : s = 228;
	{8'd124,8'd78} : s = 226;
	{8'd124,8'd79} : s = 370;
	{8'd124,8'd80} : s = 225;
	{8'd124,8'd81} : s = 369;
	{8'd124,8'd82} : s = 364;
	{8'd124,8'd83} : s = 470;
	{8'd124,8'd84} : s = 88;
	{8'd124,8'd85} : s = 216;
	{8'd124,8'd86} : s = 212;
	{8'd124,8'd87} : s = 362;
	{8'd124,8'd88} : s = 210;
	{8'd124,8'd89} : s = 361;
	{8'd124,8'd90} : s = 358;
	{8'd124,8'd91} : s = 469;
	{8'd124,8'd92} : s = 209;
	{8'd124,8'd93} : s = 357;
	{8'd124,8'd94} : s = 355;
	{8'd124,8'd95} : s = 467;
	{8'd124,8'd96} : s = 348;
	{8'd124,8'd97} : s = 462;
	{8'd124,8'd98} : s = 461;
	{8'd124,8'd99} : s = 505;
	{8'd124,8'd100} : s = 84;
	{8'd124,8'd101} : s = 204;
	{8'd124,8'd102} : s = 202;
	{8'd124,8'd103} : s = 346;
	{8'd124,8'd104} : s = 201;
	{8'd124,8'd105} : s = 345;
	{8'd124,8'd106} : s = 342;
	{8'd124,8'd107} : s = 459;
	{8'd124,8'd108} : s = 198;
	{8'd124,8'd109} : s = 341;
	{8'd124,8'd110} : s = 339;
	{8'd124,8'd111} : s = 455;
	{8'd124,8'd112} : s = 334;
	{8'd124,8'd113} : s = 444;
	{8'd124,8'd114} : s = 442;
	{8'd124,8'd115} : s = 502;
	{8'd124,8'd116} : s = 197;
	{8'd124,8'd117} : s = 333;
	{8'd124,8'd118} : s = 331;
	{8'd124,8'd119} : s = 441;
	{8'd124,8'd120} : s = 327;
	{8'd124,8'd121} : s = 438;
	{8'd124,8'd122} : s = 437;
	{8'd124,8'd123} : s = 501;
	{8'd124,8'd124} : s = 316;
	{8'd124,8'd125} : s = 435;
	{8'd124,8'd126} : s = 430;
	{8'd124,8'd127} : s = 499;
	{8'd124,8'd128} : s = 429;
	{8'd124,8'd129} : s = 494;
	{8'd124,8'd130} : s = 493;
	{8'd124,8'd131} : s = 510;
	{8'd124,8'd132} : s = 1;
	{8'd124,8'd133} : s = 18;
	{8'd124,8'd134} : s = 17;
	{8'd124,8'd135} : s = 82;
	{8'd124,8'd136} : s = 12;
	{8'd124,8'd137} : s = 81;
	{8'd124,8'd138} : s = 76;
	{8'd124,8'd139} : s = 195;
	{8'd124,8'd140} : s = 10;
	{8'd124,8'd141} : s = 74;
	{8'd124,8'd142} : s = 73;
	{8'd124,8'd143} : s = 184;
	{8'd124,8'd144} : s = 70;
	{8'd124,8'd145} : s = 180;
	{8'd124,8'd146} : s = 178;
	{8'd124,8'd147} : s = 314;
	{8'd124,8'd148} : s = 9;
	{8'd124,8'd149} : s = 69;
	{8'd124,8'd150} : s = 67;
	{8'd124,8'd151} : s = 177;
	{8'd124,8'd152} : s = 56;
	{8'd124,8'd153} : s = 172;
	{8'd124,8'd154} : s = 170;
	{8'd124,8'd155} : s = 313;
	{8'd124,8'd156} : s = 52;
	{8'd124,8'd157} : s = 169;
	{8'd124,8'd158} : s = 166;
	{8'd124,8'd159} : s = 310;
	{8'd124,8'd160} : s = 165;
	{8'd124,8'd161} : s = 309;
	{8'd124,8'd162} : s = 307;
	{8'd124,8'd163} : s = 427;
	{8'd124,8'd164} : s = 6;
	{8'd124,8'd165} : s = 50;
	{8'd124,8'd166} : s = 49;
	{8'd124,8'd167} : s = 163;
	{8'd124,8'd168} : s = 44;
	{8'd124,8'd169} : s = 156;
	{8'd124,8'd170} : s = 154;
	{8'd124,8'd171} : s = 302;
	{8'd124,8'd172} : s = 42;
	{8'd124,8'd173} : s = 153;
	{8'd124,8'd174} : s = 150;
	{8'd124,8'd175} : s = 301;
	{8'd124,8'd176} : s = 149;
	{8'd124,8'd177} : s = 299;
	{8'd124,8'd178} : s = 295;
	{8'd124,8'd179} : s = 423;
	{8'd124,8'd180} : s = 41;
	{8'd124,8'd181} : s = 147;
	{8'd124,8'd182} : s = 142;
	{8'd124,8'd183} : s = 286;
	{8'd124,8'd184} : s = 141;
	{8'd124,8'd185} : s = 285;
	{8'd124,8'd186} : s = 283;
	{8'd124,8'd187} : s = 414;
	{8'd124,8'd188} : s = 139;
	{8'd124,8'd189} : s = 279;
	{8'd124,8'd190} : s = 271;
	{8'd124,8'd191} : s = 413;
	{8'd124,8'd192} : s = 248;
	{8'd124,8'd193} : s = 411;
	{8'd124,8'd194} : s = 407;
	{8'd124,8'd195} : s = 491;
	{8'd124,8'd196} : s = 5;
	{8'd124,8'd197} : s = 38;
	{8'd124,8'd198} : s = 37;
	{8'd124,8'd199} : s = 135;
	{8'd124,8'd200} : s = 35;
	{8'd124,8'd201} : s = 120;
	{8'd124,8'd202} : s = 116;
	{8'd124,8'd203} : s = 244;
	{8'd124,8'd204} : s = 28;
	{8'd124,8'd205} : s = 114;
	{8'd124,8'd206} : s = 113;
	{8'd124,8'd207} : s = 242;
	{8'd124,8'd208} : s = 108;
	{8'd124,8'd209} : s = 241;
	{8'd124,8'd210} : s = 236;
	{8'd124,8'd211} : s = 399;
	{8'd124,8'd212} : s = 26;
	{8'd124,8'd213} : s = 106;
	{8'd124,8'd214} : s = 105;
	{8'd124,8'd215} : s = 234;
	{8'd124,8'd216} : s = 102;
	{8'd124,8'd217} : s = 233;
	{8'd124,8'd218} : s = 230;
	{8'd124,8'd219} : s = 380;
	{8'd124,8'd220} : s = 101;
	{8'd124,8'd221} : s = 229;
	{8'd124,8'd222} : s = 227;
	{8'd124,8'd223} : s = 378;
	{8'd124,8'd224} : s = 220;
	{8'd124,8'd225} : s = 377;
	{8'd124,8'd226} : s = 374;
	{8'd124,8'd227} : s = 487;
	{8'd124,8'd228} : s = 25;
	{8'd124,8'd229} : s = 99;
	{8'd124,8'd230} : s = 92;
	{8'd124,8'd231} : s = 218;
	{8'd124,8'd232} : s = 90;
	{8'd124,8'd233} : s = 217;
	{8'd124,8'd234} : s = 214;
	{8'd124,8'd235} : s = 373;
	{8'd124,8'd236} : s = 89;
	{8'd124,8'd237} : s = 213;
	{8'd124,8'd238} : s = 211;
	{8'd124,8'd239} : s = 371;
	{8'd124,8'd240} : s = 206;
	{8'd124,8'd241} : s = 366;
	{8'd124,8'd242} : s = 365;
	{8'd124,8'd243} : s = 478;
	{8'd124,8'd244} : s = 86;
	{8'd124,8'd245} : s = 205;
	{8'd124,8'd246} : s = 203;
	{8'd124,8'd247} : s = 363;
	{8'd124,8'd248} : s = 199;
	{8'd124,8'd249} : s = 359;
	{8'd124,8'd250} : s = 350;
	{8'd124,8'd251} : s = 477;
	{8'd124,8'd252} : s = 188;
	{8'd124,8'd253} : s = 349;
	{8'd124,8'd254} : s = 347;
	{8'd124,8'd255} : s = 475;
	{8'd125,8'd0} : s = 490;
	{8'd125,8'd1} : s = 489;
	{8'd125,8'd2} : s = 508;
	{8'd125,8'd3} : s = 2;
	{8'd125,8'd4} : s = 48;
	{8'd125,8'd5} : s = 40;
	{8'd125,8'd6} : s = 168;
	{8'd125,8'd7} : s = 36;
	{8'd125,8'd8} : s = 164;
	{8'd125,8'd9} : s = 162;
	{8'd125,8'd10} : s = 323;
	{8'd125,8'd11} : s = 34;
	{8'd125,8'd12} : s = 161;
	{8'd125,8'd13} : s = 152;
	{8'd125,8'd14} : s = 312;
	{8'd125,8'd15} : s = 148;
	{8'd125,8'd16} : s = 308;
	{8'd125,8'd17} : s = 306;
	{8'd125,8'd18} : s = 425;
	{8'd125,8'd19} : s = 33;
	{8'd125,8'd20} : s = 146;
	{8'd125,8'd21} : s = 145;
	{8'd125,8'd22} : s = 305;
	{8'd125,8'd23} : s = 140;
	{8'd125,8'd24} : s = 300;
	{8'd125,8'd25} : s = 298;
	{8'd125,8'd26} : s = 422;
	{8'd125,8'd27} : s = 138;
	{8'd125,8'd28} : s = 297;
	{8'd125,8'd29} : s = 294;
	{8'd125,8'd30} : s = 421;
	{8'd125,8'd31} : s = 293;
	{8'd125,8'd32} : s = 419;
	{8'd125,8'd33} : s = 412;
	{8'd125,8'd34} : s = 486;
	{8'd125,8'd35} : s = 24;
	{8'd125,8'd36} : s = 137;
	{8'd125,8'd37} : s = 134;
	{8'd125,8'd38} : s = 291;
	{8'd125,8'd39} : s = 133;
	{8'd125,8'd40} : s = 284;
	{8'd125,8'd41} : s = 282;
	{8'd125,8'd42} : s = 410;
	{8'd125,8'd43} : s = 131;
	{8'd125,8'd44} : s = 281;
	{8'd125,8'd45} : s = 278;
	{8'd125,8'd46} : s = 409;
	{8'd125,8'd47} : s = 277;
	{8'd125,8'd48} : s = 406;
	{8'd125,8'd49} : s = 405;
	{8'd125,8'd50} : s = 485;
	{8'd125,8'd51} : s = 112;
	{8'd125,8'd52} : s = 275;
	{8'd125,8'd53} : s = 270;
	{8'd125,8'd54} : s = 403;
	{8'd125,8'd55} : s = 269;
	{8'd125,8'd56} : s = 398;
	{8'd125,8'd57} : s = 397;
	{8'd125,8'd58} : s = 483;
	{8'd125,8'd59} : s = 267;
	{8'd125,8'd60} : s = 395;
	{8'd125,8'd61} : s = 391;
	{8'd125,8'd62} : s = 476;
	{8'd125,8'd63} : s = 376;
	{8'd125,8'd64} : s = 474;
	{8'd125,8'd65} : s = 473;
	{8'd125,8'd66} : s = 506;
	{8'd125,8'd67} : s = 20;
	{8'd125,8'd68} : s = 104;
	{8'd125,8'd69} : s = 100;
	{8'd125,8'd70} : s = 263;
	{8'd125,8'd71} : s = 98;
	{8'd125,8'd72} : s = 240;
	{8'd125,8'd73} : s = 232;
	{8'd125,8'd74} : s = 372;
	{8'd125,8'd75} : s = 97;
	{8'd125,8'd76} : s = 228;
	{8'd125,8'd77} : s = 226;
	{8'd125,8'd78} : s = 370;
	{8'd125,8'd79} : s = 225;
	{8'd125,8'd80} : s = 369;
	{8'd125,8'd81} : s = 364;
	{8'd125,8'd82} : s = 470;
	{8'd125,8'd83} : s = 88;
	{8'd125,8'd84} : s = 216;
	{8'd125,8'd85} : s = 212;
	{8'd125,8'd86} : s = 362;
	{8'd125,8'd87} : s = 210;
	{8'd125,8'd88} : s = 361;
	{8'd125,8'd89} : s = 358;
	{8'd125,8'd90} : s = 469;
	{8'd125,8'd91} : s = 209;
	{8'd125,8'd92} : s = 357;
	{8'd125,8'd93} : s = 355;
	{8'd125,8'd94} : s = 467;
	{8'd125,8'd95} : s = 348;
	{8'd125,8'd96} : s = 462;
	{8'd125,8'd97} : s = 461;
	{8'd125,8'd98} : s = 505;
	{8'd125,8'd99} : s = 84;
	{8'd125,8'd100} : s = 204;
	{8'd125,8'd101} : s = 202;
	{8'd125,8'd102} : s = 346;
	{8'd125,8'd103} : s = 201;
	{8'd125,8'd104} : s = 345;
	{8'd125,8'd105} : s = 342;
	{8'd125,8'd106} : s = 459;
	{8'd125,8'd107} : s = 198;
	{8'd125,8'd108} : s = 341;
	{8'd125,8'd109} : s = 339;
	{8'd125,8'd110} : s = 455;
	{8'd125,8'd111} : s = 334;
	{8'd125,8'd112} : s = 444;
	{8'd125,8'd113} : s = 442;
	{8'd125,8'd114} : s = 502;
	{8'd125,8'd115} : s = 197;
	{8'd125,8'd116} : s = 333;
	{8'd125,8'd117} : s = 331;
	{8'd125,8'd118} : s = 441;
	{8'd125,8'd119} : s = 327;
	{8'd125,8'd120} : s = 438;
	{8'd125,8'd121} : s = 437;
	{8'd125,8'd122} : s = 501;
	{8'd125,8'd123} : s = 316;
	{8'd125,8'd124} : s = 435;
	{8'd125,8'd125} : s = 430;
	{8'd125,8'd126} : s = 499;
	{8'd125,8'd127} : s = 429;
	{8'd125,8'd128} : s = 494;
	{8'd125,8'd129} : s = 493;
	{8'd125,8'd130} : s = 510;
	{8'd125,8'd131} : s = 1;
	{8'd125,8'd132} : s = 18;
	{8'd125,8'd133} : s = 17;
	{8'd125,8'd134} : s = 82;
	{8'd125,8'd135} : s = 12;
	{8'd125,8'd136} : s = 81;
	{8'd125,8'd137} : s = 76;
	{8'd125,8'd138} : s = 195;
	{8'd125,8'd139} : s = 10;
	{8'd125,8'd140} : s = 74;
	{8'd125,8'd141} : s = 73;
	{8'd125,8'd142} : s = 184;
	{8'd125,8'd143} : s = 70;
	{8'd125,8'd144} : s = 180;
	{8'd125,8'd145} : s = 178;
	{8'd125,8'd146} : s = 314;
	{8'd125,8'd147} : s = 9;
	{8'd125,8'd148} : s = 69;
	{8'd125,8'd149} : s = 67;
	{8'd125,8'd150} : s = 177;
	{8'd125,8'd151} : s = 56;
	{8'd125,8'd152} : s = 172;
	{8'd125,8'd153} : s = 170;
	{8'd125,8'd154} : s = 313;
	{8'd125,8'd155} : s = 52;
	{8'd125,8'd156} : s = 169;
	{8'd125,8'd157} : s = 166;
	{8'd125,8'd158} : s = 310;
	{8'd125,8'd159} : s = 165;
	{8'd125,8'd160} : s = 309;
	{8'd125,8'd161} : s = 307;
	{8'd125,8'd162} : s = 427;
	{8'd125,8'd163} : s = 6;
	{8'd125,8'd164} : s = 50;
	{8'd125,8'd165} : s = 49;
	{8'd125,8'd166} : s = 163;
	{8'd125,8'd167} : s = 44;
	{8'd125,8'd168} : s = 156;
	{8'd125,8'd169} : s = 154;
	{8'd125,8'd170} : s = 302;
	{8'd125,8'd171} : s = 42;
	{8'd125,8'd172} : s = 153;
	{8'd125,8'd173} : s = 150;
	{8'd125,8'd174} : s = 301;
	{8'd125,8'd175} : s = 149;
	{8'd125,8'd176} : s = 299;
	{8'd125,8'd177} : s = 295;
	{8'd125,8'd178} : s = 423;
	{8'd125,8'd179} : s = 41;
	{8'd125,8'd180} : s = 147;
	{8'd125,8'd181} : s = 142;
	{8'd125,8'd182} : s = 286;
	{8'd125,8'd183} : s = 141;
	{8'd125,8'd184} : s = 285;
	{8'd125,8'd185} : s = 283;
	{8'd125,8'd186} : s = 414;
	{8'd125,8'd187} : s = 139;
	{8'd125,8'd188} : s = 279;
	{8'd125,8'd189} : s = 271;
	{8'd125,8'd190} : s = 413;
	{8'd125,8'd191} : s = 248;
	{8'd125,8'd192} : s = 411;
	{8'd125,8'd193} : s = 407;
	{8'd125,8'd194} : s = 491;
	{8'd125,8'd195} : s = 5;
	{8'd125,8'd196} : s = 38;
	{8'd125,8'd197} : s = 37;
	{8'd125,8'd198} : s = 135;
	{8'd125,8'd199} : s = 35;
	{8'd125,8'd200} : s = 120;
	{8'd125,8'd201} : s = 116;
	{8'd125,8'd202} : s = 244;
	{8'd125,8'd203} : s = 28;
	{8'd125,8'd204} : s = 114;
	{8'd125,8'd205} : s = 113;
	{8'd125,8'd206} : s = 242;
	{8'd125,8'd207} : s = 108;
	{8'd125,8'd208} : s = 241;
	{8'd125,8'd209} : s = 236;
	{8'd125,8'd210} : s = 399;
	{8'd125,8'd211} : s = 26;
	{8'd125,8'd212} : s = 106;
	{8'd125,8'd213} : s = 105;
	{8'd125,8'd214} : s = 234;
	{8'd125,8'd215} : s = 102;
	{8'd125,8'd216} : s = 233;
	{8'd125,8'd217} : s = 230;
	{8'd125,8'd218} : s = 380;
	{8'd125,8'd219} : s = 101;
	{8'd125,8'd220} : s = 229;
	{8'd125,8'd221} : s = 227;
	{8'd125,8'd222} : s = 378;
	{8'd125,8'd223} : s = 220;
	{8'd125,8'd224} : s = 377;
	{8'd125,8'd225} : s = 374;
	{8'd125,8'd226} : s = 487;
	{8'd125,8'd227} : s = 25;
	{8'd125,8'd228} : s = 99;
	{8'd125,8'd229} : s = 92;
	{8'd125,8'd230} : s = 218;
	{8'd125,8'd231} : s = 90;
	{8'd125,8'd232} : s = 217;
	{8'd125,8'd233} : s = 214;
	{8'd125,8'd234} : s = 373;
	{8'd125,8'd235} : s = 89;
	{8'd125,8'd236} : s = 213;
	{8'd125,8'd237} : s = 211;
	{8'd125,8'd238} : s = 371;
	{8'd125,8'd239} : s = 206;
	{8'd125,8'd240} : s = 366;
	{8'd125,8'd241} : s = 365;
	{8'd125,8'd242} : s = 478;
	{8'd125,8'd243} : s = 86;
	{8'd125,8'd244} : s = 205;
	{8'd125,8'd245} : s = 203;
	{8'd125,8'd246} : s = 363;
	{8'd125,8'd247} : s = 199;
	{8'd125,8'd248} : s = 359;
	{8'd125,8'd249} : s = 350;
	{8'd125,8'd250} : s = 477;
	{8'd125,8'd251} : s = 188;
	{8'd125,8'd252} : s = 349;
	{8'd125,8'd253} : s = 347;
	{8'd125,8'd254} : s = 475;
	{8'd125,8'd255} : s = 343;
	{8'd126,8'd0} : s = 489;
	{8'd126,8'd1} : s = 508;
	{8'd126,8'd2} : s = 2;
	{8'd126,8'd3} : s = 48;
	{8'd126,8'd4} : s = 40;
	{8'd126,8'd5} : s = 168;
	{8'd126,8'd6} : s = 36;
	{8'd126,8'd7} : s = 164;
	{8'd126,8'd8} : s = 162;
	{8'd126,8'd9} : s = 323;
	{8'd126,8'd10} : s = 34;
	{8'd126,8'd11} : s = 161;
	{8'd126,8'd12} : s = 152;
	{8'd126,8'd13} : s = 312;
	{8'd126,8'd14} : s = 148;
	{8'd126,8'd15} : s = 308;
	{8'd126,8'd16} : s = 306;
	{8'd126,8'd17} : s = 425;
	{8'd126,8'd18} : s = 33;
	{8'd126,8'd19} : s = 146;
	{8'd126,8'd20} : s = 145;
	{8'd126,8'd21} : s = 305;
	{8'd126,8'd22} : s = 140;
	{8'd126,8'd23} : s = 300;
	{8'd126,8'd24} : s = 298;
	{8'd126,8'd25} : s = 422;
	{8'd126,8'd26} : s = 138;
	{8'd126,8'd27} : s = 297;
	{8'd126,8'd28} : s = 294;
	{8'd126,8'd29} : s = 421;
	{8'd126,8'd30} : s = 293;
	{8'd126,8'd31} : s = 419;
	{8'd126,8'd32} : s = 412;
	{8'd126,8'd33} : s = 486;
	{8'd126,8'd34} : s = 24;
	{8'd126,8'd35} : s = 137;
	{8'd126,8'd36} : s = 134;
	{8'd126,8'd37} : s = 291;
	{8'd126,8'd38} : s = 133;
	{8'd126,8'd39} : s = 284;
	{8'd126,8'd40} : s = 282;
	{8'd126,8'd41} : s = 410;
	{8'd126,8'd42} : s = 131;
	{8'd126,8'd43} : s = 281;
	{8'd126,8'd44} : s = 278;
	{8'd126,8'd45} : s = 409;
	{8'd126,8'd46} : s = 277;
	{8'd126,8'd47} : s = 406;
	{8'd126,8'd48} : s = 405;
	{8'd126,8'd49} : s = 485;
	{8'd126,8'd50} : s = 112;
	{8'd126,8'd51} : s = 275;
	{8'd126,8'd52} : s = 270;
	{8'd126,8'd53} : s = 403;
	{8'd126,8'd54} : s = 269;
	{8'd126,8'd55} : s = 398;
	{8'd126,8'd56} : s = 397;
	{8'd126,8'd57} : s = 483;
	{8'd126,8'd58} : s = 267;
	{8'd126,8'd59} : s = 395;
	{8'd126,8'd60} : s = 391;
	{8'd126,8'd61} : s = 476;
	{8'd126,8'd62} : s = 376;
	{8'd126,8'd63} : s = 474;
	{8'd126,8'd64} : s = 473;
	{8'd126,8'd65} : s = 506;
	{8'd126,8'd66} : s = 20;
	{8'd126,8'd67} : s = 104;
	{8'd126,8'd68} : s = 100;
	{8'd126,8'd69} : s = 263;
	{8'd126,8'd70} : s = 98;
	{8'd126,8'd71} : s = 240;
	{8'd126,8'd72} : s = 232;
	{8'd126,8'd73} : s = 372;
	{8'd126,8'd74} : s = 97;
	{8'd126,8'd75} : s = 228;
	{8'd126,8'd76} : s = 226;
	{8'd126,8'd77} : s = 370;
	{8'd126,8'd78} : s = 225;
	{8'd126,8'd79} : s = 369;
	{8'd126,8'd80} : s = 364;
	{8'd126,8'd81} : s = 470;
	{8'd126,8'd82} : s = 88;
	{8'd126,8'd83} : s = 216;
	{8'd126,8'd84} : s = 212;
	{8'd126,8'd85} : s = 362;
	{8'd126,8'd86} : s = 210;
	{8'd126,8'd87} : s = 361;
	{8'd126,8'd88} : s = 358;
	{8'd126,8'd89} : s = 469;
	{8'd126,8'd90} : s = 209;
	{8'd126,8'd91} : s = 357;
	{8'd126,8'd92} : s = 355;
	{8'd126,8'd93} : s = 467;
	{8'd126,8'd94} : s = 348;
	{8'd126,8'd95} : s = 462;
	{8'd126,8'd96} : s = 461;
	{8'd126,8'd97} : s = 505;
	{8'd126,8'd98} : s = 84;
	{8'd126,8'd99} : s = 204;
	{8'd126,8'd100} : s = 202;
	{8'd126,8'd101} : s = 346;
	{8'd126,8'd102} : s = 201;
	{8'd126,8'd103} : s = 345;
	{8'd126,8'd104} : s = 342;
	{8'd126,8'd105} : s = 459;
	{8'd126,8'd106} : s = 198;
	{8'd126,8'd107} : s = 341;
	{8'd126,8'd108} : s = 339;
	{8'd126,8'd109} : s = 455;
	{8'd126,8'd110} : s = 334;
	{8'd126,8'd111} : s = 444;
	{8'd126,8'd112} : s = 442;
	{8'd126,8'd113} : s = 502;
	{8'd126,8'd114} : s = 197;
	{8'd126,8'd115} : s = 333;
	{8'd126,8'd116} : s = 331;
	{8'd126,8'd117} : s = 441;
	{8'd126,8'd118} : s = 327;
	{8'd126,8'd119} : s = 438;
	{8'd126,8'd120} : s = 437;
	{8'd126,8'd121} : s = 501;
	{8'd126,8'd122} : s = 316;
	{8'd126,8'd123} : s = 435;
	{8'd126,8'd124} : s = 430;
	{8'd126,8'd125} : s = 499;
	{8'd126,8'd126} : s = 429;
	{8'd126,8'd127} : s = 494;
	{8'd126,8'd128} : s = 493;
	{8'd126,8'd129} : s = 510;
	{8'd126,8'd130} : s = 1;
	{8'd126,8'd131} : s = 18;
	{8'd126,8'd132} : s = 17;
	{8'd126,8'd133} : s = 82;
	{8'd126,8'd134} : s = 12;
	{8'd126,8'd135} : s = 81;
	{8'd126,8'd136} : s = 76;
	{8'd126,8'd137} : s = 195;
	{8'd126,8'd138} : s = 10;
	{8'd126,8'd139} : s = 74;
	{8'd126,8'd140} : s = 73;
	{8'd126,8'd141} : s = 184;
	{8'd126,8'd142} : s = 70;
	{8'd126,8'd143} : s = 180;
	{8'd126,8'd144} : s = 178;
	{8'd126,8'd145} : s = 314;
	{8'd126,8'd146} : s = 9;
	{8'd126,8'd147} : s = 69;
	{8'd126,8'd148} : s = 67;
	{8'd126,8'd149} : s = 177;
	{8'd126,8'd150} : s = 56;
	{8'd126,8'd151} : s = 172;
	{8'd126,8'd152} : s = 170;
	{8'd126,8'd153} : s = 313;
	{8'd126,8'd154} : s = 52;
	{8'd126,8'd155} : s = 169;
	{8'd126,8'd156} : s = 166;
	{8'd126,8'd157} : s = 310;
	{8'd126,8'd158} : s = 165;
	{8'd126,8'd159} : s = 309;
	{8'd126,8'd160} : s = 307;
	{8'd126,8'd161} : s = 427;
	{8'd126,8'd162} : s = 6;
	{8'd126,8'd163} : s = 50;
	{8'd126,8'd164} : s = 49;
	{8'd126,8'd165} : s = 163;
	{8'd126,8'd166} : s = 44;
	{8'd126,8'd167} : s = 156;
	{8'd126,8'd168} : s = 154;
	{8'd126,8'd169} : s = 302;
	{8'd126,8'd170} : s = 42;
	{8'd126,8'd171} : s = 153;
	{8'd126,8'd172} : s = 150;
	{8'd126,8'd173} : s = 301;
	{8'd126,8'd174} : s = 149;
	{8'd126,8'd175} : s = 299;
	{8'd126,8'd176} : s = 295;
	{8'd126,8'd177} : s = 423;
	{8'd126,8'd178} : s = 41;
	{8'd126,8'd179} : s = 147;
	{8'd126,8'd180} : s = 142;
	{8'd126,8'd181} : s = 286;
	{8'd126,8'd182} : s = 141;
	{8'd126,8'd183} : s = 285;
	{8'd126,8'd184} : s = 283;
	{8'd126,8'd185} : s = 414;
	{8'd126,8'd186} : s = 139;
	{8'd126,8'd187} : s = 279;
	{8'd126,8'd188} : s = 271;
	{8'd126,8'd189} : s = 413;
	{8'd126,8'd190} : s = 248;
	{8'd126,8'd191} : s = 411;
	{8'd126,8'd192} : s = 407;
	{8'd126,8'd193} : s = 491;
	{8'd126,8'd194} : s = 5;
	{8'd126,8'd195} : s = 38;
	{8'd126,8'd196} : s = 37;
	{8'd126,8'd197} : s = 135;
	{8'd126,8'd198} : s = 35;
	{8'd126,8'd199} : s = 120;
	{8'd126,8'd200} : s = 116;
	{8'd126,8'd201} : s = 244;
	{8'd126,8'd202} : s = 28;
	{8'd126,8'd203} : s = 114;
	{8'd126,8'd204} : s = 113;
	{8'd126,8'd205} : s = 242;
	{8'd126,8'd206} : s = 108;
	{8'd126,8'd207} : s = 241;
	{8'd126,8'd208} : s = 236;
	{8'd126,8'd209} : s = 399;
	{8'd126,8'd210} : s = 26;
	{8'd126,8'd211} : s = 106;
	{8'd126,8'd212} : s = 105;
	{8'd126,8'd213} : s = 234;
	{8'd126,8'd214} : s = 102;
	{8'd126,8'd215} : s = 233;
	{8'd126,8'd216} : s = 230;
	{8'd126,8'd217} : s = 380;
	{8'd126,8'd218} : s = 101;
	{8'd126,8'd219} : s = 229;
	{8'd126,8'd220} : s = 227;
	{8'd126,8'd221} : s = 378;
	{8'd126,8'd222} : s = 220;
	{8'd126,8'd223} : s = 377;
	{8'd126,8'd224} : s = 374;
	{8'd126,8'd225} : s = 487;
	{8'd126,8'd226} : s = 25;
	{8'd126,8'd227} : s = 99;
	{8'd126,8'd228} : s = 92;
	{8'd126,8'd229} : s = 218;
	{8'd126,8'd230} : s = 90;
	{8'd126,8'd231} : s = 217;
	{8'd126,8'd232} : s = 214;
	{8'd126,8'd233} : s = 373;
	{8'd126,8'd234} : s = 89;
	{8'd126,8'd235} : s = 213;
	{8'd126,8'd236} : s = 211;
	{8'd126,8'd237} : s = 371;
	{8'd126,8'd238} : s = 206;
	{8'd126,8'd239} : s = 366;
	{8'd126,8'd240} : s = 365;
	{8'd126,8'd241} : s = 478;
	{8'd126,8'd242} : s = 86;
	{8'd126,8'd243} : s = 205;
	{8'd126,8'd244} : s = 203;
	{8'd126,8'd245} : s = 363;
	{8'd126,8'd246} : s = 199;
	{8'd126,8'd247} : s = 359;
	{8'd126,8'd248} : s = 350;
	{8'd126,8'd249} : s = 477;
	{8'd126,8'd250} : s = 188;
	{8'd126,8'd251} : s = 349;
	{8'd126,8'd252} : s = 347;
	{8'd126,8'd253} : s = 475;
	{8'd126,8'd254} : s = 343;
	{8'd126,8'd255} : s = 471;
	{8'd127,8'd0} : s = 508;
	{8'd127,8'd1} : s = 2;
	{8'd127,8'd2} : s = 48;
	{8'd127,8'd3} : s = 40;
	{8'd127,8'd4} : s = 168;
	{8'd127,8'd5} : s = 36;
	{8'd127,8'd6} : s = 164;
	{8'd127,8'd7} : s = 162;
	{8'd127,8'd8} : s = 323;
	{8'd127,8'd9} : s = 34;
	{8'd127,8'd10} : s = 161;
	{8'd127,8'd11} : s = 152;
	{8'd127,8'd12} : s = 312;
	{8'd127,8'd13} : s = 148;
	{8'd127,8'd14} : s = 308;
	{8'd127,8'd15} : s = 306;
	{8'd127,8'd16} : s = 425;
	{8'd127,8'd17} : s = 33;
	{8'd127,8'd18} : s = 146;
	{8'd127,8'd19} : s = 145;
	{8'd127,8'd20} : s = 305;
	{8'd127,8'd21} : s = 140;
	{8'd127,8'd22} : s = 300;
	{8'd127,8'd23} : s = 298;
	{8'd127,8'd24} : s = 422;
	{8'd127,8'd25} : s = 138;
	{8'd127,8'd26} : s = 297;
	{8'd127,8'd27} : s = 294;
	{8'd127,8'd28} : s = 421;
	{8'd127,8'd29} : s = 293;
	{8'd127,8'd30} : s = 419;
	{8'd127,8'd31} : s = 412;
	{8'd127,8'd32} : s = 486;
	{8'd127,8'd33} : s = 24;
	{8'd127,8'd34} : s = 137;
	{8'd127,8'd35} : s = 134;
	{8'd127,8'd36} : s = 291;
	{8'd127,8'd37} : s = 133;
	{8'd127,8'd38} : s = 284;
	{8'd127,8'd39} : s = 282;
	{8'd127,8'd40} : s = 410;
	{8'd127,8'd41} : s = 131;
	{8'd127,8'd42} : s = 281;
	{8'd127,8'd43} : s = 278;
	{8'd127,8'd44} : s = 409;
	{8'd127,8'd45} : s = 277;
	{8'd127,8'd46} : s = 406;
	{8'd127,8'd47} : s = 405;
	{8'd127,8'd48} : s = 485;
	{8'd127,8'd49} : s = 112;
	{8'd127,8'd50} : s = 275;
	{8'd127,8'd51} : s = 270;
	{8'd127,8'd52} : s = 403;
	{8'd127,8'd53} : s = 269;
	{8'd127,8'd54} : s = 398;
	{8'd127,8'd55} : s = 397;
	{8'd127,8'd56} : s = 483;
	{8'd127,8'd57} : s = 267;
	{8'd127,8'd58} : s = 395;
	{8'd127,8'd59} : s = 391;
	{8'd127,8'd60} : s = 476;
	{8'd127,8'd61} : s = 376;
	{8'd127,8'd62} : s = 474;
	{8'd127,8'd63} : s = 473;
	{8'd127,8'd64} : s = 506;
	{8'd127,8'd65} : s = 20;
	{8'd127,8'd66} : s = 104;
	{8'd127,8'd67} : s = 100;
	{8'd127,8'd68} : s = 263;
	{8'd127,8'd69} : s = 98;
	{8'd127,8'd70} : s = 240;
	{8'd127,8'd71} : s = 232;
	{8'd127,8'd72} : s = 372;
	{8'd127,8'd73} : s = 97;
	{8'd127,8'd74} : s = 228;
	{8'd127,8'd75} : s = 226;
	{8'd127,8'd76} : s = 370;
	{8'd127,8'd77} : s = 225;
	{8'd127,8'd78} : s = 369;
	{8'd127,8'd79} : s = 364;
	{8'd127,8'd80} : s = 470;
	{8'd127,8'd81} : s = 88;
	{8'd127,8'd82} : s = 216;
	{8'd127,8'd83} : s = 212;
	{8'd127,8'd84} : s = 362;
	{8'd127,8'd85} : s = 210;
	{8'd127,8'd86} : s = 361;
	{8'd127,8'd87} : s = 358;
	{8'd127,8'd88} : s = 469;
	{8'd127,8'd89} : s = 209;
	{8'd127,8'd90} : s = 357;
	{8'd127,8'd91} : s = 355;
	{8'd127,8'd92} : s = 467;
	{8'd127,8'd93} : s = 348;
	{8'd127,8'd94} : s = 462;
	{8'd127,8'd95} : s = 461;
	{8'd127,8'd96} : s = 505;
	{8'd127,8'd97} : s = 84;
	{8'd127,8'd98} : s = 204;
	{8'd127,8'd99} : s = 202;
	{8'd127,8'd100} : s = 346;
	{8'd127,8'd101} : s = 201;
	{8'd127,8'd102} : s = 345;
	{8'd127,8'd103} : s = 342;
	{8'd127,8'd104} : s = 459;
	{8'd127,8'd105} : s = 198;
	{8'd127,8'd106} : s = 341;
	{8'd127,8'd107} : s = 339;
	{8'd127,8'd108} : s = 455;
	{8'd127,8'd109} : s = 334;
	{8'd127,8'd110} : s = 444;
	{8'd127,8'd111} : s = 442;
	{8'd127,8'd112} : s = 502;
	{8'd127,8'd113} : s = 197;
	{8'd127,8'd114} : s = 333;
	{8'd127,8'd115} : s = 331;
	{8'd127,8'd116} : s = 441;
	{8'd127,8'd117} : s = 327;
	{8'd127,8'd118} : s = 438;
	{8'd127,8'd119} : s = 437;
	{8'd127,8'd120} : s = 501;
	{8'd127,8'd121} : s = 316;
	{8'd127,8'd122} : s = 435;
	{8'd127,8'd123} : s = 430;
	{8'd127,8'd124} : s = 499;
	{8'd127,8'd125} : s = 429;
	{8'd127,8'd126} : s = 494;
	{8'd127,8'd127} : s = 493;
	{8'd127,8'd128} : s = 510;
	{8'd127,8'd129} : s = 1;
	{8'd127,8'd130} : s = 18;
	{8'd127,8'd131} : s = 17;
	{8'd127,8'd132} : s = 82;
	{8'd127,8'd133} : s = 12;
	{8'd127,8'd134} : s = 81;
	{8'd127,8'd135} : s = 76;
	{8'd127,8'd136} : s = 195;
	{8'd127,8'd137} : s = 10;
	{8'd127,8'd138} : s = 74;
	{8'd127,8'd139} : s = 73;
	{8'd127,8'd140} : s = 184;
	{8'd127,8'd141} : s = 70;
	{8'd127,8'd142} : s = 180;
	{8'd127,8'd143} : s = 178;
	{8'd127,8'd144} : s = 314;
	{8'd127,8'd145} : s = 9;
	{8'd127,8'd146} : s = 69;
	{8'd127,8'd147} : s = 67;
	{8'd127,8'd148} : s = 177;
	{8'd127,8'd149} : s = 56;
	{8'd127,8'd150} : s = 172;
	{8'd127,8'd151} : s = 170;
	{8'd127,8'd152} : s = 313;
	{8'd127,8'd153} : s = 52;
	{8'd127,8'd154} : s = 169;
	{8'd127,8'd155} : s = 166;
	{8'd127,8'd156} : s = 310;
	{8'd127,8'd157} : s = 165;
	{8'd127,8'd158} : s = 309;
	{8'd127,8'd159} : s = 307;
	{8'd127,8'd160} : s = 427;
	{8'd127,8'd161} : s = 6;
	{8'd127,8'd162} : s = 50;
	{8'd127,8'd163} : s = 49;
	{8'd127,8'd164} : s = 163;
	{8'd127,8'd165} : s = 44;
	{8'd127,8'd166} : s = 156;
	{8'd127,8'd167} : s = 154;
	{8'd127,8'd168} : s = 302;
	{8'd127,8'd169} : s = 42;
	{8'd127,8'd170} : s = 153;
	{8'd127,8'd171} : s = 150;
	{8'd127,8'd172} : s = 301;
	{8'd127,8'd173} : s = 149;
	{8'd127,8'd174} : s = 299;
	{8'd127,8'd175} : s = 295;
	{8'd127,8'd176} : s = 423;
	{8'd127,8'd177} : s = 41;
	{8'd127,8'd178} : s = 147;
	{8'd127,8'd179} : s = 142;
	{8'd127,8'd180} : s = 286;
	{8'd127,8'd181} : s = 141;
	{8'd127,8'd182} : s = 285;
	{8'd127,8'd183} : s = 283;
	{8'd127,8'd184} : s = 414;
	{8'd127,8'd185} : s = 139;
	{8'd127,8'd186} : s = 279;
	{8'd127,8'd187} : s = 271;
	{8'd127,8'd188} : s = 413;
	{8'd127,8'd189} : s = 248;
	{8'd127,8'd190} : s = 411;
	{8'd127,8'd191} : s = 407;
	{8'd127,8'd192} : s = 491;
	{8'd127,8'd193} : s = 5;
	{8'd127,8'd194} : s = 38;
	{8'd127,8'd195} : s = 37;
	{8'd127,8'd196} : s = 135;
	{8'd127,8'd197} : s = 35;
	{8'd127,8'd198} : s = 120;
	{8'd127,8'd199} : s = 116;
	{8'd127,8'd200} : s = 244;
	{8'd127,8'd201} : s = 28;
	{8'd127,8'd202} : s = 114;
	{8'd127,8'd203} : s = 113;
	{8'd127,8'd204} : s = 242;
	{8'd127,8'd205} : s = 108;
	{8'd127,8'd206} : s = 241;
	{8'd127,8'd207} : s = 236;
	{8'd127,8'd208} : s = 399;
	{8'd127,8'd209} : s = 26;
	{8'd127,8'd210} : s = 106;
	{8'd127,8'd211} : s = 105;
	{8'd127,8'd212} : s = 234;
	{8'd127,8'd213} : s = 102;
	{8'd127,8'd214} : s = 233;
	{8'd127,8'd215} : s = 230;
	{8'd127,8'd216} : s = 380;
	{8'd127,8'd217} : s = 101;
	{8'd127,8'd218} : s = 229;
	{8'd127,8'd219} : s = 227;
	{8'd127,8'd220} : s = 378;
	{8'd127,8'd221} : s = 220;
	{8'd127,8'd222} : s = 377;
	{8'd127,8'd223} : s = 374;
	{8'd127,8'd224} : s = 487;
	{8'd127,8'd225} : s = 25;
	{8'd127,8'd226} : s = 99;
	{8'd127,8'd227} : s = 92;
	{8'd127,8'd228} : s = 218;
	{8'd127,8'd229} : s = 90;
	{8'd127,8'd230} : s = 217;
	{8'd127,8'd231} : s = 214;
	{8'd127,8'd232} : s = 373;
	{8'd127,8'd233} : s = 89;
	{8'd127,8'd234} : s = 213;
	{8'd127,8'd235} : s = 211;
	{8'd127,8'd236} : s = 371;
	{8'd127,8'd237} : s = 206;
	{8'd127,8'd238} : s = 366;
	{8'd127,8'd239} : s = 365;
	{8'd127,8'd240} : s = 478;
	{8'd127,8'd241} : s = 86;
	{8'd127,8'd242} : s = 205;
	{8'd127,8'd243} : s = 203;
	{8'd127,8'd244} : s = 363;
	{8'd127,8'd245} : s = 199;
	{8'd127,8'd246} : s = 359;
	{8'd127,8'd247} : s = 350;
	{8'd127,8'd248} : s = 477;
	{8'd127,8'd249} : s = 188;
	{8'd127,8'd250} : s = 349;
	{8'd127,8'd251} : s = 347;
	{8'd127,8'd252} : s = 475;
	{8'd127,8'd253} : s = 343;
	{8'd127,8'd254} : s = 471;
	{8'd127,8'd255} : s = 463;
	{8'd128,8'd0} : s = 2;
	{8'd128,8'd1} : s = 48;
	{8'd128,8'd2} : s = 40;
	{8'd128,8'd3} : s = 168;
	{8'd128,8'd4} : s = 36;
	{8'd128,8'd5} : s = 164;
	{8'd128,8'd6} : s = 162;
	{8'd128,8'd7} : s = 323;
	{8'd128,8'd8} : s = 34;
	{8'd128,8'd9} : s = 161;
	{8'd128,8'd10} : s = 152;
	{8'd128,8'd11} : s = 312;
	{8'd128,8'd12} : s = 148;
	{8'd128,8'd13} : s = 308;
	{8'd128,8'd14} : s = 306;
	{8'd128,8'd15} : s = 425;
	{8'd128,8'd16} : s = 33;
	{8'd128,8'd17} : s = 146;
	{8'd128,8'd18} : s = 145;
	{8'd128,8'd19} : s = 305;
	{8'd128,8'd20} : s = 140;
	{8'd128,8'd21} : s = 300;
	{8'd128,8'd22} : s = 298;
	{8'd128,8'd23} : s = 422;
	{8'd128,8'd24} : s = 138;
	{8'd128,8'd25} : s = 297;
	{8'd128,8'd26} : s = 294;
	{8'd128,8'd27} : s = 421;
	{8'd128,8'd28} : s = 293;
	{8'd128,8'd29} : s = 419;
	{8'd128,8'd30} : s = 412;
	{8'd128,8'd31} : s = 486;
	{8'd128,8'd32} : s = 24;
	{8'd128,8'd33} : s = 137;
	{8'd128,8'd34} : s = 134;
	{8'd128,8'd35} : s = 291;
	{8'd128,8'd36} : s = 133;
	{8'd128,8'd37} : s = 284;
	{8'd128,8'd38} : s = 282;
	{8'd128,8'd39} : s = 410;
	{8'd128,8'd40} : s = 131;
	{8'd128,8'd41} : s = 281;
	{8'd128,8'd42} : s = 278;
	{8'd128,8'd43} : s = 409;
	{8'd128,8'd44} : s = 277;
	{8'd128,8'd45} : s = 406;
	{8'd128,8'd46} : s = 405;
	{8'd128,8'd47} : s = 485;
	{8'd128,8'd48} : s = 112;
	{8'd128,8'd49} : s = 275;
	{8'd128,8'd50} : s = 270;
	{8'd128,8'd51} : s = 403;
	{8'd128,8'd52} : s = 269;
	{8'd128,8'd53} : s = 398;
	{8'd128,8'd54} : s = 397;
	{8'd128,8'd55} : s = 483;
	{8'd128,8'd56} : s = 267;
	{8'd128,8'd57} : s = 395;
	{8'd128,8'd58} : s = 391;
	{8'd128,8'd59} : s = 476;
	{8'd128,8'd60} : s = 376;
	{8'd128,8'd61} : s = 474;
	{8'd128,8'd62} : s = 473;
	{8'd128,8'd63} : s = 506;
	{8'd128,8'd64} : s = 20;
	{8'd128,8'd65} : s = 104;
	{8'd128,8'd66} : s = 100;
	{8'd128,8'd67} : s = 263;
	{8'd128,8'd68} : s = 98;
	{8'd128,8'd69} : s = 240;
	{8'd128,8'd70} : s = 232;
	{8'd128,8'd71} : s = 372;
	{8'd128,8'd72} : s = 97;
	{8'd128,8'd73} : s = 228;
	{8'd128,8'd74} : s = 226;
	{8'd128,8'd75} : s = 370;
	{8'd128,8'd76} : s = 225;
	{8'd128,8'd77} : s = 369;
	{8'd128,8'd78} : s = 364;
	{8'd128,8'd79} : s = 470;
	{8'd128,8'd80} : s = 88;
	{8'd128,8'd81} : s = 216;
	{8'd128,8'd82} : s = 212;
	{8'd128,8'd83} : s = 362;
	{8'd128,8'd84} : s = 210;
	{8'd128,8'd85} : s = 361;
	{8'd128,8'd86} : s = 358;
	{8'd128,8'd87} : s = 469;
	{8'd128,8'd88} : s = 209;
	{8'd128,8'd89} : s = 357;
	{8'd128,8'd90} : s = 355;
	{8'd128,8'd91} : s = 467;
	{8'd128,8'd92} : s = 348;
	{8'd128,8'd93} : s = 462;
	{8'd128,8'd94} : s = 461;
	{8'd128,8'd95} : s = 505;
	{8'd128,8'd96} : s = 84;
	{8'd128,8'd97} : s = 204;
	{8'd128,8'd98} : s = 202;
	{8'd128,8'd99} : s = 346;
	{8'd128,8'd100} : s = 201;
	{8'd128,8'd101} : s = 345;
	{8'd128,8'd102} : s = 342;
	{8'd128,8'd103} : s = 459;
	{8'd128,8'd104} : s = 198;
	{8'd128,8'd105} : s = 341;
	{8'd128,8'd106} : s = 339;
	{8'd128,8'd107} : s = 455;
	{8'd128,8'd108} : s = 334;
	{8'd128,8'd109} : s = 444;
	{8'd128,8'd110} : s = 442;
	{8'd128,8'd111} : s = 502;
	{8'd128,8'd112} : s = 197;
	{8'd128,8'd113} : s = 333;
	{8'd128,8'd114} : s = 331;
	{8'd128,8'd115} : s = 441;
	{8'd128,8'd116} : s = 327;
	{8'd128,8'd117} : s = 438;
	{8'd128,8'd118} : s = 437;
	{8'd128,8'd119} : s = 501;
	{8'd128,8'd120} : s = 316;
	{8'd128,8'd121} : s = 435;
	{8'd128,8'd122} : s = 430;
	{8'd128,8'd123} : s = 499;
	{8'd128,8'd124} : s = 429;
	{8'd128,8'd125} : s = 494;
	{8'd128,8'd126} : s = 493;
	{8'd128,8'd127} : s = 510;
	{8'd128,8'd128} : s = 1;
	{8'd128,8'd129} : s = 18;
	{8'd128,8'd130} : s = 17;
	{8'd128,8'd131} : s = 82;
	{8'd128,8'd132} : s = 12;
	{8'd128,8'd133} : s = 81;
	{8'd128,8'd134} : s = 76;
	{8'd128,8'd135} : s = 195;
	{8'd128,8'd136} : s = 10;
	{8'd128,8'd137} : s = 74;
	{8'd128,8'd138} : s = 73;
	{8'd128,8'd139} : s = 184;
	{8'd128,8'd140} : s = 70;
	{8'd128,8'd141} : s = 180;
	{8'd128,8'd142} : s = 178;
	{8'd128,8'd143} : s = 314;
	{8'd128,8'd144} : s = 9;
	{8'd128,8'd145} : s = 69;
	{8'd128,8'd146} : s = 67;
	{8'd128,8'd147} : s = 177;
	{8'd128,8'd148} : s = 56;
	{8'd128,8'd149} : s = 172;
	{8'd128,8'd150} : s = 170;
	{8'd128,8'd151} : s = 313;
	{8'd128,8'd152} : s = 52;
	{8'd128,8'd153} : s = 169;
	{8'd128,8'd154} : s = 166;
	{8'd128,8'd155} : s = 310;
	{8'd128,8'd156} : s = 165;
	{8'd128,8'd157} : s = 309;
	{8'd128,8'd158} : s = 307;
	{8'd128,8'd159} : s = 427;
	{8'd128,8'd160} : s = 6;
	{8'd128,8'd161} : s = 50;
	{8'd128,8'd162} : s = 49;
	{8'd128,8'd163} : s = 163;
	{8'd128,8'd164} : s = 44;
	{8'd128,8'd165} : s = 156;
	{8'd128,8'd166} : s = 154;
	{8'd128,8'd167} : s = 302;
	{8'd128,8'd168} : s = 42;
	{8'd128,8'd169} : s = 153;
	{8'd128,8'd170} : s = 150;
	{8'd128,8'd171} : s = 301;
	{8'd128,8'd172} : s = 149;
	{8'd128,8'd173} : s = 299;
	{8'd128,8'd174} : s = 295;
	{8'd128,8'd175} : s = 423;
	{8'd128,8'd176} : s = 41;
	{8'd128,8'd177} : s = 147;
	{8'd128,8'd178} : s = 142;
	{8'd128,8'd179} : s = 286;
	{8'd128,8'd180} : s = 141;
	{8'd128,8'd181} : s = 285;
	{8'd128,8'd182} : s = 283;
	{8'd128,8'd183} : s = 414;
	{8'd128,8'd184} : s = 139;
	{8'd128,8'd185} : s = 279;
	{8'd128,8'd186} : s = 271;
	{8'd128,8'd187} : s = 413;
	{8'd128,8'd188} : s = 248;
	{8'd128,8'd189} : s = 411;
	{8'd128,8'd190} : s = 407;
	{8'd128,8'd191} : s = 491;
	{8'd128,8'd192} : s = 5;
	{8'd128,8'd193} : s = 38;
	{8'd128,8'd194} : s = 37;
	{8'd128,8'd195} : s = 135;
	{8'd128,8'd196} : s = 35;
	{8'd128,8'd197} : s = 120;
	{8'd128,8'd198} : s = 116;
	{8'd128,8'd199} : s = 244;
	{8'd128,8'd200} : s = 28;
	{8'd128,8'd201} : s = 114;
	{8'd128,8'd202} : s = 113;
	{8'd128,8'd203} : s = 242;
	{8'd128,8'd204} : s = 108;
	{8'd128,8'd205} : s = 241;
	{8'd128,8'd206} : s = 236;
	{8'd128,8'd207} : s = 399;
	{8'd128,8'd208} : s = 26;
	{8'd128,8'd209} : s = 106;
	{8'd128,8'd210} : s = 105;
	{8'd128,8'd211} : s = 234;
	{8'd128,8'd212} : s = 102;
	{8'd128,8'd213} : s = 233;
	{8'd128,8'd214} : s = 230;
	{8'd128,8'd215} : s = 380;
	{8'd128,8'd216} : s = 101;
	{8'd128,8'd217} : s = 229;
	{8'd128,8'd218} : s = 227;
	{8'd128,8'd219} : s = 378;
	{8'd128,8'd220} : s = 220;
	{8'd128,8'd221} : s = 377;
	{8'd128,8'd222} : s = 374;
	{8'd128,8'd223} : s = 487;
	{8'd128,8'd224} : s = 25;
	{8'd128,8'd225} : s = 99;
	{8'd128,8'd226} : s = 92;
	{8'd128,8'd227} : s = 218;
	{8'd128,8'd228} : s = 90;
	{8'd128,8'd229} : s = 217;
	{8'd128,8'd230} : s = 214;
	{8'd128,8'd231} : s = 373;
	{8'd128,8'd232} : s = 89;
	{8'd128,8'd233} : s = 213;
	{8'd128,8'd234} : s = 211;
	{8'd128,8'd235} : s = 371;
	{8'd128,8'd236} : s = 206;
	{8'd128,8'd237} : s = 366;
	{8'd128,8'd238} : s = 365;
	{8'd128,8'd239} : s = 478;
	{8'd128,8'd240} : s = 86;
	{8'd128,8'd241} : s = 205;
	{8'd128,8'd242} : s = 203;
	{8'd128,8'd243} : s = 363;
	{8'd128,8'd244} : s = 199;
	{8'd128,8'd245} : s = 359;
	{8'd128,8'd246} : s = 350;
	{8'd128,8'd247} : s = 477;
	{8'd128,8'd248} : s = 188;
	{8'd128,8'd249} : s = 349;
	{8'd128,8'd250} : s = 347;
	{8'd128,8'd251} : s = 475;
	{8'd128,8'd252} : s = 343;
	{8'd128,8'd253} : s = 471;
	{8'd128,8'd254} : s = 463;
	{8'd128,8'd255} : s = 509;
	{8'd129,8'd0} : s = 48;
	{8'd129,8'd1} : s = 40;
	{8'd129,8'd2} : s = 168;
	{8'd129,8'd3} : s = 36;
	{8'd129,8'd4} : s = 164;
	{8'd129,8'd5} : s = 162;
	{8'd129,8'd6} : s = 323;
	{8'd129,8'd7} : s = 34;
	{8'd129,8'd8} : s = 161;
	{8'd129,8'd9} : s = 152;
	{8'd129,8'd10} : s = 312;
	{8'd129,8'd11} : s = 148;
	{8'd129,8'd12} : s = 308;
	{8'd129,8'd13} : s = 306;
	{8'd129,8'd14} : s = 425;
	{8'd129,8'd15} : s = 33;
	{8'd129,8'd16} : s = 146;
	{8'd129,8'd17} : s = 145;
	{8'd129,8'd18} : s = 305;
	{8'd129,8'd19} : s = 140;
	{8'd129,8'd20} : s = 300;
	{8'd129,8'd21} : s = 298;
	{8'd129,8'd22} : s = 422;
	{8'd129,8'd23} : s = 138;
	{8'd129,8'd24} : s = 297;
	{8'd129,8'd25} : s = 294;
	{8'd129,8'd26} : s = 421;
	{8'd129,8'd27} : s = 293;
	{8'd129,8'd28} : s = 419;
	{8'd129,8'd29} : s = 412;
	{8'd129,8'd30} : s = 486;
	{8'd129,8'd31} : s = 24;
	{8'd129,8'd32} : s = 137;
	{8'd129,8'd33} : s = 134;
	{8'd129,8'd34} : s = 291;
	{8'd129,8'd35} : s = 133;
	{8'd129,8'd36} : s = 284;
	{8'd129,8'd37} : s = 282;
	{8'd129,8'd38} : s = 410;
	{8'd129,8'd39} : s = 131;
	{8'd129,8'd40} : s = 281;
	{8'd129,8'd41} : s = 278;
	{8'd129,8'd42} : s = 409;
	{8'd129,8'd43} : s = 277;
	{8'd129,8'd44} : s = 406;
	{8'd129,8'd45} : s = 405;
	{8'd129,8'd46} : s = 485;
	{8'd129,8'd47} : s = 112;
	{8'd129,8'd48} : s = 275;
	{8'd129,8'd49} : s = 270;
	{8'd129,8'd50} : s = 403;
	{8'd129,8'd51} : s = 269;
	{8'd129,8'd52} : s = 398;
	{8'd129,8'd53} : s = 397;
	{8'd129,8'd54} : s = 483;
	{8'd129,8'd55} : s = 267;
	{8'd129,8'd56} : s = 395;
	{8'd129,8'd57} : s = 391;
	{8'd129,8'd58} : s = 476;
	{8'd129,8'd59} : s = 376;
	{8'd129,8'd60} : s = 474;
	{8'd129,8'd61} : s = 473;
	{8'd129,8'd62} : s = 506;
	{8'd129,8'd63} : s = 20;
	{8'd129,8'd64} : s = 104;
	{8'd129,8'd65} : s = 100;
	{8'd129,8'd66} : s = 263;
	{8'd129,8'd67} : s = 98;
	{8'd129,8'd68} : s = 240;
	{8'd129,8'd69} : s = 232;
	{8'd129,8'd70} : s = 372;
	{8'd129,8'd71} : s = 97;
	{8'd129,8'd72} : s = 228;
	{8'd129,8'd73} : s = 226;
	{8'd129,8'd74} : s = 370;
	{8'd129,8'd75} : s = 225;
	{8'd129,8'd76} : s = 369;
	{8'd129,8'd77} : s = 364;
	{8'd129,8'd78} : s = 470;
	{8'd129,8'd79} : s = 88;
	{8'd129,8'd80} : s = 216;
	{8'd129,8'd81} : s = 212;
	{8'd129,8'd82} : s = 362;
	{8'd129,8'd83} : s = 210;
	{8'd129,8'd84} : s = 361;
	{8'd129,8'd85} : s = 358;
	{8'd129,8'd86} : s = 469;
	{8'd129,8'd87} : s = 209;
	{8'd129,8'd88} : s = 357;
	{8'd129,8'd89} : s = 355;
	{8'd129,8'd90} : s = 467;
	{8'd129,8'd91} : s = 348;
	{8'd129,8'd92} : s = 462;
	{8'd129,8'd93} : s = 461;
	{8'd129,8'd94} : s = 505;
	{8'd129,8'd95} : s = 84;
	{8'd129,8'd96} : s = 204;
	{8'd129,8'd97} : s = 202;
	{8'd129,8'd98} : s = 346;
	{8'd129,8'd99} : s = 201;
	{8'd129,8'd100} : s = 345;
	{8'd129,8'd101} : s = 342;
	{8'd129,8'd102} : s = 459;
	{8'd129,8'd103} : s = 198;
	{8'd129,8'd104} : s = 341;
	{8'd129,8'd105} : s = 339;
	{8'd129,8'd106} : s = 455;
	{8'd129,8'd107} : s = 334;
	{8'd129,8'd108} : s = 444;
	{8'd129,8'd109} : s = 442;
	{8'd129,8'd110} : s = 502;
	{8'd129,8'd111} : s = 197;
	{8'd129,8'd112} : s = 333;
	{8'd129,8'd113} : s = 331;
	{8'd129,8'd114} : s = 441;
	{8'd129,8'd115} : s = 327;
	{8'd129,8'd116} : s = 438;
	{8'd129,8'd117} : s = 437;
	{8'd129,8'd118} : s = 501;
	{8'd129,8'd119} : s = 316;
	{8'd129,8'd120} : s = 435;
	{8'd129,8'd121} : s = 430;
	{8'd129,8'd122} : s = 499;
	{8'd129,8'd123} : s = 429;
	{8'd129,8'd124} : s = 494;
	{8'd129,8'd125} : s = 493;
	{8'd129,8'd126} : s = 510;
	{8'd129,8'd127} : s = 1;
	{8'd129,8'd128} : s = 18;
	{8'd129,8'd129} : s = 17;
	{8'd129,8'd130} : s = 82;
	{8'd129,8'd131} : s = 12;
	{8'd129,8'd132} : s = 81;
	{8'd129,8'd133} : s = 76;
	{8'd129,8'd134} : s = 195;
	{8'd129,8'd135} : s = 10;
	{8'd129,8'd136} : s = 74;
	{8'd129,8'd137} : s = 73;
	{8'd129,8'd138} : s = 184;
	{8'd129,8'd139} : s = 70;
	{8'd129,8'd140} : s = 180;
	{8'd129,8'd141} : s = 178;
	{8'd129,8'd142} : s = 314;
	{8'd129,8'd143} : s = 9;
	{8'd129,8'd144} : s = 69;
	{8'd129,8'd145} : s = 67;
	{8'd129,8'd146} : s = 177;
	{8'd129,8'd147} : s = 56;
	{8'd129,8'd148} : s = 172;
	{8'd129,8'd149} : s = 170;
	{8'd129,8'd150} : s = 313;
	{8'd129,8'd151} : s = 52;
	{8'd129,8'd152} : s = 169;
	{8'd129,8'd153} : s = 166;
	{8'd129,8'd154} : s = 310;
	{8'd129,8'd155} : s = 165;
	{8'd129,8'd156} : s = 309;
	{8'd129,8'd157} : s = 307;
	{8'd129,8'd158} : s = 427;
	{8'd129,8'd159} : s = 6;
	{8'd129,8'd160} : s = 50;
	{8'd129,8'd161} : s = 49;
	{8'd129,8'd162} : s = 163;
	{8'd129,8'd163} : s = 44;
	{8'd129,8'd164} : s = 156;
	{8'd129,8'd165} : s = 154;
	{8'd129,8'd166} : s = 302;
	{8'd129,8'd167} : s = 42;
	{8'd129,8'd168} : s = 153;
	{8'd129,8'd169} : s = 150;
	{8'd129,8'd170} : s = 301;
	{8'd129,8'd171} : s = 149;
	{8'd129,8'd172} : s = 299;
	{8'd129,8'd173} : s = 295;
	{8'd129,8'd174} : s = 423;
	{8'd129,8'd175} : s = 41;
	{8'd129,8'd176} : s = 147;
	{8'd129,8'd177} : s = 142;
	{8'd129,8'd178} : s = 286;
	{8'd129,8'd179} : s = 141;
	{8'd129,8'd180} : s = 285;
	{8'd129,8'd181} : s = 283;
	{8'd129,8'd182} : s = 414;
	{8'd129,8'd183} : s = 139;
	{8'd129,8'd184} : s = 279;
	{8'd129,8'd185} : s = 271;
	{8'd129,8'd186} : s = 413;
	{8'd129,8'd187} : s = 248;
	{8'd129,8'd188} : s = 411;
	{8'd129,8'd189} : s = 407;
	{8'd129,8'd190} : s = 491;
	{8'd129,8'd191} : s = 5;
	{8'd129,8'd192} : s = 38;
	{8'd129,8'd193} : s = 37;
	{8'd129,8'd194} : s = 135;
	{8'd129,8'd195} : s = 35;
	{8'd129,8'd196} : s = 120;
	{8'd129,8'd197} : s = 116;
	{8'd129,8'd198} : s = 244;
	{8'd129,8'd199} : s = 28;
	{8'd129,8'd200} : s = 114;
	{8'd129,8'd201} : s = 113;
	{8'd129,8'd202} : s = 242;
	{8'd129,8'd203} : s = 108;
	{8'd129,8'd204} : s = 241;
	{8'd129,8'd205} : s = 236;
	{8'd129,8'd206} : s = 399;
	{8'd129,8'd207} : s = 26;
	{8'd129,8'd208} : s = 106;
	{8'd129,8'd209} : s = 105;
	{8'd129,8'd210} : s = 234;
	{8'd129,8'd211} : s = 102;
	{8'd129,8'd212} : s = 233;
	{8'd129,8'd213} : s = 230;
	{8'd129,8'd214} : s = 380;
	{8'd129,8'd215} : s = 101;
	{8'd129,8'd216} : s = 229;
	{8'd129,8'd217} : s = 227;
	{8'd129,8'd218} : s = 378;
	{8'd129,8'd219} : s = 220;
	{8'd129,8'd220} : s = 377;
	{8'd129,8'd221} : s = 374;
	{8'd129,8'd222} : s = 487;
	{8'd129,8'd223} : s = 25;
	{8'd129,8'd224} : s = 99;
	{8'd129,8'd225} : s = 92;
	{8'd129,8'd226} : s = 218;
	{8'd129,8'd227} : s = 90;
	{8'd129,8'd228} : s = 217;
	{8'd129,8'd229} : s = 214;
	{8'd129,8'd230} : s = 373;
	{8'd129,8'd231} : s = 89;
	{8'd129,8'd232} : s = 213;
	{8'd129,8'd233} : s = 211;
	{8'd129,8'd234} : s = 371;
	{8'd129,8'd235} : s = 206;
	{8'd129,8'd236} : s = 366;
	{8'd129,8'd237} : s = 365;
	{8'd129,8'd238} : s = 478;
	{8'd129,8'd239} : s = 86;
	{8'd129,8'd240} : s = 205;
	{8'd129,8'd241} : s = 203;
	{8'd129,8'd242} : s = 363;
	{8'd129,8'd243} : s = 199;
	{8'd129,8'd244} : s = 359;
	{8'd129,8'd245} : s = 350;
	{8'd129,8'd246} : s = 477;
	{8'd129,8'd247} : s = 188;
	{8'd129,8'd248} : s = 349;
	{8'd129,8'd249} : s = 347;
	{8'd129,8'd250} : s = 475;
	{8'd129,8'd251} : s = 343;
	{8'd129,8'd252} : s = 471;
	{8'd129,8'd253} : s = 463;
	{8'd129,8'd254} : s = 509;
	{8'd129,8'd255} : s = 3;
	{8'd130,8'd0} : s = 40;
	{8'd130,8'd1} : s = 168;
	{8'd130,8'd2} : s = 36;
	{8'd130,8'd3} : s = 164;
	{8'd130,8'd4} : s = 162;
	{8'd130,8'd5} : s = 323;
	{8'd130,8'd6} : s = 34;
	{8'd130,8'd7} : s = 161;
	{8'd130,8'd8} : s = 152;
	{8'd130,8'd9} : s = 312;
	{8'd130,8'd10} : s = 148;
	{8'd130,8'd11} : s = 308;
	{8'd130,8'd12} : s = 306;
	{8'd130,8'd13} : s = 425;
	{8'd130,8'd14} : s = 33;
	{8'd130,8'd15} : s = 146;
	{8'd130,8'd16} : s = 145;
	{8'd130,8'd17} : s = 305;
	{8'd130,8'd18} : s = 140;
	{8'd130,8'd19} : s = 300;
	{8'd130,8'd20} : s = 298;
	{8'd130,8'd21} : s = 422;
	{8'd130,8'd22} : s = 138;
	{8'd130,8'd23} : s = 297;
	{8'd130,8'd24} : s = 294;
	{8'd130,8'd25} : s = 421;
	{8'd130,8'd26} : s = 293;
	{8'd130,8'd27} : s = 419;
	{8'd130,8'd28} : s = 412;
	{8'd130,8'd29} : s = 486;
	{8'd130,8'd30} : s = 24;
	{8'd130,8'd31} : s = 137;
	{8'd130,8'd32} : s = 134;
	{8'd130,8'd33} : s = 291;
	{8'd130,8'd34} : s = 133;
	{8'd130,8'd35} : s = 284;
	{8'd130,8'd36} : s = 282;
	{8'd130,8'd37} : s = 410;
	{8'd130,8'd38} : s = 131;
	{8'd130,8'd39} : s = 281;
	{8'd130,8'd40} : s = 278;
	{8'd130,8'd41} : s = 409;
	{8'd130,8'd42} : s = 277;
	{8'd130,8'd43} : s = 406;
	{8'd130,8'd44} : s = 405;
	{8'd130,8'd45} : s = 485;
	{8'd130,8'd46} : s = 112;
	{8'd130,8'd47} : s = 275;
	{8'd130,8'd48} : s = 270;
	{8'd130,8'd49} : s = 403;
	{8'd130,8'd50} : s = 269;
	{8'd130,8'd51} : s = 398;
	{8'd130,8'd52} : s = 397;
	{8'd130,8'd53} : s = 483;
	{8'd130,8'd54} : s = 267;
	{8'd130,8'd55} : s = 395;
	{8'd130,8'd56} : s = 391;
	{8'd130,8'd57} : s = 476;
	{8'd130,8'd58} : s = 376;
	{8'd130,8'd59} : s = 474;
	{8'd130,8'd60} : s = 473;
	{8'd130,8'd61} : s = 506;
	{8'd130,8'd62} : s = 20;
	{8'd130,8'd63} : s = 104;
	{8'd130,8'd64} : s = 100;
	{8'd130,8'd65} : s = 263;
	{8'd130,8'd66} : s = 98;
	{8'd130,8'd67} : s = 240;
	{8'd130,8'd68} : s = 232;
	{8'd130,8'd69} : s = 372;
	{8'd130,8'd70} : s = 97;
	{8'd130,8'd71} : s = 228;
	{8'd130,8'd72} : s = 226;
	{8'd130,8'd73} : s = 370;
	{8'd130,8'd74} : s = 225;
	{8'd130,8'd75} : s = 369;
	{8'd130,8'd76} : s = 364;
	{8'd130,8'd77} : s = 470;
	{8'd130,8'd78} : s = 88;
	{8'd130,8'd79} : s = 216;
	{8'd130,8'd80} : s = 212;
	{8'd130,8'd81} : s = 362;
	{8'd130,8'd82} : s = 210;
	{8'd130,8'd83} : s = 361;
	{8'd130,8'd84} : s = 358;
	{8'd130,8'd85} : s = 469;
	{8'd130,8'd86} : s = 209;
	{8'd130,8'd87} : s = 357;
	{8'd130,8'd88} : s = 355;
	{8'd130,8'd89} : s = 467;
	{8'd130,8'd90} : s = 348;
	{8'd130,8'd91} : s = 462;
	{8'd130,8'd92} : s = 461;
	{8'd130,8'd93} : s = 505;
	{8'd130,8'd94} : s = 84;
	{8'd130,8'd95} : s = 204;
	{8'd130,8'd96} : s = 202;
	{8'd130,8'd97} : s = 346;
	{8'd130,8'd98} : s = 201;
	{8'd130,8'd99} : s = 345;
	{8'd130,8'd100} : s = 342;
	{8'd130,8'd101} : s = 459;
	{8'd130,8'd102} : s = 198;
	{8'd130,8'd103} : s = 341;
	{8'd130,8'd104} : s = 339;
	{8'd130,8'd105} : s = 455;
	{8'd130,8'd106} : s = 334;
	{8'd130,8'd107} : s = 444;
	{8'd130,8'd108} : s = 442;
	{8'd130,8'd109} : s = 502;
	{8'd130,8'd110} : s = 197;
	{8'd130,8'd111} : s = 333;
	{8'd130,8'd112} : s = 331;
	{8'd130,8'd113} : s = 441;
	{8'd130,8'd114} : s = 327;
	{8'd130,8'd115} : s = 438;
	{8'd130,8'd116} : s = 437;
	{8'd130,8'd117} : s = 501;
	{8'd130,8'd118} : s = 316;
	{8'd130,8'd119} : s = 435;
	{8'd130,8'd120} : s = 430;
	{8'd130,8'd121} : s = 499;
	{8'd130,8'd122} : s = 429;
	{8'd130,8'd123} : s = 494;
	{8'd130,8'd124} : s = 493;
	{8'd130,8'd125} : s = 510;
	{8'd130,8'd126} : s = 1;
	{8'd130,8'd127} : s = 18;
	{8'd130,8'd128} : s = 17;
	{8'd130,8'd129} : s = 82;
	{8'd130,8'd130} : s = 12;
	{8'd130,8'd131} : s = 81;
	{8'd130,8'd132} : s = 76;
	{8'd130,8'd133} : s = 195;
	{8'd130,8'd134} : s = 10;
	{8'd130,8'd135} : s = 74;
	{8'd130,8'd136} : s = 73;
	{8'd130,8'd137} : s = 184;
	{8'd130,8'd138} : s = 70;
	{8'd130,8'd139} : s = 180;
	{8'd130,8'd140} : s = 178;
	{8'd130,8'd141} : s = 314;
	{8'd130,8'd142} : s = 9;
	{8'd130,8'd143} : s = 69;
	{8'd130,8'd144} : s = 67;
	{8'd130,8'd145} : s = 177;
	{8'd130,8'd146} : s = 56;
	{8'd130,8'd147} : s = 172;
	{8'd130,8'd148} : s = 170;
	{8'd130,8'd149} : s = 313;
	{8'd130,8'd150} : s = 52;
	{8'd130,8'd151} : s = 169;
	{8'd130,8'd152} : s = 166;
	{8'd130,8'd153} : s = 310;
	{8'd130,8'd154} : s = 165;
	{8'd130,8'd155} : s = 309;
	{8'd130,8'd156} : s = 307;
	{8'd130,8'd157} : s = 427;
	{8'd130,8'd158} : s = 6;
	{8'd130,8'd159} : s = 50;
	{8'd130,8'd160} : s = 49;
	{8'd130,8'd161} : s = 163;
	{8'd130,8'd162} : s = 44;
	{8'd130,8'd163} : s = 156;
	{8'd130,8'd164} : s = 154;
	{8'd130,8'd165} : s = 302;
	{8'd130,8'd166} : s = 42;
	{8'd130,8'd167} : s = 153;
	{8'd130,8'd168} : s = 150;
	{8'd130,8'd169} : s = 301;
	{8'd130,8'd170} : s = 149;
	{8'd130,8'd171} : s = 299;
	{8'd130,8'd172} : s = 295;
	{8'd130,8'd173} : s = 423;
	{8'd130,8'd174} : s = 41;
	{8'd130,8'd175} : s = 147;
	{8'd130,8'd176} : s = 142;
	{8'd130,8'd177} : s = 286;
	{8'd130,8'd178} : s = 141;
	{8'd130,8'd179} : s = 285;
	{8'd130,8'd180} : s = 283;
	{8'd130,8'd181} : s = 414;
	{8'd130,8'd182} : s = 139;
	{8'd130,8'd183} : s = 279;
	{8'd130,8'd184} : s = 271;
	{8'd130,8'd185} : s = 413;
	{8'd130,8'd186} : s = 248;
	{8'd130,8'd187} : s = 411;
	{8'd130,8'd188} : s = 407;
	{8'd130,8'd189} : s = 491;
	{8'd130,8'd190} : s = 5;
	{8'd130,8'd191} : s = 38;
	{8'd130,8'd192} : s = 37;
	{8'd130,8'd193} : s = 135;
	{8'd130,8'd194} : s = 35;
	{8'd130,8'd195} : s = 120;
	{8'd130,8'd196} : s = 116;
	{8'd130,8'd197} : s = 244;
	{8'd130,8'd198} : s = 28;
	{8'd130,8'd199} : s = 114;
	{8'd130,8'd200} : s = 113;
	{8'd130,8'd201} : s = 242;
	{8'd130,8'd202} : s = 108;
	{8'd130,8'd203} : s = 241;
	{8'd130,8'd204} : s = 236;
	{8'd130,8'd205} : s = 399;
	{8'd130,8'd206} : s = 26;
	{8'd130,8'd207} : s = 106;
	{8'd130,8'd208} : s = 105;
	{8'd130,8'd209} : s = 234;
	{8'd130,8'd210} : s = 102;
	{8'd130,8'd211} : s = 233;
	{8'd130,8'd212} : s = 230;
	{8'd130,8'd213} : s = 380;
	{8'd130,8'd214} : s = 101;
	{8'd130,8'd215} : s = 229;
	{8'd130,8'd216} : s = 227;
	{8'd130,8'd217} : s = 378;
	{8'd130,8'd218} : s = 220;
	{8'd130,8'd219} : s = 377;
	{8'd130,8'd220} : s = 374;
	{8'd130,8'd221} : s = 487;
	{8'd130,8'd222} : s = 25;
	{8'd130,8'd223} : s = 99;
	{8'd130,8'd224} : s = 92;
	{8'd130,8'd225} : s = 218;
	{8'd130,8'd226} : s = 90;
	{8'd130,8'd227} : s = 217;
	{8'd130,8'd228} : s = 214;
	{8'd130,8'd229} : s = 373;
	{8'd130,8'd230} : s = 89;
	{8'd130,8'd231} : s = 213;
	{8'd130,8'd232} : s = 211;
	{8'd130,8'd233} : s = 371;
	{8'd130,8'd234} : s = 206;
	{8'd130,8'd235} : s = 366;
	{8'd130,8'd236} : s = 365;
	{8'd130,8'd237} : s = 478;
	{8'd130,8'd238} : s = 86;
	{8'd130,8'd239} : s = 205;
	{8'd130,8'd240} : s = 203;
	{8'd130,8'd241} : s = 363;
	{8'd130,8'd242} : s = 199;
	{8'd130,8'd243} : s = 359;
	{8'd130,8'd244} : s = 350;
	{8'd130,8'd245} : s = 477;
	{8'd130,8'd246} : s = 188;
	{8'd130,8'd247} : s = 349;
	{8'd130,8'd248} : s = 347;
	{8'd130,8'd249} : s = 475;
	{8'd130,8'd250} : s = 343;
	{8'd130,8'd251} : s = 471;
	{8'd130,8'd252} : s = 463;
	{8'd130,8'd253} : s = 509;
	{8'd130,8'd254} : s = 3;
	{8'd130,8'd255} : s = 22;
	{8'd131,8'd0} : s = 168;
	{8'd131,8'd1} : s = 36;
	{8'd131,8'd2} : s = 164;
	{8'd131,8'd3} : s = 162;
	{8'd131,8'd4} : s = 323;
	{8'd131,8'd5} : s = 34;
	{8'd131,8'd6} : s = 161;
	{8'd131,8'd7} : s = 152;
	{8'd131,8'd8} : s = 312;
	{8'd131,8'd9} : s = 148;
	{8'd131,8'd10} : s = 308;
	{8'd131,8'd11} : s = 306;
	{8'd131,8'd12} : s = 425;
	{8'd131,8'd13} : s = 33;
	{8'd131,8'd14} : s = 146;
	{8'd131,8'd15} : s = 145;
	{8'd131,8'd16} : s = 305;
	{8'd131,8'd17} : s = 140;
	{8'd131,8'd18} : s = 300;
	{8'd131,8'd19} : s = 298;
	{8'd131,8'd20} : s = 422;
	{8'd131,8'd21} : s = 138;
	{8'd131,8'd22} : s = 297;
	{8'd131,8'd23} : s = 294;
	{8'd131,8'd24} : s = 421;
	{8'd131,8'd25} : s = 293;
	{8'd131,8'd26} : s = 419;
	{8'd131,8'd27} : s = 412;
	{8'd131,8'd28} : s = 486;
	{8'd131,8'd29} : s = 24;
	{8'd131,8'd30} : s = 137;
	{8'd131,8'd31} : s = 134;
	{8'd131,8'd32} : s = 291;
	{8'd131,8'd33} : s = 133;
	{8'd131,8'd34} : s = 284;
	{8'd131,8'd35} : s = 282;
	{8'd131,8'd36} : s = 410;
	{8'd131,8'd37} : s = 131;
	{8'd131,8'd38} : s = 281;
	{8'd131,8'd39} : s = 278;
	{8'd131,8'd40} : s = 409;
	{8'd131,8'd41} : s = 277;
	{8'd131,8'd42} : s = 406;
	{8'd131,8'd43} : s = 405;
	{8'd131,8'd44} : s = 485;
	{8'd131,8'd45} : s = 112;
	{8'd131,8'd46} : s = 275;
	{8'd131,8'd47} : s = 270;
	{8'd131,8'd48} : s = 403;
	{8'd131,8'd49} : s = 269;
	{8'd131,8'd50} : s = 398;
	{8'd131,8'd51} : s = 397;
	{8'd131,8'd52} : s = 483;
	{8'd131,8'd53} : s = 267;
	{8'd131,8'd54} : s = 395;
	{8'd131,8'd55} : s = 391;
	{8'd131,8'd56} : s = 476;
	{8'd131,8'd57} : s = 376;
	{8'd131,8'd58} : s = 474;
	{8'd131,8'd59} : s = 473;
	{8'd131,8'd60} : s = 506;
	{8'd131,8'd61} : s = 20;
	{8'd131,8'd62} : s = 104;
	{8'd131,8'd63} : s = 100;
	{8'd131,8'd64} : s = 263;
	{8'd131,8'd65} : s = 98;
	{8'd131,8'd66} : s = 240;
	{8'd131,8'd67} : s = 232;
	{8'd131,8'd68} : s = 372;
	{8'd131,8'd69} : s = 97;
	{8'd131,8'd70} : s = 228;
	{8'd131,8'd71} : s = 226;
	{8'd131,8'd72} : s = 370;
	{8'd131,8'd73} : s = 225;
	{8'd131,8'd74} : s = 369;
	{8'd131,8'd75} : s = 364;
	{8'd131,8'd76} : s = 470;
	{8'd131,8'd77} : s = 88;
	{8'd131,8'd78} : s = 216;
	{8'd131,8'd79} : s = 212;
	{8'd131,8'd80} : s = 362;
	{8'd131,8'd81} : s = 210;
	{8'd131,8'd82} : s = 361;
	{8'd131,8'd83} : s = 358;
	{8'd131,8'd84} : s = 469;
	{8'd131,8'd85} : s = 209;
	{8'd131,8'd86} : s = 357;
	{8'd131,8'd87} : s = 355;
	{8'd131,8'd88} : s = 467;
	{8'd131,8'd89} : s = 348;
	{8'd131,8'd90} : s = 462;
	{8'd131,8'd91} : s = 461;
	{8'd131,8'd92} : s = 505;
	{8'd131,8'd93} : s = 84;
	{8'd131,8'd94} : s = 204;
	{8'd131,8'd95} : s = 202;
	{8'd131,8'd96} : s = 346;
	{8'd131,8'd97} : s = 201;
	{8'd131,8'd98} : s = 345;
	{8'd131,8'd99} : s = 342;
	{8'd131,8'd100} : s = 459;
	{8'd131,8'd101} : s = 198;
	{8'd131,8'd102} : s = 341;
	{8'd131,8'd103} : s = 339;
	{8'd131,8'd104} : s = 455;
	{8'd131,8'd105} : s = 334;
	{8'd131,8'd106} : s = 444;
	{8'd131,8'd107} : s = 442;
	{8'd131,8'd108} : s = 502;
	{8'd131,8'd109} : s = 197;
	{8'd131,8'd110} : s = 333;
	{8'd131,8'd111} : s = 331;
	{8'd131,8'd112} : s = 441;
	{8'd131,8'd113} : s = 327;
	{8'd131,8'd114} : s = 438;
	{8'd131,8'd115} : s = 437;
	{8'd131,8'd116} : s = 501;
	{8'd131,8'd117} : s = 316;
	{8'd131,8'd118} : s = 435;
	{8'd131,8'd119} : s = 430;
	{8'd131,8'd120} : s = 499;
	{8'd131,8'd121} : s = 429;
	{8'd131,8'd122} : s = 494;
	{8'd131,8'd123} : s = 493;
	{8'd131,8'd124} : s = 510;
	{8'd131,8'd125} : s = 1;
	{8'd131,8'd126} : s = 18;
	{8'd131,8'd127} : s = 17;
	{8'd131,8'd128} : s = 82;
	{8'd131,8'd129} : s = 12;
	{8'd131,8'd130} : s = 81;
	{8'd131,8'd131} : s = 76;
	{8'd131,8'd132} : s = 195;
	{8'd131,8'd133} : s = 10;
	{8'd131,8'd134} : s = 74;
	{8'd131,8'd135} : s = 73;
	{8'd131,8'd136} : s = 184;
	{8'd131,8'd137} : s = 70;
	{8'd131,8'd138} : s = 180;
	{8'd131,8'd139} : s = 178;
	{8'd131,8'd140} : s = 314;
	{8'd131,8'd141} : s = 9;
	{8'd131,8'd142} : s = 69;
	{8'd131,8'd143} : s = 67;
	{8'd131,8'd144} : s = 177;
	{8'd131,8'd145} : s = 56;
	{8'd131,8'd146} : s = 172;
	{8'd131,8'd147} : s = 170;
	{8'd131,8'd148} : s = 313;
	{8'd131,8'd149} : s = 52;
	{8'd131,8'd150} : s = 169;
	{8'd131,8'd151} : s = 166;
	{8'd131,8'd152} : s = 310;
	{8'd131,8'd153} : s = 165;
	{8'd131,8'd154} : s = 309;
	{8'd131,8'd155} : s = 307;
	{8'd131,8'd156} : s = 427;
	{8'd131,8'd157} : s = 6;
	{8'd131,8'd158} : s = 50;
	{8'd131,8'd159} : s = 49;
	{8'd131,8'd160} : s = 163;
	{8'd131,8'd161} : s = 44;
	{8'd131,8'd162} : s = 156;
	{8'd131,8'd163} : s = 154;
	{8'd131,8'd164} : s = 302;
	{8'd131,8'd165} : s = 42;
	{8'd131,8'd166} : s = 153;
	{8'd131,8'd167} : s = 150;
	{8'd131,8'd168} : s = 301;
	{8'd131,8'd169} : s = 149;
	{8'd131,8'd170} : s = 299;
	{8'd131,8'd171} : s = 295;
	{8'd131,8'd172} : s = 423;
	{8'd131,8'd173} : s = 41;
	{8'd131,8'd174} : s = 147;
	{8'd131,8'd175} : s = 142;
	{8'd131,8'd176} : s = 286;
	{8'd131,8'd177} : s = 141;
	{8'd131,8'd178} : s = 285;
	{8'd131,8'd179} : s = 283;
	{8'd131,8'd180} : s = 414;
	{8'd131,8'd181} : s = 139;
	{8'd131,8'd182} : s = 279;
	{8'd131,8'd183} : s = 271;
	{8'd131,8'd184} : s = 413;
	{8'd131,8'd185} : s = 248;
	{8'd131,8'd186} : s = 411;
	{8'd131,8'd187} : s = 407;
	{8'd131,8'd188} : s = 491;
	{8'd131,8'd189} : s = 5;
	{8'd131,8'd190} : s = 38;
	{8'd131,8'd191} : s = 37;
	{8'd131,8'd192} : s = 135;
	{8'd131,8'd193} : s = 35;
	{8'd131,8'd194} : s = 120;
	{8'd131,8'd195} : s = 116;
	{8'd131,8'd196} : s = 244;
	{8'd131,8'd197} : s = 28;
	{8'd131,8'd198} : s = 114;
	{8'd131,8'd199} : s = 113;
	{8'd131,8'd200} : s = 242;
	{8'd131,8'd201} : s = 108;
	{8'd131,8'd202} : s = 241;
	{8'd131,8'd203} : s = 236;
	{8'd131,8'd204} : s = 399;
	{8'd131,8'd205} : s = 26;
	{8'd131,8'd206} : s = 106;
	{8'd131,8'd207} : s = 105;
	{8'd131,8'd208} : s = 234;
	{8'd131,8'd209} : s = 102;
	{8'd131,8'd210} : s = 233;
	{8'd131,8'd211} : s = 230;
	{8'd131,8'd212} : s = 380;
	{8'd131,8'd213} : s = 101;
	{8'd131,8'd214} : s = 229;
	{8'd131,8'd215} : s = 227;
	{8'd131,8'd216} : s = 378;
	{8'd131,8'd217} : s = 220;
	{8'd131,8'd218} : s = 377;
	{8'd131,8'd219} : s = 374;
	{8'd131,8'd220} : s = 487;
	{8'd131,8'd221} : s = 25;
	{8'd131,8'd222} : s = 99;
	{8'd131,8'd223} : s = 92;
	{8'd131,8'd224} : s = 218;
	{8'd131,8'd225} : s = 90;
	{8'd131,8'd226} : s = 217;
	{8'd131,8'd227} : s = 214;
	{8'd131,8'd228} : s = 373;
	{8'd131,8'd229} : s = 89;
	{8'd131,8'd230} : s = 213;
	{8'd131,8'd231} : s = 211;
	{8'd131,8'd232} : s = 371;
	{8'd131,8'd233} : s = 206;
	{8'd131,8'd234} : s = 366;
	{8'd131,8'd235} : s = 365;
	{8'd131,8'd236} : s = 478;
	{8'd131,8'd237} : s = 86;
	{8'd131,8'd238} : s = 205;
	{8'd131,8'd239} : s = 203;
	{8'd131,8'd240} : s = 363;
	{8'd131,8'd241} : s = 199;
	{8'd131,8'd242} : s = 359;
	{8'd131,8'd243} : s = 350;
	{8'd131,8'd244} : s = 477;
	{8'd131,8'd245} : s = 188;
	{8'd131,8'd246} : s = 349;
	{8'd131,8'd247} : s = 347;
	{8'd131,8'd248} : s = 475;
	{8'd131,8'd249} : s = 343;
	{8'd131,8'd250} : s = 471;
	{8'd131,8'd251} : s = 463;
	{8'd131,8'd252} : s = 509;
	{8'd131,8'd253} : s = 3;
	{8'd131,8'd254} : s = 22;
	{8'd131,8'd255} : s = 21;
	{8'd132,8'd0} : s = 36;
	{8'd132,8'd1} : s = 164;
	{8'd132,8'd2} : s = 162;
	{8'd132,8'd3} : s = 323;
	{8'd132,8'd4} : s = 34;
	{8'd132,8'd5} : s = 161;
	{8'd132,8'd6} : s = 152;
	{8'd132,8'd7} : s = 312;
	{8'd132,8'd8} : s = 148;
	{8'd132,8'd9} : s = 308;
	{8'd132,8'd10} : s = 306;
	{8'd132,8'd11} : s = 425;
	{8'd132,8'd12} : s = 33;
	{8'd132,8'd13} : s = 146;
	{8'd132,8'd14} : s = 145;
	{8'd132,8'd15} : s = 305;
	{8'd132,8'd16} : s = 140;
	{8'd132,8'd17} : s = 300;
	{8'd132,8'd18} : s = 298;
	{8'd132,8'd19} : s = 422;
	{8'd132,8'd20} : s = 138;
	{8'd132,8'd21} : s = 297;
	{8'd132,8'd22} : s = 294;
	{8'd132,8'd23} : s = 421;
	{8'd132,8'd24} : s = 293;
	{8'd132,8'd25} : s = 419;
	{8'd132,8'd26} : s = 412;
	{8'd132,8'd27} : s = 486;
	{8'd132,8'd28} : s = 24;
	{8'd132,8'd29} : s = 137;
	{8'd132,8'd30} : s = 134;
	{8'd132,8'd31} : s = 291;
	{8'd132,8'd32} : s = 133;
	{8'd132,8'd33} : s = 284;
	{8'd132,8'd34} : s = 282;
	{8'd132,8'd35} : s = 410;
	{8'd132,8'd36} : s = 131;
	{8'd132,8'd37} : s = 281;
	{8'd132,8'd38} : s = 278;
	{8'd132,8'd39} : s = 409;
	{8'd132,8'd40} : s = 277;
	{8'd132,8'd41} : s = 406;
	{8'd132,8'd42} : s = 405;
	{8'd132,8'd43} : s = 485;
	{8'd132,8'd44} : s = 112;
	{8'd132,8'd45} : s = 275;
	{8'd132,8'd46} : s = 270;
	{8'd132,8'd47} : s = 403;
	{8'd132,8'd48} : s = 269;
	{8'd132,8'd49} : s = 398;
	{8'd132,8'd50} : s = 397;
	{8'd132,8'd51} : s = 483;
	{8'd132,8'd52} : s = 267;
	{8'd132,8'd53} : s = 395;
	{8'd132,8'd54} : s = 391;
	{8'd132,8'd55} : s = 476;
	{8'd132,8'd56} : s = 376;
	{8'd132,8'd57} : s = 474;
	{8'd132,8'd58} : s = 473;
	{8'd132,8'd59} : s = 506;
	{8'd132,8'd60} : s = 20;
	{8'd132,8'd61} : s = 104;
	{8'd132,8'd62} : s = 100;
	{8'd132,8'd63} : s = 263;
	{8'd132,8'd64} : s = 98;
	{8'd132,8'd65} : s = 240;
	{8'd132,8'd66} : s = 232;
	{8'd132,8'd67} : s = 372;
	{8'd132,8'd68} : s = 97;
	{8'd132,8'd69} : s = 228;
	{8'd132,8'd70} : s = 226;
	{8'd132,8'd71} : s = 370;
	{8'd132,8'd72} : s = 225;
	{8'd132,8'd73} : s = 369;
	{8'd132,8'd74} : s = 364;
	{8'd132,8'd75} : s = 470;
	{8'd132,8'd76} : s = 88;
	{8'd132,8'd77} : s = 216;
	{8'd132,8'd78} : s = 212;
	{8'd132,8'd79} : s = 362;
	{8'd132,8'd80} : s = 210;
	{8'd132,8'd81} : s = 361;
	{8'd132,8'd82} : s = 358;
	{8'd132,8'd83} : s = 469;
	{8'd132,8'd84} : s = 209;
	{8'd132,8'd85} : s = 357;
	{8'd132,8'd86} : s = 355;
	{8'd132,8'd87} : s = 467;
	{8'd132,8'd88} : s = 348;
	{8'd132,8'd89} : s = 462;
	{8'd132,8'd90} : s = 461;
	{8'd132,8'd91} : s = 505;
	{8'd132,8'd92} : s = 84;
	{8'd132,8'd93} : s = 204;
	{8'd132,8'd94} : s = 202;
	{8'd132,8'd95} : s = 346;
	{8'd132,8'd96} : s = 201;
	{8'd132,8'd97} : s = 345;
	{8'd132,8'd98} : s = 342;
	{8'd132,8'd99} : s = 459;
	{8'd132,8'd100} : s = 198;
	{8'd132,8'd101} : s = 341;
	{8'd132,8'd102} : s = 339;
	{8'd132,8'd103} : s = 455;
	{8'd132,8'd104} : s = 334;
	{8'd132,8'd105} : s = 444;
	{8'd132,8'd106} : s = 442;
	{8'd132,8'd107} : s = 502;
	{8'd132,8'd108} : s = 197;
	{8'd132,8'd109} : s = 333;
	{8'd132,8'd110} : s = 331;
	{8'd132,8'd111} : s = 441;
	{8'd132,8'd112} : s = 327;
	{8'd132,8'd113} : s = 438;
	{8'd132,8'd114} : s = 437;
	{8'd132,8'd115} : s = 501;
	{8'd132,8'd116} : s = 316;
	{8'd132,8'd117} : s = 435;
	{8'd132,8'd118} : s = 430;
	{8'd132,8'd119} : s = 499;
	{8'd132,8'd120} : s = 429;
	{8'd132,8'd121} : s = 494;
	{8'd132,8'd122} : s = 493;
	{8'd132,8'd123} : s = 510;
	{8'd132,8'd124} : s = 1;
	{8'd132,8'd125} : s = 18;
	{8'd132,8'd126} : s = 17;
	{8'd132,8'd127} : s = 82;
	{8'd132,8'd128} : s = 12;
	{8'd132,8'd129} : s = 81;
	{8'd132,8'd130} : s = 76;
	{8'd132,8'd131} : s = 195;
	{8'd132,8'd132} : s = 10;
	{8'd132,8'd133} : s = 74;
	{8'd132,8'd134} : s = 73;
	{8'd132,8'd135} : s = 184;
	{8'd132,8'd136} : s = 70;
	{8'd132,8'd137} : s = 180;
	{8'd132,8'd138} : s = 178;
	{8'd132,8'd139} : s = 314;
	{8'd132,8'd140} : s = 9;
	{8'd132,8'd141} : s = 69;
	{8'd132,8'd142} : s = 67;
	{8'd132,8'd143} : s = 177;
	{8'd132,8'd144} : s = 56;
	{8'd132,8'd145} : s = 172;
	{8'd132,8'd146} : s = 170;
	{8'd132,8'd147} : s = 313;
	{8'd132,8'd148} : s = 52;
	{8'd132,8'd149} : s = 169;
	{8'd132,8'd150} : s = 166;
	{8'd132,8'd151} : s = 310;
	{8'd132,8'd152} : s = 165;
	{8'd132,8'd153} : s = 309;
	{8'd132,8'd154} : s = 307;
	{8'd132,8'd155} : s = 427;
	{8'd132,8'd156} : s = 6;
	{8'd132,8'd157} : s = 50;
	{8'd132,8'd158} : s = 49;
	{8'd132,8'd159} : s = 163;
	{8'd132,8'd160} : s = 44;
	{8'd132,8'd161} : s = 156;
	{8'd132,8'd162} : s = 154;
	{8'd132,8'd163} : s = 302;
	{8'd132,8'd164} : s = 42;
	{8'd132,8'd165} : s = 153;
	{8'd132,8'd166} : s = 150;
	{8'd132,8'd167} : s = 301;
	{8'd132,8'd168} : s = 149;
	{8'd132,8'd169} : s = 299;
	{8'd132,8'd170} : s = 295;
	{8'd132,8'd171} : s = 423;
	{8'd132,8'd172} : s = 41;
	{8'd132,8'd173} : s = 147;
	{8'd132,8'd174} : s = 142;
	{8'd132,8'd175} : s = 286;
	{8'd132,8'd176} : s = 141;
	{8'd132,8'd177} : s = 285;
	{8'd132,8'd178} : s = 283;
	{8'd132,8'd179} : s = 414;
	{8'd132,8'd180} : s = 139;
	{8'd132,8'd181} : s = 279;
	{8'd132,8'd182} : s = 271;
	{8'd132,8'd183} : s = 413;
	{8'd132,8'd184} : s = 248;
	{8'd132,8'd185} : s = 411;
	{8'd132,8'd186} : s = 407;
	{8'd132,8'd187} : s = 491;
	{8'd132,8'd188} : s = 5;
	{8'd132,8'd189} : s = 38;
	{8'd132,8'd190} : s = 37;
	{8'd132,8'd191} : s = 135;
	{8'd132,8'd192} : s = 35;
	{8'd132,8'd193} : s = 120;
	{8'd132,8'd194} : s = 116;
	{8'd132,8'd195} : s = 244;
	{8'd132,8'd196} : s = 28;
	{8'd132,8'd197} : s = 114;
	{8'd132,8'd198} : s = 113;
	{8'd132,8'd199} : s = 242;
	{8'd132,8'd200} : s = 108;
	{8'd132,8'd201} : s = 241;
	{8'd132,8'd202} : s = 236;
	{8'd132,8'd203} : s = 399;
	{8'd132,8'd204} : s = 26;
	{8'd132,8'd205} : s = 106;
	{8'd132,8'd206} : s = 105;
	{8'd132,8'd207} : s = 234;
	{8'd132,8'd208} : s = 102;
	{8'd132,8'd209} : s = 233;
	{8'd132,8'd210} : s = 230;
	{8'd132,8'd211} : s = 380;
	{8'd132,8'd212} : s = 101;
	{8'd132,8'd213} : s = 229;
	{8'd132,8'd214} : s = 227;
	{8'd132,8'd215} : s = 378;
	{8'd132,8'd216} : s = 220;
	{8'd132,8'd217} : s = 377;
	{8'd132,8'd218} : s = 374;
	{8'd132,8'd219} : s = 487;
	{8'd132,8'd220} : s = 25;
	{8'd132,8'd221} : s = 99;
	{8'd132,8'd222} : s = 92;
	{8'd132,8'd223} : s = 218;
	{8'd132,8'd224} : s = 90;
	{8'd132,8'd225} : s = 217;
	{8'd132,8'd226} : s = 214;
	{8'd132,8'd227} : s = 373;
	{8'd132,8'd228} : s = 89;
	{8'd132,8'd229} : s = 213;
	{8'd132,8'd230} : s = 211;
	{8'd132,8'd231} : s = 371;
	{8'd132,8'd232} : s = 206;
	{8'd132,8'd233} : s = 366;
	{8'd132,8'd234} : s = 365;
	{8'd132,8'd235} : s = 478;
	{8'd132,8'd236} : s = 86;
	{8'd132,8'd237} : s = 205;
	{8'd132,8'd238} : s = 203;
	{8'd132,8'd239} : s = 363;
	{8'd132,8'd240} : s = 199;
	{8'd132,8'd241} : s = 359;
	{8'd132,8'd242} : s = 350;
	{8'd132,8'd243} : s = 477;
	{8'd132,8'd244} : s = 188;
	{8'd132,8'd245} : s = 349;
	{8'd132,8'd246} : s = 347;
	{8'd132,8'd247} : s = 475;
	{8'd132,8'd248} : s = 343;
	{8'd132,8'd249} : s = 471;
	{8'd132,8'd250} : s = 463;
	{8'd132,8'd251} : s = 509;
	{8'd132,8'd252} : s = 3;
	{8'd132,8'd253} : s = 22;
	{8'd132,8'd254} : s = 21;
	{8'd132,8'd255} : s = 85;
	{8'd133,8'd0} : s = 164;
	{8'd133,8'd1} : s = 162;
	{8'd133,8'd2} : s = 323;
	{8'd133,8'd3} : s = 34;
	{8'd133,8'd4} : s = 161;
	{8'd133,8'd5} : s = 152;
	{8'd133,8'd6} : s = 312;
	{8'd133,8'd7} : s = 148;
	{8'd133,8'd8} : s = 308;
	{8'd133,8'd9} : s = 306;
	{8'd133,8'd10} : s = 425;
	{8'd133,8'd11} : s = 33;
	{8'd133,8'd12} : s = 146;
	{8'd133,8'd13} : s = 145;
	{8'd133,8'd14} : s = 305;
	{8'd133,8'd15} : s = 140;
	{8'd133,8'd16} : s = 300;
	{8'd133,8'd17} : s = 298;
	{8'd133,8'd18} : s = 422;
	{8'd133,8'd19} : s = 138;
	{8'd133,8'd20} : s = 297;
	{8'd133,8'd21} : s = 294;
	{8'd133,8'd22} : s = 421;
	{8'd133,8'd23} : s = 293;
	{8'd133,8'd24} : s = 419;
	{8'd133,8'd25} : s = 412;
	{8'd133,8'd26} : s = 486;
	{8'd133,8'd27} : s = 24;
	{8'd133,8'd28} : s = 137;
	{8'd133,8'd29} : s = 134;
	{8'd133,8'd30} : s = 291;
	{8'd133,8'd31} : s = 133;
	{8'd133,8'd32} : s = 284;
	{8'd133,8'd33} : s = 282;
	{8'd133,8'd34} : s = 410;
	{8'd133,8'd35} : s = 131;
	{8'd133,8'd36} : s = 281;
	{8'd133,8'd37} : s = 278;
	{8'd133,8'd38} : s = 409;
	{8'd133,8'd39} : s = 277;
	{8'd133,8'd40} : s = 406;
	{8'd133,8'd41} : s = 405;
	{8'd133,8'd42} : s = 485;
	{8'd133,8'd43} : s = 112;
	{8'd133,8'd44} : s = 275;
	{8'd133,8'd45} : s = 270;
	{8'd133,8'd46} : s = 403;
	{8'd133,8'd47} : s = 269;
	{8'd133,8'd48} : s = 398;
	{8'd133,8'd49} : s = 397;
	{8'd133,8'd50} : s = 483;
	{8'd133,8'd51} : s = 267;
	{8'd133,8'd52} : s = 395;
	{8'd133,8'd53} : s = 391;
	{8'd133,8'd54} : s = 476;
	{8'd133,8'd55} : s = 376;
	{8'd133,8'd56} : s = 474;
	{8'd133,8'd57} : s = 473;
	{8'd133,8'd58} : s = 506;
	{8'd133,8'd59} : s = 20;
	{8'd133,8'd60} : s = 104;
	{8'd133,8'd61} : s = 100;
	{8'd133,8'd62} : s = 263;
	{8'd133,8'd63} : s = 98;
	{8'd133,8'd64} : s = 240;
	{8'd133,8'd65} : s = 232;
	{8'd133,8'd66} : s = 372;
	{8'd133,8'd67} : s = 97;
	{8'd133,8'd68} : s = 228;
	{8'd133,8'd69} : s = 226;
	{8'd133,8'd70} : s = 370;
	{8'd133,8'd71} : s = 225;
	{8'd133,8'd72} : s = 369;
	{8'd133,8'd73} : s = 364;
	{8'd133,8'd74} : s = 470;
	{8'd133,8'd75} : s = 88;
	{8'd133,8'd76} : s = 216;
	{8'd133,8'd77} : s = 212;
	{8'd133,8'd78} : s = 362;
	{8'd133,8'd79} : s = 210;
	{8'd133,8'd80} : s = 361;
	{8'd133,8'd81} : s = 358;
	{8'd133,8'd82} : s = 469;
	{8'd133,8'd83} : s = 209;
	{8'd133,8'd84} : s = 357;
	{8'd133,8'd85} : s = 355;
	{8'd133,8'd86} : s = 467;
	{8'd133,8'd87} : s = 348;
	{8'd133,8'd88} : s = 462;
	{8'd133,8'd89} : s = 461;
	{8'd133,8'd90} : s = 505;
	{8'd133,8'd91} : s = 84;
	{8'd133,8'd92} : s = 204;
	{8'd133,8'd93} : s = 202;
	{8'd133,8'd94} : s = 346;
	{8'd133,8'd95} : s = 201;
	{8'd133,8'd96} : s = 345;
	{8'd133,8'd97} : s = 342;
	{8'd133,8'd98} : s = 459;
	{8'd133,8'd99} : s = 198;
	{8'd133,8'd100} : s = 341;
	{8'd133,8'd101} : s = 339;
	{8'd133,8'd102} : s = 455;
	{8'd133,8'd103} : s = 334;
	{8'd133,8'd104} : s = 444;
	{8'd133,8'd105} : s = 442;
	{8'd133,8'd106} : s = 502;
	{8'd133,8'd107} : s = 197;
	{8'd133,8'd108} : s = 333;
	{8'd133,8'd109} : s = 331;
	{8'd133,8'd110} : s = 441;
	{8'd133,8'd111} : s = 327;
	{8'd133,8'd112} : s = 438;
	{8'd133,8'd113} : s = 437;
	{8'd133,8'd114} : s = 501;
	{8'd133,8'd115} : s = 316;
	{8'd133,8'd116} : s = 435;
	{8'd133,8'd117} : s = 430;
	{8'd133,8'd118} : s = 499;
	{8'd133,8'd119} : s = 429;
	{8'd133,8'd120} : s = 494;
	{8'd133,8'd121} : s = 493;
	{8'd133,8'd122} : s = 510;
	{8'd133,8'd123} : s = 1;
	{8'd133,8'd124} : s = 18;
	{8'd133,8'd125} : s = 17;
	{8'd133,8'd126} : s = 82;
	{8'd133,8'd127} : s = 12;
	{8'd133,8'd128} : s = 81;
	{8'd133,8'd129} : s = 76;
	{8'd133,8'd130} : s = 195;
	{8'd133,8'd131} : s = 10;
	{8'd133,8'd132} : s = 74;
	{8'd133,8'd133} : s = 73;
	{8'd133,8'd134} : s = 184;
	{8'd133,8'd135} : s = 70;
	{8'd133,8'd136} : s = 180;
	{8'd133,8'd137} : s = 178;
	{8'd133,8'd138} : s = 314;
	{8'd133,8'd139} : s = 9;
	{8'd133,8'd140} : s = 69;
	{8'd133,8'd141} : s = 67;
	{8'd133,8'd142} : s = 177;
	{8'd133,8'd143} : s = 56;
	{8'd133,8'd144} : s = 172;
	{8'd133,8'd145} : s = 170;
	{8'd133,8'd146} : s = 313;
	{8'd133,8'd147} : s = 52;
	{8'd133,8'd148} : s = 169;
	{8'd133,8'd149} : s = 166;
	{8'd133,8'd150} : s = 310;
	{8'd133,8'd151} : s = 165;
	{8'd133,8'd152} : s = 309;
	{8'd133,8'd153} : s = 307;
	{8'd133,8'd154} : s = 427;
	{8'd133,8'd155} : s = 6;
	{8'd133,8'd156} : s = 50;
	{8'd133,8'd157} : s = 49;
	{8'd133,8'd158} : s = 163;
	{8'd133,8'd159} : s = 44;
	{8'd133,8'd160} : s = 156;
	{8'd133,8'd161} : s = 154;
	{8'd133,8'd162} : s = 302;
	{8'd133,8'd163} : s = 42;
	{8'd133,8'd164} : s = 153;
	{8'd133,8'd165} : s = 150;
	{8'd133,8'd166} : s = 301;
	{8'd133,8'd167} : s = 149;
	{8'd133,8'd168} : s = 299;
	{8'd133,8'd169} : s = 295;
	{8'd133,8'd170} : s = 423;
	{8'd133,8'd171} : s = 41;
	{8'd133,8'd172} : s = 147;
	{8'd133,8'd173} : s = 142;
	{8'd133,8'd174} : s = 286;
	{8'd133,8'd175} : s = 141;
	{8'd133,8'd176} : s = 285;
	{8'd133,8'd177} : s = 283;
	{8'd133,8'd178} : s = 414;
	{8'd133,8'd179} : s = 139;
	{8'd133,8'd180} : s = 279;
	{8'd133,8'd181} : s = 271;
	{8'd133,8'd182} : s = 413;
	{8'd133,8'd183} : s = 248;
	{8'd133,8'd184} : s = 411;
	{8'd133,8'd185} : s = 407;
	{8'd133,8'd186} : s = 491;
	{8'd133,8'd187} : s = 5;
	{8'd133,8'd188} : s = 38;
	{8'd133,8'd189} : s = 37;
	{8'd133,8'd190} : s = 135;
	{8'd133,8'd191} : s = 35;
	{8'd133,8'd192} : s = 120;
	{8'd133,8'd193} : s = 116;
	{8'd133,8'd194} : s = 244;
	{8'd133,8'd195} : s = 28;
	{8'd133,8'd196} : s = 114;
	{8'd133,8'd197} : s = 113;
	{8'd133,8'd198} : s = 242;
	{8'd133,8'd199} : s = 108;
	{8'd133,8'd200} : s = 241;
	{8'd133,8'd201} : s = 236;
	{8'd133,8'd202} : s = 399;
	{8'd133,8'd203} : s = 26;
	{8'd133,8'd204} : s = 106;
	{8'd133,8'd205} : s = 105;
	{8'd133,8'd206} : s = 234;
	{8'd133,8'd207} : s = 102;
	{8'd133,8'd208} : s = 233;
	{8'd133,8'd209} : s = 230;
	{8'd133,8'd210} : s = 380;
	{8'd133,8'd211} : s = 101;
	{8'd133,8'd212} : s = 229;
	{8'd133,8'd213} : s = 227;
	{8'd133,8'd214} : s = 378;
	{8'd133,8'd215} : s = 220;
	{8'd133,8'd216} : s = 377;
	{8'd133,8'd217} : s = 374;
	{8'd133,8'd218} : s = 487;
	{8'd133,8'd219} : s = 25;
	{8'd133,8'd220} : s = 99;
	{8'd133,8'd221} : s = 92;
	{8'd133,8'd222} : s = 218;
	{8'd133,8'd223} : s = 90;
	{8'd133,8'd224} : s = 217;
	{8'd133,8'd225} : s = 214;
	{8'd133,8'd226} : s = 373;
	{8'd133,8'd227} : s = 89;
	{8'd133,8'd228} : s = 213;
	{8'd133,8'd229} : s = 211;
	{8'd133,8'd230} : s = 371;
	{8'd133,8'd231} : s = 206;
	{8'd133,8'd232} : s = 366;
	{8'd133,8'd233} : s = 365;
	{8'd133,8'd234} : s = 478;
	{8'd133,8'd235} : s = 86;
	{8'd133,8'd236} : s = 205;
	{8'd133,8'd237} : s = 203;
	{8'd133,8'd238} : s = 363;
	{8'd133,8'd239} : s = 199;
	{8'd133,8'd240} : s = 359;
	{8'd133,8'd241} : s = 350;
	{8'd133,8'd242} : s = 477;
	{8'd133,8'd243} : s = 188;
	{8'd133,8'd244} : s = 349;
	{8'd133,8'd245} : s = 347;
	{8'd133,8'd246} : s = 475;
	{8'd133,8'd247} : s = 343;
	{8'd133,8'd248} : s = 471;
	{8'd133,8'd249} : s = 463;
	{8'd133,8'd250} : s = 509;
	{8'd133,8'd251} : s = 3;
	{8'd133,8'd252} : s = 22;
	{8'd133,8'd253} : s = 21;
	{8'd133,8'd254} : s = 85;
	{8'd133,8'd255} : s = 19;
	{8'd134,8'd0} : s = 162;
	{8'd134,8'd1} : s = 323;
	{8'd134,8'd2} : s = 34;
	{8'd134,8'd3} : s = 161;
	{8'd134,8'd4} : s = 152;
	{8'd134,8'd5} : s = 312;
	{8'd134,8'd6} : s = 148;
	{8'd134,8'd7} : s = 308;
	{8'd134,8'd8} : s = 306;
	{8'd134,8'd9} : s = 425;
	{8'd134,8'd10} : s = 33;
	{8'd134,8'd11} : s = 146;
	{8'd134,8'd12} : s = 145;
	{8'd134,8'd13} : s = 305;
	{8'd134,8'd14} : s = 140;
	{8'd134,8'd15} : s = 300;
	{8'd134,8'd16} : s = 298;
	{8'd134,8'd17} : s = 422;
	{8'd134,8'd18} : s = 138;
	{8'd134,8'd19} : s = 297;
	{8'd134,8'd20} : s = 294;
	{8'd134,8'd21} : s = 421;
	{8'd134,8'd22} : s = 293;
	{8'd134,8'd23} : s = 419;
	{8'd134,8'd24} : s = 412;
	{8'd134,8'd25} : s = 486;
	{8'd134,8'd26} : s = 24;
	{8'd134,8'd27} : s = 137;
	{8'd134,8'd28} : s = 134;
	{8'd134,8'd29} : s = 291;
	{8'd134,8'd30} : s = 133;
	{8'd134,8'd31} : s = 284;
	{8'd134,8'd32} : s = 282;
	{8'd134,8'd33} : s = 410;
	{8'd134,8'd34} : s = 131;
	{8'd134,8'd35} : s = 281;
	{8'd134,8'd36} : s = 278;
	{8'd134,8'd37} : s = 409;
	{8'd134,8'd38} : s = 277;
	{8'd134,8'd39} : s = 406;
	{8'd134,8'd40} : s = 405;
	{8'd134,8'd41} : s = 485;
	{8'd134,8'd42} : s = 112;
	{8'd134,8'd43} : s = 275;
	{8'd134,8'd44} : s = 270;
	{8'd134,8'd45} : s = 403;
	{8'd134,8'd46} : s = 269;
	{8'd134,8'd47} : s = 398;
	{8'd134,8'd48} : s = 397;
	{8'd134,8'd49} : s = 483;
	{8'd134,8'd50} : s = 267;
	{8'd134,8'd51} : s = 395;
	{8'd134,8'd52} : s = 391;
	{8'd134,8'd53} : s = 476;
	{8'd134,8'd54} : s = 376;
	{8'd134,8'd55} : s = 474;
	{8'd134,8'd56} : s = 473;
	{8'd134,8'd57} : s = 506;
	{8'd134,8'd58} : s = 20;
	{8'd134,8'd59} : s = 104;
	{8'd134,8'd60} : s = 100;
	{8'd134,8'd61} : s = 263;
	{8'd134,8'd62} : s = 98;
	{8'd134,8'd63} : s = 240;
	{8'd134,8'd64} : s = 232;
	{8'd134,8'd65} : s = 372;
	{8'd134,8'd66} : s = 97;
	{8'd134,8'd67} : s = 228;
	{8'd134,8'd68} : s = 226;
	{8'd134,8'd69} : s = 370;
	{8'd134,8'd70} : s = 225;
	{8'd134,8'd71} : s = 369;
	{8'd134,8'd72} : s = 364;
	{8'd134,8'd73} : s = 470;
	{8'd134,8'd74} : s = 88;
	{8'd134,8'd75} : s = 216;
	{8'd134,8'd76} : s = 212;
	{8'd134,8'd77} : s = 362;
	{8'd134,8'd78} : s = 210;
	{8'd134,8'd79} : s = 361;
	{8'd134,8'd80} : s = 358;
	{8'd134,8'd81} : s = 469;
	{8'd134,8'd82} : s = 209;
	{8'd134,8'd83} : s = 357;
	{8'd134,8'd84} : s = 355;
	{8'd134,8'd85} : s = 467;
	{8'd134,8'd86} : s = 348;
	{8'd134,8'd87} : s = 462;
	{8'd134,8'd88} : s = 461;
	{8'd134,8'd89} : s = 505;
	{8'd134,8'd90} : s = 84;
	{8'd134,8'd91} : s = 204;
	{8'd134,8'd92} : s = 202;
	{8'd134,8'd93} : s = 346;
	{8'd134,8'd94} : s = 201;
	{8'd134,8'd95} : s = 345;
	{8'd134,8'd96} : s = 342;
	{8'd134,8'd97} : s = 459;
	{8'd134,8'd98} : s = 198;
	{8'd134,8'd99} : s = 341;
	{8'd134,8'd100} : s = 339;
	{8'd134,8'd101} : s = 455;
	{8'd134,8'd102} : s = 334;
	{8'd134,8'd103} : s = 444;
	{8'd134,8'd104} : s = 442;
	{8'd134,8'd105} : s = 502;
	{8'd134,8'd106} : s = 197;
	{8'd134,8'd107} : s = 333;
	{8'd134,8'd108} : s = 331;
	{8'd134,8'd109} : s = 441;
	{8'd134,8'd110} : s = 327;
	{8'd134,8'd111} : s = 438;
	{8'd134,8'd112} : s = 437;
	{8'd134,8'd113} : s = 501;
	{8'd134,8'd114} : s = 316;
	{8'd134,8'd115} : s = 435;
	{8'd134,8'd116} : s = 430;
	{8'd134,8'd117} : s = 499;
	{8'd134,8'd118} : s = 429;
	{8'd134,8'd119} : s = 494;
	{8'd134,8'd120} : s = 493;
	{8'd134,8'd121} : s = 510;
	{8'd134,8'd122} : s = 1;
	{8'd134,8'd123} : s = 18;
	{8'd134,8'd124} : s = 17;
	{8'd134,8'd125} : s = 82;
	{8'd134,8'd126} : s = 12;
	{8'd134,8'd127} : s = 81;
	{8'd134,8'd128} : s = 76;
	{8'd134,8'd129} : s = 195;
	{8'd134,8'd130} : s = 10;
	{8'd134,8'd131} : s = 74;
	{8'd134,8'd132} : s = 73;
	{8'd134,8'd133} : s = 184;
	{8'd134,8'd134} : s = 70;
	{8'd134,8'd135} : s = 180;
	{8'd134,8'd136} : s = 178;
	{8'd134,8'd137} : s = 314;
	{8'd134,8'd138} : s = 9;
	{8'd134,8'd139} : s = 69;
	{8'd134,8'd140} : s = 67;
	{8'd134,8'd141} : s = 177;
	{8'd134,8'd142} : s = 56;
	{8'd134,8'd143} : s = 172;
	{8'd134,8'd144} : s = 170;
	{8'd134,8'd145} : s = 313;
	{8'd134,8'd146} : s = 52;
	{8'd134,8'd147} : s = 169;
	{8'd134,8'd148} : s = 166;
	{8'd134,8'd149} : s = 310;
	{8'd134,8'd150} : s = 165;
	{8'd134,8'd151} : s = 309;
	{8'd134,8'd152} : s = 307;
	{8'd134,8'd153} : s = 427;
	{8'd134,8'd154} : s = 6;
	{8'd134,8'd155} : s = 50;
	{8'd134,8'd156} : s = 49;
	{8'd134,8'd157} : s = 163;
	{8'd134,8'd158} : s = 44;
	{8'd134,8'd159} : s = 156;
	{8'd134,8'd160} : s = 154;
	{8'd134,8'd161} : s = 302;
	{8'd134,8'd162} : s = 42;
	{8'd134,8'd163} : s = 153;
	{8'd134,8'd164} : s = 150;
	{8'd134,8'd165} : s = 301;
	{8'd134,8'd166} : s = 149;
	{8'd134,8'd167} : s = 299;
	{8'd134,8'd168} : s = 295;
	{8'd134,8'd169} : s = 423;
	{8'd134,8'd170} : s = 41;
	{8'd134,8'd171} : s = 147;
	{8'd134,8'd172} : s = 142;
	{8'd134,8'd173} : s = 286;
	{8'd134,8'd174} : s = 141;
	{8'd134,8'd175} : s = 285;
	{8'd134,8'd176} : s = 283;
	{8'd134,8'd177} : s = 414;
	{8'd134,8'd178} : s = 139;
	{8'd134,8'd179} : s = 279;
	{8'd134,8'd180} : s = 271;
	{8'd134,8'd181} : s = 413;
	{8'd134,8'd182} : s = 248;
	{8'd134,8'd183} : s = 411;
	{8'd134,8'd184} : s = 407;
	{8'd134,8'd185} : s = 491;
	{8'd134,8'd186} : s = 5;
	{8'd134,8'd187} : s = 38;
	{8'd134,8'd188} : s = 37;
	{8'd134,8'd189} : s = 135;
	{8'd134,8'd190} : s = 35;
	{8'd134,8'd191} : s = 120;
	{8'd134,8'd192} : s = 116;
	{8'd134,8'd193} : s = 244;
	{8'd134,8'd194} : s = 28;
	{8'd134,8'd195} : s = 114;
	{8'd134,8'd196} : s = 113;
	{8'd134,8'd197} : s = 242;
	{8'd134,8'd198} : s = 108;
	{8'd134,8'd199} : s = 241;
	{8'd134,8'd200} : s = 236;
	{8'd134,8'd201} : s = 399;
	{8'd134,8'd202} : s = 26;
	{8'd134,8'd203} : s = 106;
	{8'd134,8'd204} : s = 105;
	{8'd134,8'd205} : s = 234;
	{8'd134,8'd206} : s = 102;
	{8'd134,8'd207} : s = 233;
	{8'd134,8'd208} : s = 230;
	{8'd134,8'd209} : s = 380;
	{8'd134,8'd210} : s = 101;
	{8'd134,8'd211} : s = 229;
	{8'd134,8'd212} : s = 227;
	{8'd134,8'd213} : s = 378;
	{8'd134,8'd214} : s = 220;
	{8'd134,8'd215} : s = 377;
	{8'd134,8'd216} : s = 374;
	{8'd134,8'd217} : s = 487;
	{8'd134,8'd218} : s = 25;
	{8'd134,8'd219} : s = 99;
	{8'd134,8'd220} : s = 92;
	{8'd134,8'd221} : s = 218;
	{8'd134,8'd222} : s = 90;
	{8'd134,8'd223} : s = 217;
	{8'd134,8'd224} : s = 214;
	{8'd134,8'd225} : s = 373;
	{8'd134,8'd226} : s = 89;
	{8'd134,8'd227} : s = 213;
	{8'd134,8'd228} : s = 211;
	{8'd134,8'd229} : s = 371;
	{8'd134,8'd230} : s = 206;
	{8'd134,8'd231} : s = 366;
	{8'd134,8'd232} : s = 365;
	{8'd134,8'd233} : s = 478;
	{8'd134,8'd234} : s = 86;
	{8'd134,8'd235} : s = 205;
	{8'd134,8'd236} : s = 203;
	{8'd134,8'd237} : s = 363;
	{8'd134,8'd238} : s = 199;
	{8'd134,8'd239} : s = 359;
	{8'd134,8'd240} : s = 350;
	{8'd134,8'd241} : s = 477;
	{8'd134,8'd242} : s = 188;
	{8'd134,8'd243} : s = 349;
	{8'd134,8'd244} : s = 347;
	{8'd134,8'd245} : s = 475;
	{8'd134,8'd246} : s = 343;
	{8'd134,8'd247} : s = 471;
	{8'd134,8'd248} : s = 463;
	{8'd134,8'd249} : s = 509;
	{8'd134,8'd250} : s = 3;
	{8'd134,8'd251} : s = 22;
	{8'd134,8'd252} : s = 21;
	{8'd134,8'd253} : s = 85;
	{8'd134,8'd254} : s = 19;
	{8'd134,8'd255} : s = 83;
	{8'd135,8'd0} : s = 323;
	{8'd135,8'd1} : s = 34;
	{8'd135,8'd2} : s = 161;
	{8'd135,8'd3} : s = 152;
	{8'd135,8'd4} : s = 312;
	{8'd135,8'd5} : s = 148;
	{8'd135,8'd6} : s = 308;
	{8'd135,8'd7} : s = 306;
	{8'd135,8'd8} : s = 425;
	{8'd135,8'd9} : s = 33;
	{8'd135,8'd10} : s = 146;
	{8'd135,8'd11} : s = 145;
	{8'd135,8'd12} : s = 305;
	{8'd135,8'd13} : s = 140;
	{8'd135,8'd14} : s = 300;
	{8'd135,8'd15} : s = 298;
	{8'd135,8'd16} : s = 422;
	{8'd135,8'd17} : s = 138;
	{8'd135,8'd18} : s = 297;
	{8'd135,8'd19} : s = 294;
	{8'd135,8'd20} : s = 421;
	{8'd135,8'd21} : s = 293;
	{8'd135,8'd22} : s = 419;
	{8'd135,8'd23} : s = 412;
	{8'd135,8'd24} : s = 486;
	{8'd135,8'd25} : s = 24;
	{8'd135,8'd26} : s = 137;
	{8'd135,8'd27} : s = 134;
	{8'd135,8'd28} : s = 291;
	{8'd135,8'd29} : s = 133;
	{8'd135,8'd30} : s = 284;
	{8'd135,8'd31} : s = 282;
	{8'd135,8'd32} : s = 410;
	{8'd135,8'd33} : s = 131;
	{8'd135,8'd34} : s = 281;
	{8'd135,8'd35} : s = 278;
	{8'd135,8'd36} : s = 409;
	{8'd135,8'd37} : s = 277;
	{8'd135,8'd38} : s = 406;
	{8'd135,8'd39} : s = 405;
	{8'd135,8'd40} : s = 485;
	{8'd135,8'd41} : s = 112;
	{8'd135,8'd42} : s = 275;
	{8'd135,8'd43} : s = 270;
	{8'd135,8'd44} : s = 403;
	{8'd135,8'd45} : s = 269;
	{8'd135,8'd46} : s = 398;
	{8'd135,8'd47} : s = 397;
	{8'd135,8'd48} : s = 483;
	{8'd135,8'd49} : s = 267;
	{8'd135,8'd50} : s = 395;
	{8'd135,8'd51} : s = 391;
	{8'd135,8'd52} : s = 476;
	{8'd135,8'd53} : s = 376;
	{8'd135,8'd54} : s = 474;
	{8'd135,8'd55} : s = 473;
	{8'd135,8'd56} : s = 506;
	{8'd135,8'd57} : s = 20;
	{8'd135,8'd58} : s = 104;
	{8'd135,8'd59} : s = 100;
	{8'd135,8'd60} : s = 263;
	{8'd135,8'd61} : s = 98;
	{8'd135,8'd62} : s = 240;
	{8'd135,8'd63} : s = 232;
	{8'd135,8'd64} : s = 372;
	{8'd135,8'd65} : s = 97;
	{8'd135,8'd66} : s = 228;
	{8'd135,8'd67} : s = 226;
	{8'd135,8'd68} : s = 370;
	{8'd135,8'd69} : s = 225;
	{8'd135,8'd70} : s = 369;
	{8'd135,8'd71} : s = 364;
	{8'd135,8'd72} : s = 470;
	{8'd135,8'd73} : s = 88;
	{8'd135,8'd74} : s = 216;
	{8'd135,8'd75} : s = 212;
	{8'd135,8'd76} : s = 362;
	{8'd135,8'd77} : s = 210;
	{8'd135,8'd78} : s = 361;
	{8'd135,8'd79} : s = 358;
	{8'd135,8'd80} : s = 469;
	{8'd135,8'd81} : s = 209;
	{8'd135,8'd82} : s = 357;
	{8'd135,8'd83} : s = 355;
	{8'd135,8'd84} : s = 467;
	{8'd135,8'd85} : s = 348;
	{8'd135,8'd86} : s = 462;
	{8'd135,8'd87} : s = 461;
	{8'd135,8'd88} : s = 505;
	{8'd135,8'd89} : s = 84;
	{8'd135,8'd90} : s = 204;
	{8'd135,8'd91} : s = 202;
	{8'd135,8'd92} : s = 346;
	{8'd135,8'd93} : s = 201;
	{8'd135,8'd94} : s = 345;
	{8'd135,8'd95} : s = 342;
	{8'd135,8'd96} : s = 459;
	{8'd135,8'd97} : s = 198;
	{8'd135,8'd98} : s = 341;
	{8'd135,8'd99} : s = 339;
	{8'd135,8'd100} : s = 455;
	{8'd135,8'd101} : s = 334;
	{8'd135,8'd102} : s = 444;
	{8'd135,8'd103} : s = 442;
	{8'd135,8'd104} : s = 502;
	{8'd135,8'd105} : s = 197;
	{8'd135,8'd106} : s = 333;
	{8'd135,8'd107} : s = 331;
	{8'd135,8'd108} : s = 441;
	{8'd135,8'd109} : s = 327;
	{8'd135,8'd110} : s = 438;
	{8'd135,8'd111} : s = 437;
	{8'd135,8'd112} : s = 501;
	{8'd135,8'd113} : s = 316;
	{8'd135,8'd114} : s = 435;
	{8'd135,8'd115} : s = 430;
	{8'd135,8'd116} : s = 499;
	{8'd135,8'd117} : s = 429;
	{8'd135,8'd118} : s = 494;
	{8'd135,8'd119} : s = 493;
	{8'd135,8'd120} : s = 510;
	{8'd135,8'd121} : s = 1;
	{8'd135,8'd122} : s = 18;
	{8'd135,8'd123} : s = 17;
	{8'd135,8'd124} : s = 82;
	{8'd135,8'd125} : s = 12;
	{8'd135,8'd126} : s = 81;
	{8'd135,8'd127} : s = 76;
	{8'd135,8'd128} : s = 195;
	{8'd135,8'd129} : s = 10;
	{8'd135,8'd130} : s = 74;
	{8'd135,8'd131} : s = 73;
	{8'd135,8'd132} : s = 184;
	{8'd135,8'd133} : s = 70;
	{8'd135,8'd134} : s = 180;
	{8'd135,8'd135} : s = 178;
	{8'd135,8'd136} : s = 314;
	{8'd135,8'd137} : s = 9;
	{8'd135,8'd138} : s = 69;
	{8'd135,8'd139} : s = 67;
	{8'd135,8'd140} : s = 177;
	{8'd135,8'd141} : s = 56;
	{8'd135,8'd142} : s = 172;
	{8'd135,8'd143} : s = 170;
	{8'd135,8'd144} : s = 313;
	{8'd135,8'd145} : s = 52;
	{8'd135,8'd146} : s = 169;
	{8'd135,8'd147} : s = 166;
	{8'd135,8'd148} : s = 310;
	{8'd135,8'd149} : s = 165;
	{8'd135,8'd150} : s = 309;
	{8'd135,8'd151} : s = 307;
	{8'd135,8'd152} : s = 427;
	{8'd135,8'd153} : s = 6;
	{8'd135,8'd154} : s = 50;
	{8'd135,8'd155} : s = 49;
	{8'd135,8'd156} : s = 163;
	{8'd135,8'd157} : s = 44;
	{8'd135,8'd158} : s = 156;
	{8'd135,8'd159} : s = 154;
	{8'd135,8'd160} : s = 302;
	{8'd135,8'd161} : s = 42;
	{8'd135,8'd162} : s = 153;
	{8'd135,8'd163} : s = 150;
	{8'd135,8'd164} : s = 301;
	{8'd135,8'd165} : s = 149;
	{8'd135,8'd166} : s = 299;
	{8'd135,8'd167} : s = 295;
	{8'd135,8'd168} : s = 423;
	{8'd135,8'd169} : s = 41;
	{8'd135,8'd170} : s = 147;
	{8'd135,8'd171} : s = 142;
	{8'd135,8'd172} : s = 286;
	{8'd135,8'd173} : s = 141;
	{8'd135,8'd174} : s = 285;
	{8'd135,8'd175} : s = 283;
	{8'd135,8'd176} : s = 414;
	{8'd135,8'd177} : s = 139;
	{8'd135,8'd178} : s = 279;
	{8'd135,8'd179} : s = 271;
	{8'd135,8'd180} : s = 413;
	{8'd135,8'd181} : s = 248;
	{8'd135,8'd182} : s = 411;
	{8'd135,8'd183} : s = 407;
	{8'd135,8'd184} : s = 491;
	{8'd135,8'd185} : s = 5;
	{8'd135,8'd186} : s = 38;
	{8'd135,8'd187} : s = 37;
	{8'd135,8'd188} : s = 135;
	{8'd135,8'd189} : s = 35;
	{8'd135,8'd190} : s = 120;
	{8'd135,8'd191} : s = 116;
	{8'd135,8'd192} : s = 244;
	{8'd135,8'd193} : s = 28;
	{8'd135,8'd194} : s = 114;
	{8'd135,8'd195} : s = 113;
	{8'd135,8'd196} : s = 242;
	{8'd135,8'd197} : s = 108;
	{8'd135,8'd198} : s = 241;
	{8'd135,8'd199} : s = 236;
	{8'd135,8'd200} : s = 399;
	{8'd135,8'd201} : s = 26;
	{8'd135,8'd202} : s = 106;
	{8'd135,8'd203} : s = 105;
	{8'd135,8'd204} : s = 234;
	{8'd135,8'd205} : s = 102;
	{8'd135,8'd206} : s = 233;
	{8'd135,8'd207} : s = 230;
	{8'd135,8'd208} : s = 380;
	{8'd135,8'd209} : s = 101;
	{8'd135,8'd210} : s = 229;
	{8'd135,8'd211} : s = 227;
	{8'd135,8'd212} : s = 378;
	{8'd135,8'd213} : s = 220;
	{8'd135,8'd214} : s = 377;
	{8'd135,8'd215} : s = 374;
	{8'd135,8'd216} : s = 487;
	{8'd135,8'd217} : s = 25;
	{8'd135,8'd218} : s = 99;
	{8'd135,8'd219} : s = 92;
	{8'd135,8'd220} : s = 218;
	{8'd135,8'd221} : s = 90;
	{8'd135,8'd222} : s = 217;
	{8'd135,8'd223} : s = 214;
	{8'd135,8'd224} : s = 373;
	{8'd135,8'd225} : s = 89;
	{8'd135,8'd226} : s = 213;
	{8'd135,8'd227} : s = 211;
	{8'd135,8'd228} : s = 371;
	{8'd135,8'd229} : s = 206;
	{8'd135,8'd230} : s = 366;
	{8'd135,8'd231} : s = 365;
	{8'd135,8'd232} : s = 478;
	{8'd135,8'd233} : s = 86;
	{8'd135,8'd234} : s = 205;
	{8'd135,8'd235} : s = 203;
	{8'd135,8'd236} : s = 363;
	{8'd135,8'd237} : s = 199;
	{8'd135,8'd238} : s = 359;
	{8'd135,8'd239} : s = 350;
	{8'd135,8'd240} : s = 477;
	{8'd135,8'd241} : s = 188;
	{8'd135,8'd242} : s = 349;
	{8'd135,8'd243} : s = 347;
	{8'd135,8'd244} : s = 475;
	{8'd135,8'd245} : s = 343;
	{8'd135,8'd246} : s = 471;
	{8'd135,8'd247} : s = 463;
	{8'd135,8'd248} : s = 509;
	{8'd135,8'd249} : s = 3;
	{8'd135,8'd250} : s = 22;
	{8'd135,8'd251} : s = 21;
	{8'd135,8'd252} : s = 85;
	{8'd135,8'd253} : s = 19;
	{8'd135,8'd254} : s = 83;
	{8'd135,8'd255} : s = 78;
	{8'd136,8'd0} : s = 34;
	{8'd136,8'd1} : s = 161;
	{8'd136,8'd2} : s = 152;
	{8'd136,8'd3} : s = 312;
	{8'd136,8'd4} : s = 148;
	{8'd136,8'd5} : s = 308;
	{8'd136,8'd6} : s = 306;
	{8'd136,8'd7} : s = 425;
	{8'd136,8'd8} : s = 33;
	{8'd136,8'd9} : s = 146;
	{8'd136,8'd10} : s = 145;
	{8'd136,8'd11} : s = 305;
	{8'd136,8'd12} : s = 140;
	{8'd136,8'd13} : s = 300;
	{8'd136,8'd14} : s = 298;
	{8'd136,8'd15} : s = 422;
	{8'd136,8'd16} : s = 138;
	{8'd136,8'd17} : s = 297;
	{8'd136,8'd18} : s = 294;
	{8'd136,8'd19} : s = 421;
	{8'd136,8'd20} : s = 293;
	{8'd136,8'd21} : s = 419;
	{8'd136,8'd22} : s = 412;
	{8'd136,8'd23} : s = 486;
	{8'd136,8'd24} : s = 24;
	{8'd136,8'd25} : s = 137;
	{8'd136,8'd26} : s = 134;
	{8'd136,8'd27} : s = 291;
	{8'd136,8'd28} : s = 133;
	{8'd136,8'd29} : s = 284;
	{8'd136,8'd30} : s = 282;
	{8'd136,8'd31} : s = 410;
	{8'd136,8'd32} : s = 131;
	{8'd136,8'd33} : s = 281;
	{8'd136,8'd34} : s = 278;
	{8'd136,8'd35} : s = 409;
	{8'd136,8'd36} : s = 277;
	{8'd136,8'd37} : s = 406;
	{8'd136,8'd38} : s = 405;
	{8'd136,8'd39} : s = 485;
	{8'd136,8'd40} : s = 112;
	{8'd136,8'd41} : s = 275;
	{8'd136,8'd42} : s = 270;
	{8'd136,8'd43} : s = 403;
	{8'd136,8'd44} : s = 269;
	{8'd136,8'd45} : s = 398;
	{8'd136,8'd46} : s = 397;
	{8'd136,8'd47} : s = 483;
	{8'd136,8'd48} : s = 267;
	{8'd136,8'd49} : s = 395;
	{8'd136,8'd50} : s = 391;
	{8'd136,8'd51} : s = 476;
	{8'd136,8'd52} : s = 376;
	{8'd136,8'd53} : s = 474;
	{8'd136,8'd54} : s = 473;
	{8'd136,8'd55} : s = 506;
	{8'd136,8'd56} : s = 20;
	{8'd136,8'd57} : s = 104;
	{8'd136,8'd58} : s = 100;
	{8'd136,8'd59} : s = 263;
	{8'd136,8'd60} : s = 98;
	{8'd136,8'd61} : s = 240;
	{8'd136,8'd62} : s = 232;
	{8'd136,8'd63} : s = 372;
	{8'd136,8'd64} : s = 97;
	{8'd136,8'd65} : s = 228;
	{8'd136,8'd66} : s = 226;
	{8'd136,8'd67} : s = 370;
	{8'd136,8'd68} : s = 225;
	{8'd136,8'd69} : s = 369;
	{8'd136,8'd70} : s = 364;
	{8'd136,8'd71} : s = 470;
	{8'd136,8'd72} : s = 88;
	{8'd136,8'd73} : s = 216;
	{8'd136,8'd74} : s = 212;
	{8'd136,8'd75} : s = 362;
	{8'd136,8'd76} : s = 210;
	{8'd136,8'd77} : s = 361;
	{8'd136,8'd78} : s = 358;
	{8'd136,8'd79} : s = 469;
	{8'd136,8'd80} : s = 209;
	{8'd136,8'd81} : s = 357;
	{8'd136,8'd82} : s = 355;
	{8'd136,8'd83} : s = 467;
	{8'd136,8'd84} : s = 348;
	{8'd136,8'd85} : s = 462;
	{8'd136,8'd86} : s = 461;
	{8'd136,8'd87} : s = 505;
	{8'd136,8'd88} : s = 84;
	{8'd136,8'd89} : s = 204;
	{8'd136,8'd90} : s = 202;
	{8'd136,8'd91} : s = 346;
	{8'd136,8'd92} : s = 201;
	{8'd136,8'd93} : s = 345;
	{8'd136,8'd94} : s = 342;
	{8'd136,8'd95} : s = 459;
	{8'd136,8'd96} : s = 198;
	{8'd136,8'd97} : s = 341;
	{8'd136,8'd98} : s = 339;
	{8'd136,8'd99} : s = 455;
	{8'd136,8'd100} : s = 334;
	{8'd136,8'd101} : s = 444;
	{8'd136,8'd102} : s = 442;
	{8'd136,8'd103} : s = 502;
	{8'd136,8'd104} : s = 197;
	{8'd136,8'd105} : s = 333;
	{8'd136,8'd106} : s = 331;
	{8'd136,8'd107} : s = 441;
	{8'd136,8'd108} : s = 327;
	{8'd136,8'd109} : s = 438;
	{8'd136,8'd110} : s = 437;
	{8'd136,8'd111} : s = 501;
	{8'd136,8'd112} : s = 316;
	{8'd136,8'd113} : s = 435;
	{8'd136,8'd114} : s = 430;
	{8'd136,8'd115} : s = 499;
	{8'd136,8'd116} : s = 429;
	{8'd136,8'd117} : s = 494;
	{8'd136,8'd118} : s = 493;
	{8'd136,8'd119} : s = 510;
	{8'd136,8'd120} : s = 1;
	{8'd136,8'd121} : s = 18;
	{8'd136,8'd122} : s = 17;
	{8'd136,8'd123} : s = 82;
	{8'd136,8'd124} : s = 12;
	{8'd136,8'd125} : s = 81;
	{8'd136,8'd126} : s = 76;
	{8'd136,8'd127} : s = 195;
	{8'd136,8'd128} : s = 10;
	{8'd136,8'd129} : s = 74;
	{8'd136,8'd130} : s = 73;
	{8'd136,8'd131} : s = 184;
	{8'd136,8'd132} : s = 70;
	{8'd136,8'd133} : s = 180;
	{8'd136,8'd134} : s = 178;
	{8'd136,8'd135} : s = 314;
	{8'd136,8'd136} : s = 9;
	{8'd136,8'd137} : s = 69;
	{8'd136,8'd138} : s = 67;
	{8'd136,8'd139} : s = 177;
	{8'd136,8'd140} : s = 56;
	{8'd136,8'd141} : s = 172;
	{8'd136,8'd142} : s = 170;
	{8'd136,8'd143} : s = 313;
	{8'd136,8'd144} : s = 52;
	{8'd136,8'd145} : s = 169;
	{8'd136,8'd146} : s = 166;
	{8'd136,8'd147} : s = 310;
	{8'd136,8'd148} : s = 165;
	{8'd136,8'd149} : s = 309;
	{8'd136,8'd150} : s = 307;
	{8'd136,8'd151} : s = 427;
	{8'd136,8'd152} : s = 6;
	{8'd136,8'd153} : s = 50;
	{8'd136,8'd154} : s = 49;
	{8'd136,8'd155} : s = 163;
	{8'd136,8'd156} : s = 44;
	{8'd136,8'd157} : s = 156;
	{8'd136,8'd158} : s = 154;
	{8'd136,8'd159} : s = 302;
	{8'd136,8'd160} : s = 42;
	{8'd136,8'd161} : s = 153;
	{8'd136,8'd162} : s = 150;
	{8'd136,8'd163} : s = 301;
	{8'd136,8'd164} : s = 149;
	{8'd136,8'd165} : s = 299;
	{8'd136,8'd166} : s = 295;
	{8'd136,8'd167} : s = 423;
	{8'd136,8'd168} : s = 41;
	{8'd136,8'd169} : s = 147;
	{8'd136,8'd170} : s = 142;
	{8'd136,8'd171} : s = 286;
	{8'd136,8'd172} : s = 141;
	{8'd136,8'd173} : s = 285;
	{8'd136,8'd174} : s = 283;
	{8'd136,8'd175} : s = 414;
	{8'd136,8'd176} : s = 139;
	{8'd136,8'd177} : s = 279;
	{8'd136,8'd178} : s = 271;
	{8'd136,8'd179} : s = 413;
	{8'd136,8'd180} : s = 248;
	{8'd136,8'd181} : s = 411;
	{8'd136,8'd182} : s = 407;
	{8'd136,8'd183} : s = 491;
	{8'd136,8'd184} : s = 5;
	{8'd136,8'd185} : s = 38;
	{8'd136,8'd186} : s = 37;
	{8'd136,8'd187} : s = 135;
	{8'd136,8'd188} : s = 35;
	{8'd136,8'd189} : s = 120;
	{8'd136,8'd190} : s = 116;
	{8'd136,8'd191} : s = 244;
	{8'd136,8'd192} : s = 28;
	{8'd136,8'd193} : s = 114;
	{8'd136,8'd194} : s = 113;
	{8'd136,8'd195} : s = 242;
	{8'd136,8'd196} : s = 108;
	{8'd136,8'd197} : s = 241;
	{8'd136,8'd198} : s = 236;
	{8'd136,8'd199} : s = 399;
	{8'd136,8'd200} : s = 26;
	{8'd136,8'd201} : s = 106;
	{8'd136,8'd202} : s = 105;
	{8'd136,8'd203} : s = 234;
	{8'd136,8'd204} : s = 102;
	{8'd136,8'd205} : s = 233;
	{8'd136,8'd206} : s = 230;
	{8'd136,8'd207} : s = 380;
	{8'd136,8'd208} : s = 101;
	{8'd136,8'd209} : s = 229;
	{8'd136,8'd210} : s = 227;
	{8'd136,8'd211} : s = 378;
	{8'd136,8'd212} : s = 220;
	{8'd136,8'd213} : s = 377;
	{8'd136,8'd214} : s = 374;
	{8'd136,8'd215} : s = 487;
	{8'd136,8'd216} : s = 25;
	{8'd136,8'd217} : s = 99;
	{8'd136,8'd218} : s = 92;
	{8'd136,8'd219} : s = 218;
	{8'd136,8'd220} : s = 90;
	{8'd136,8'd221} : s = 217;
	{8'd136,8'd222} : s = 214;
	{8'd136,8'd223} : s = 373;
	{8'd136,8'd224} : s = 89;
	{8'd136,8'd225} : s = 213;
	{8'd136,8'd226} : s = 211;
	{8'd136,8'd227} : s = 371;
	{8'd136,8'd228} : s = 206;
	{8'd136,8'd229} : s = 366;
	{8'd136,8'd230} : s = 365;
	{8'd136,8'd231} : s = 478;
	{8'd136,8'd232} : s = 86;
	{8'd136,8'd233} : s = 205;
	{8'd136,8'd234} : s = 203;
	{8'd136,8'd235} : s = 363;
	{8'd136,8'd236} : s = 199;
	{8'd136,8'd237} : s = 359;
	{8'd136,8'd238} : s = 350;
	{8'd136,8'd239} : s = 477;
	{8'd136,8'd240} : s = 188;
	{8'd136,8'd241} : s = 349;
	{8'd136,8'd242} : s = 347;
	{8'd136,8'd243} : s = 475;
	{8'd136,8'd244} : s = 343;
	{8'd136,8'd245} : s = 471;
	{8'd136,8'd246} : s = 463;
	{8'd136,8'd247} : s = 509;
	{8'd136,8'd248} : s = 3;
	{8'd136,8'd249} : s = 22;
	{8'd136,8'd250} : s = 21;
	{8'd136,8'd251} : s = 85;
	{8'd136,8'd252} : s = 19;
	{8'd136,8'd253} : s = 83;
	{8'd136,8'd254} : s = 78;
	{8'd136,8'd255} : s = 186;
	{8'd137,8'd0} : s = 161;
	{8'd137,8'd1} : s = 152;
	{8'd137,8'd2} : s = 312;
	{8'd137,8'd3} : s = 148;
	{8'd137,8'd4} : s = 308;
	{8'd137,8'd5} : s = 306;
	{8'd137,8'd6} : s = 425;
	{8'd137,8'd7} : s = 33;
	{8'd137,8'd8} : s = 146;
	{8'd137,8'd9} : s = 145;
	{8'd137,8'd10} : s = 305;
	{8'd137,8'd11} : s = 140;
	{8'd137,8'd12} : s = 300;
	{8'd137,8'd13} : s = 298;
	{8'd137,8'd14} : s = 422;
	{8'd137,8'd15} : s = 138;
	{8'd137,8'd16} : s = 297;
	{8'd137,8'd17} : s = 294;
	{8'd137,8'd18} : s = 421;
	{8'd137,8'd19} : s = 293;
	{8'd137,8'd20} : s = 419;
	{8'd137,8'd21} : s = 412;
	{8'd137,8'd22} : s = 486;
	{8'd137,8'd23} : s = 24;
	{8'd137,8'd24} : s = 137;
	{8'd137,8'd25} : s = 134;
	{8'd137,8'd26} : s = 291;
	{8'd137,8'd27} : s = 133;
	{8'd137,8'd28} : s = 284;
	{8'd137,8'd29} : s = 282;
	{8'd137,8'd30} : s = 410;
	{8'd137,8'd31} : s = 131;
	{8'd137,8'd32} : s = 281;
	{8'd137,8'd33} : s = 278;
	{8'd137,8'd34} : s = 409;
	{8'd137,8'd35} : s = 277;
	{8'd137,8'd36} : s = 406;
	{8'd137,8'd37} : s = 405;
	{8'd137,8'd38} : s = 485;
	{8'd137,8'd39} : s = 112;
	{8'd137,8'd40} : s = 275;
	{8'd137,8'd41} : s = 270;
	{8'd137,8'd42} : s = 403;
	{8'd137,8'd43} : s = 269;
	{8'd137,8'd44} : s = 398;
	{8'd137,8'd45} : s = 397;
	{8'd137,8'd46} : s = 483;
	{8'd137,8'd47} : s = 267;
	{8'd137,8'd48} : s = 395;
	{8'd137,8'd49} : s = 391;
	{8'd137,8'd50} : s = 476;
	{8'd137,8'd51} : s = 376;
	{8'd137,8'd52} : s = 474;
	{8'd137,8'd53} : s = 473;
	{8'd137,8'd54} : s = 506;
	{8'd137,8'd55} : s = 20;
	{8'd137,8'd56} : s = 104;
	{8'd137,8'd57} : s = 100;
	{8'd137,8'd58} : s = 263;
	{8'd137,8'd59} : s = 98;
	{8'd137,8'd60} : s = 240;
	{8'd137,8'd61} : s = 232;
	{8'd137,8'd62} : s = 372;
	{8'd137,8'd63} : s = 97;
	{8'd137,8'd64} : s = 228;
	{8'd137,8'd65} : s = 226;
	{8'd137,8'd66} : s = 370;
	{8'd137,8'd67} : s = 225;
	{8'd137,8'd68} : s = 369;
	{8'd137,8'd69} : s = 364;
	{8'd137,8'd70} : s = 470;
	{8'd137,8'd71} : s = 88;
	{8'd137,8'd72} : s = 216;
	{8'd137,8'd73} : s = 212;
	{8'd137,8'd74} : s = 362;
	{8'd137,8'd75} : s = 210;
	{8'd137,8'd76} : s = 361;
	{8'd137,8'd77} : s = 358;
	{8'd137,8'd78} : s = 469;
	{8'd137,8'd79} : s = 209;
	{8'd137,8'd80} : s = 357;
	{8'd137,8'd81} : s = 355;
	{8'd137,8'd82} : s = 467;
	{8'd137,8'd83} : s = 348;
	{8'd137,8'd84} : s = 462;
	{8'd137,8'd85} : s = 461;
	{8'd137,8'd86} : s = 505;
	{8'd137,8'd87} : s = 84;
	{8'd137,8'd88} : s = 204;
	{8'd137,8'd89} : s = 202;
	{8'd137,8'd90} : s = 346;
	{8'd137,8'd91} : s = 201;
	{8'd137,8'd92} : s = 345;
	{8'd137,8'd93} : s = 342;
	{8'd137,8'd94} : s = 459;
	{8'd137,8'd95} : s = 198;
	{8'd137,8'd96} : s = 341;
	{8'd137,8'd97} : s = 339;
	{8'd137,8'd98} : s = 455;
	{8'd137,8'd99} : s = 334;
	{8'd137,8'd100} : s = 444;
	{8'd137,8'd101} : s = 442;
	{8'd137,8'd102} : s = 502;
	{8'd137,8'd103} : s = 197;
	{8'd137,8'd104} : s = 333;
	{8'd137,8'd105} : s = 331;
	{8'd137,8'd106} : s = 441;
	{8'd137,8'd107} : s = 327;
	{8'd137,8'd108} : s = 438;
	{8'd137,8'd109} : s = 437;
	{8'd137,8'd110} : s = 501;
	{8'd137,8'd111} : s = 316;
	{8'd137,8'd112} : s = 435;
	{8'd137,8'd113} : s = 430;
	{8'd137,8'd114} : s = 499;
	{8'd137,8'd115} : s = 429;
	{8'd137,8'd116} : s = 494;
	{8'd137,8'd117} : s = 493;
	{8'd137,8'd118} : s = 510;
	{8'd137,8'd119} : s = 1;
	{8'd137,8'd120} : s = 18;
	{8'd137,8'd121} : s = 17;
	{8'd137,8'd122} : s = 82;
	{8'd137,8'd123} : s = 12;
	{8'd137,8'd124} : s = 81;
	{8'd137,8'd125} : s = 76;
	{8'd137,8'd126} : s = 195;
	{8'd137,8'd127} : s = 10;
	{8'd137,8'd128} : s = 74;
	{8'd137,8'd129} : s = 73;
	{8'd137,8'd130} : s = 184;
	{8'd137,8'd131} : s = 70;
	{8'd137,8'd132} : s = 180;
	{8'd137,8'd133} : s = 178;
	{8'd137,8'd134} : s = 314;
	{8'd137,8'd135} : s = 9;
	{8'd137,8'd136} : s = 69;
	{8'd137,8'd137} : s = 67;
	{8'd137,8'd138} : s = 177;
	{8'd137,8'd139} : s = 56;
	{8'd137,8'd140} : s = 172;
	{8'd137,8'd141} : s = 170;
	{8'd137,8'd142} : s = 313;
	{8'd137,8'd143} : s = 52;
	{8'd137,8'd144} : s = 169;
	{8'd137,8'd145} : s = 166;
	{8'd137,8'd146} : s = 310;
	{8'd137,8'd147} : s = 165;
	{8'd137,8'd148} : s = 309;
	{8'd137,8'd149} : s = 307;
	{8'd137,8'd150} : s = 427;
	{8'd137,8'd151} : s = 6;
	{8'd137,8'd152} : s = 50;
	{8'd137,8'd153} : s = 49;
	{8'd137,8'd154} : s = 163;
	{8'd137,8'd155} : s = 44;
	{8'd137,8'd156} : s = 156;
	{8'd137,8'd157} : s = 154;
	{8'd137,8'd158} : s = 302;
	{8'd137,8'd159} : s = 42;
	{8'd137,8'd160} : s = 153;
	{8'd137,8'd161} : s = 150;
	{8'd137,8'd162} : s = 301;
	{8'd137,8'd163} : s = 149;
	{8'd137,8'd164} : s = 299;
	{8'd137,8'd165} : s = 295;
	{8'd137,8'd166} : s = 423;
	{8'd137,8'd167} : s = 41;
	{8'd137,8'd168} : s = 147;
	{8'd137,8'd169} : s = 142;
	{8'd137,8'd170} : s = 286;
	{8'd137,8'd171} : s = 141;
	{8'd137,8'd172} : s = 285;
	{8'd137,8'd173} : s = 283;
	{8'd137,8'd174} : s = 414;
	{8'd137,8'd175} : s = 139;
	{8'd137,8'd176} : s = 279;
	{8'd137,8'd177} : s = 271;
	{8'd137,8'd178} : s = 413;
	{8'd137,8'd179} : s = 248;
	{8'd137,8'd180} : s = 411;
	{8'd137,8'd181} : s = 407;
	{8'd137,8'd182} : s = 491;
	{8'd137,8'd183} : s = 5;
	{8'd137,8'd184} : s = 38;
	{8'd137,8'd185} : s = 37;
	{8'd137,8'd186} : s = 135;
	{8'd137,8'd187} : s = 35;
	{8'd137,8'd188} : s = 120;
	{8'd137,8'd189} : s = 116;
	{8'd137,8'd190} : s = 244;
	{8'd137,8'd191} : s = 28;
	{8'd137,8'd192} : s = 114;
	{8'd137,8'd193} : s = 113;
	{8'd137,8'd194} : s = 242;
	{8'd137,8'd195} : s = 108;
	{8'd137,8'd196} : s = 241;
	{8'd137,8'd197} : s = 236;
	{8'd137,8'd198} : s = 399;
	{8'd137,8'd199} : s = 26;
	{8'd137,8'd200} : s = 106;
	{8'd137,8'd201} : s = 105;
	{8'd137,8'd202} : s = 234;
	{8'd137,8'd203} : s = 102;
	{8'd137,8'd204} : s = 233;
	{8'd137,8'd205} : s = 230;
	{8'd137,8'd206} : s = 380;
	{8'd137,8'd207} : s = 101;
	{8'd137,8'd208} : s = 229;
	{8'd137,8'd209} : s = 227;
	{8'd137,8'd210} : s = 378;
	{8'd137,8'd211} : s = 220;
	{8'd137,8'd212} : s = 377;
	{8'd137,8'd213} : s = 374;
	{8'd137,8'd214} : s = 487;
	{8'd137,8'd215} : s = 25;
	{8'd137,8'd216} : s = 99;
	{8'd137,8'd217} : s = 92;
	{8'd137,8'd218} : s = 218;
	{8'd137,8'd219} : s = 90;
	{8'd137,8'd220} : s = 217;
	{8'd137,8'd221} : s = 214;
	{8'd137,8'd222} : s = 373;
	{8'd137,8'd223} : s = 89;
	{8'd137,8'd224} : s = 213;
	{8'd137,8'd225} : s = 211;
	{8'd137,8'd226} : s = 371;
	{8'd137,8'd227} : s = 206;
	{8'd137,8'd228} : s = 366;
	{8'd137,8'd229} : s = 365;
	{8'd137,8'd230} : s = 478;
	{8'd137,8'd231} : s = 86;
	{8'd137,8'd232} : s = 205;
	{8'd137,8'd233} : s = 203;
	{8'd137,8'd234} : s = 363;
	{8'd137,8'd235} : s = 199;
	{8'd137,8'd236} : s = 359;
	{8'd137,8'd237} : s = 350;
	{8'd137,8'd238} : s = 477;
	{8'd137,8'd239} : s = 188;
	{8'd137,8'd240} : s = 349;
	{8'd137,8'd241} : s = 347;
	{8'd137,8'd242} : s = 475;
	{8'd137,8'd243} : s = 343;
	{8'd137,8'd244} : s = 471;
	{8'd137,8'd245} : s = 463;
	{8'd137,8'd246} : s = 509;
	{8'd137,8'd247} : s = 3;
	{8'd137,8'd248} : s = 22;
	{8'd137,8'd249} : s = 21;
	{8'd137,8'd250} : s = 85;
	{8'd137,8'd251} : s = 19;
	{8'd137,8'd252} : s = 83;
	{8'd137,8'd253} : s = 78;
	{8'd137,8'd254} : s = 186;
	{8'd137,8'd255} : s = 14;
	{8'd138,8'd0} : s = 152;
	{8'd138,8'd1} : s = 312;
	{8'd138,8'd2} : s = 148;
	{8'd138,8'd3} : s = 308;
	{8'd138,8'd4} : s = 306;
	{8'd138,8'd5} : s = 425;
	{8'd138,8'd6} : s = 33;
	{8'd138,8'd7} : s = 146;
	{8'd138,8'd8} : s = 145;
	{8'd138,8'd9} : s = 305;
	{8'd138,8'd10} : s = 140;
	{8'd138,8'd11} : s = 300;
	{8'd138,8'd12} : s = 298;
	{8'd138,8'd13} : s = 422;
	{8'd138,8'd14} : s = 138;
	{8'd138,8'd15} : s = 297;
	{8'd138,8'd16} : s = 294;
	{8'd138,8'd17} : s = 421;
	{8'd138,8'd18} : s = 293;
	{8'd138,8'd19} : s = 419;
	{8'd138,8'd20} : s = 412;
	{8'd138,8'd21} : s = 486;
	{8'd138,8'd22} : s = 24;
	{8'd138,8'd23} : s = 137;
	{8'd138,8'd24} : s = 134;
	{8'd138,8'd25} : s = 291;
	{8'd138,8'd26} : s = 133;
	{8'd138,8'd27} : s = 284;
	{8'd138,8'd28} : s = 282;
	{8'd138,8'd29} : s = 410;
	{8'd138,8'd30} : s = 131;
	{8'd138,8'd31} : s = 281;
	{8'd138,8'd32} : s = 278;
	{8'd138,8'd33} : s = 409;
	{8'd138,8'd34} : s = 277;
	{8'd138,8'd35} : s = 406;
	{8'd138,8'd36} : s = 405;
	{8'd138,8'd37} : s = 485;
	{8'd138,8'd38} : s = 112;
	{8'd138,8'd39} : s = 275;
	{8'd138,8'd40} : s = 270;
	{8'd138,8'd41} : s = 403;
	{8'd138,8'd42} : s = 269;
	{8'd138,8'd43} : s = 398;
	{8'd138,8'd44} : s = 397;
	{8'd138,8'd45} : s = 483;
	{8'd138,8'd46} : s = 267;
	{8'd138,8'd47} : s = 395;
	{8'd138,8'd48} : s = 391;
	{8'd138,8'd49} : s = 476;
	{8'd138,8'd50} : s = 376;
	{8'd138,8'd51} : s = 474;
	{8'd138,8'd52} : s = 473;
	{8'd138,8'd53} : s = 506;
	{8'd138,8'd54} : s = 20;
	{8'd138,8'd55} : s = 104;
	{8'd138,8'd56} : s = 100;
	{8'd138,8'd57} : s = 263;
	{8'd138,8'd58} : s = 98;
	{8'd138,8'd59} : s = 240;
	{8'd138,8'd60} : s = 232;
	{8'd138,8'd61} : s = 372;
	{8'd138,8'd62} : s = 97;
	{8'd138,8'd63} : s = 228;
	{8'd138,8'd64} : s = 226;
	{8'd138,8'd65} : s = 370;
	{8'd138,8'd66} : s = 225;
	{8'd138,8'd67} : s = 369;
	{8'd138,8'd68} : s = 364;
	{8'd138,8'd69} : s = 470;
	{8'd138,8'd70} : s = 88;
	{8'd138,8'd71} : s = 216;
	{8'd138,8'd72} : s = 212;
	{8'd138,8'd73} : s = 362;
	{8'd138,8'd74} : s = 210;
	{8'd138,8'd75} : s = 361;
	{8'd138,8'd76} : s = 358;
	{8'd138,8'd77} : s = 469;
	{8'd138,8'd78} : s = 209;
	{8'd138,8'd79} : s = 357;
	{8'd138,8'd80} : s = 355;
	{8'd138,8'd81} : s = 467;
	{8'd138,8'd82} : s = 348;
	{8'd138,8'd83} : s = 462;
	{8'd138,8'd84} : s = 461;
	{8'd138,8'd85} : s = 505;
	{8'd138,8'd86} : s = 84;
	{8'd138,8'd87} : s = 204;
	{8'd138,8'd88} : s = 202;
	{8'd138,8'd89} : s = 346;
	{8'd138,8'd90} : s = 201;
	{8'd138,8'd91} : s = 345;
	{8'd138,8'd92} : s = 342;
	{8'd138,8'd93} : s = 459;
	{8'd138,8'd94} : s = 198;
	{8'd138,8'd95} : s = 341;
	{8'd138,8'd96} : s = 339;
	{8'd138,8'd97} : s = 455;
	{8'd138,8'd98} : s = 334;
	{8'd138,8'd99} : s = 444;
	{8'd138,8'd100} : s = 442;
	{8'd138,8'd101} : s = 502;
	{8'd138,8'd102} : s = 197;
	{8'd138,8'd103} : s = 333;
	{8'd138,8'd104} : s = 331;
	{8'd138,8'd105} : s = 441;
	{8'd138,8'd106} : s = 327;
	{8'd138,8'd107} : s = 438;
	{8'd138,8'd108} : s = 437;
	{8'd138,8'd109} : s = 501;
	{8'd138,8'd110} : s = 316;
	{8'd138,8'd111} : s = 435;
	{8'd138,8'd112} : s = 430;
	{8'd138,8'd113} : s = 499;
	{8'd138,8'd114} : s = 429;
	{8'd138,8'd115} : s = 494;
	{8'd138,8'd116} : s = 493;
	{8'd138,8'd117} : s = 510;
	{8'd138,8'd118} : s = 1;
	{8'd138,8'd119} : s = 18;
	{8'd138,8'd120} : s = 17;
	{8'd138,8'd121} : s = 82;
	{8'd138,8'd122} : s = 12;
	{8'd138,8'd123} : s = 81;
	{8'd138,8'd124} : s = 76;
	{8'd138,8'd125} : s = 195;
	{8'd138,8'd126} : s = 10;
	{8'd138,8'd127} : s = 74;
	{8'd138,8'd128} : s = 73;
	{8'd138,8'd129} : s = 184;
	{8'd138,8'd130} : s = 70;
	{8'd138,8'd131} : s = 180;
	{8'd138,8'd132} : s = 178;
	{8'd138,8'd133} : s = 314;
	{8'd138,8'd134} : s = 9;
	{8'd138,8'd135} : s = 69;
	{8'd138,8'd136} : s = 67;
	{8'd138,8'd137} : s = 177;
	{8'd138,8'd138} : s = 56;
	{8'd138,8'd139} : s = 172;
	{8'd138,8'd140} : s = 170;
	{8'd138,8'd141} : s = 313;
	{8'd138,8'd142} : s = 52;
	{8'd138,8'd143} : s = 169;
	{8'd138,8'd144} : s = 166;
	{8'd138,8'd145} : s = 310;
	{8'd138,8'd146} : s = 165;
	{8'd138,8'd147} : s = 309;
	{8'd138,8'd148} : s = 307;
	{8'd138,8'd149} : s = 427;
	{8'd138,8'd150} : s = 6;
	{8'd138,8'd151} : s = 50;
	{8'd138,8'd152} : s = 49;
	{8'd138,8'd153} : s = 163;
	{8'd138,8'd154} : s = 44;
	{8'd138,8'd155} : s = 156;
	{8'd138,8'd156} : s = 154;
	{8'd138,8'd157} : s = 302;
	{8'd138,8'd158} : s = 42;
	{8'd138,8'd159} : s = 153;
	{8'd138,8'd160} : s = 150;
	{8'd138,8'd161} : s = 301;
	{8'd138,8'd162} : s = 149;
	{8'd138,8'd163} : s = 299;
	{8'd138,8'd164} : s = 295;
	{8'd138,8'd165} : s = 423;
	{8'd138,8'd166} : s = 41;
	{8'd138,8'd167} : s = 147;
	{8'd138,8'd168} : s = 142;
	{8'd138,8'd169} : s = 286;
	{8'd138,8'd170} : s = 141;
	{8'd138,8'd171} : s = 285;
	{8'd138,8'd172} : s = 283;
	{8'd138,8'd173} : s = 414;
	{8'd138,8'd174} : s = 139;
	{8'd138,8'd175} : s = 279;
	{8'd138,8'd176} : s = 271;
	{8'd138,8'd177} : s = 413;
	{8'd138,8'd178} : s = 248;
	{8'd138,8'd179} : s = 411;
	{8'd138,8'd180} : s = 407;
	{8'd138,8'd181} : s = 491;
	{8'd138,8'd182} : s = 5;
	{8'd138,8'd183} : s = 38;
	{8'd138,8'd184} : s = 37;
	{8'd138,8'd185} : s = 135;
	{8'd138,8'd186} : s = 35;
	{8'd138,8'd187} : s = 120;
	{8'd138,8'd188} : s = 116;
	{8'd138,8'd189} : s = 244;
	{8'd138,8'd190} : s = 28;
	{8'd138,8'd191} : s = 114;
	{8'd138,8'd192} : s = 113;
	{8'd138,8'd193} : s = 242;
	{8'd138,8'd194} : s = 108;
	{8'd138,8'd195} : s = 241;
	{8'd138,8'd196} : s = 236;
	{8'd138,8'd197} : s = 399;
	{8'd138,8'd198} : s = 26;
	{8'd138,8'd199} : s = 106;
	{8'd138,8'd200} : s = 105;
	{8'd138,8'd201} : s = 234;
	{8'd138,8'd202} : s = 102;
	{8'd138,8'd203} : s = 233;
	{8'd138,8'd204} : s = 230;
	{8'd138,8'd205} : s = 380;
	{8'd138,8'd206} : s = 101;
	{8'd138,8'd207} : s = 229;
	{8'd138,8'd208} : s = 227;
	{8'd138,8'd209} : s = 378;
	{8'd138,8'd210} : s = 220;
	{8'd138,8'd211} : s = 377;
	{8'd138,8'd212} : s = 374;
	{8'd138,8'd213} : s = 487;
	{8'd138,8'd214} : s = 25;
	{8'd138,8'd215} : s = 99;
	{8'd138,8'd216} : s = 92;
	{8'd138,8'd217} : s = 218;
	{8'd138,8'd218} : s = 90;
	{8'd138,8'd219} : s = 217;
	{8'd138,8'd220} : s = 214;
	{8'd138,8'd221} : s = 373;
	{8'd138,8'd222} : s = 89;
	{8'd138,8'd223} : s = 213;
	{8'd138,8'd224} : s = 211;
	{8'd138,8'd225} : s = 371;
	{8'd138,8'd226} : s = 206;
	{8'd138,8'd227} : s = 366;
	{8'd138,8'd228} : s = 365;
	{8'd138,8'd229} : s = 478;
	{8'd138,8'd230} : s = 86;
	{8'd138,8'd231} : s = 205;
	{8'd138,8'd232} : s = 203;
	{8'd138,8'd233} : s = 363;
	{8'd138,8'd234} : s = 199;
	{8'd138,8'd235} : s = 359;
	{8'd138,8'd236} : s = 350;
	{8'd138,8'd237} : s = 477;
	{8'd138,8'd238} : s = 188;
	{8'd138,8'd239} : s = 349;
	{8'd138,8'd240} : s = 347;
	{8'd138,8'd241} : s = 475;
	{8'd138,8'd242} : s = 343;
	{8'd138,8'd243} : s = 471;
	{8'd138,8'd244} : s = 463;
	{8'd138,8'd245} : s = 509;
	{8'd138,8'd246} : s = 3;
	{8'd138,8'd247} : s = 22;
	{8'd138,8'd248} : s = 21;
	{8'd138,8'd249} : s = 85;
	{8'd138,8'd250} : s = 19;
	{8'd138,8'd251} : s = 83;
	{8'd138,8'd252} : s = 78;
	{8'd138,8'd253} : s = 186;
	{8'd138,8'd254} : s = 14;
	{8'd138,8'd255} : s = 77;
	{8'd139,8'd0} : s = 312;
	{8'd139,8'd1} : s = 148;
	{8'd139,8'd2} : s = 308;
	{8'd139,8'd3} : s = 306;
	{8'd139,8'd4} : s = 425;
	{8'd139,8'd5} : s = 33;
	{8'd139,8'd6} : s = 146;
	{8'd139,8'd7} : s = 145;
	{8'd139,8'd8} : s = 305;
	{8'd139,8'd9} : s = 140;
	{8'd139,8'd10} : s = 300;
	{8'd139,8'd11} : s = 298;
	{8'd139,8'd12} : s = 422;
	{8'd139,8'd13} : s = 138;
	{8'd139,8'd14} : s = 297;
	{8'd139,8'd15} : s = 294;
	{8'd139,8'd16} : s = 421;
	{8'd139,8'd17} : s = 293;
	{8'd139,8'd18} : s = 419;
	{8'd139,8'd19} : s = 412;
	{8'd139,8'd20} : s = 486;
	{8'd139,8'd21} : s = 24;
	{8'd139,8'd22} : s = 137;
	{8'd139,8'd23} : s = 134;
	{8'd139,8'd24} : s = 291;
	{8'd139,8'd25} : s = 133;
	{8'd139,8'd26} : s = 284;
	{8'd139,8'd27} : s = 282;
	{8'd139,8'd28} : s = 410;
	{8'd139,8'd29} : s = 131;
	{8'd139,8'd30} : s = 281;
	{8'd139,8'd31} : s = 278;
	{8'd139,8'd32} : s = 409;
	{8'd139,8'd33} : s = 277;
	{8'd139,8'd34} : s = 406;
	{8'd139,8'd35} : s = 405;
	{8'd139,8'd36} : s = 485;
	{8'd139,8'd37} : s = 112;
	{8'd139,8'd38} : s = 275;
	{8'd139,8'd39} : s = 270;
	{8'd139,8'd40} : s = 403;
	{8'd139,8'd41} : s = 269;
	{8'd139,8'd42} : s = 398;
	{8'd139,8'd43} : s = 397;
	{8'd139,8'd44} : s = 483;
	{8'd139,8'd45} : s = 267;
	{8'd139,8'd46} : s = 395;
	{8'd139,8'd47} : s = 391;
	{8'd139,8'd48} : s = 476;
	{8'd139,8'd49} : s = 376;
	{8'd139,8'd50} : s = 474;
	{8'd139,8'd51} : s = 473;
	{8'd139,8'd52} : s = 506;
	{8'd139,8'd53} : s = 20;
	{8'd139,8'd54} : s = 104;
	{8'd139,8'd55} : s = 100;
	{8'd139,8'd56} : s = 263;
	{8'd139,8'd57} : s = 98;
	{8'd139,8'd58} : s = 240;
	{8'd139,8'd59} : s = 232;
	{8'd139,8'd60} : s = 372;
	{8'd139,8'd61} : s = 97;
	{8'd139,8'd62} : s = 228;
	{8'd139,8'd63} : s = 226;
	{8'd139,8'd64} : s = 370;
	{8'd139,8'd65} : s = 225;
	{8'd139,8'd66} : s = 369;
	{8'd139,8'd67} : s = 364;
	{8'd139,8'd68} : s = 470;
	{8'd139,8'd69} : s = 88;
	{8'd139,8'd70} : s = 216;
	{8'd139,8'd71} : s = 212;
	{8'd139,8'd72} : s = 362;
	{8'd139,8'd73} : s = 210;
	{8'd139,8'd74} : s = 361;
	{8'd139,8'd75} : s = 358;
	{8'd139,8'd76} : s = 469;
	{8'd139,8'd77} : s = 209;
	{8'd139,8'd78} : s = 357;
	{8'd139,8'd79} : s = 355;
	{8'd139,8'd80} : s = 467;
	{8'd139,8'd81} : s = 348;
	{8'd139,8'd82} : s = 462;
	{8'd139,8'd83} : s = 461;
	{8'd139,8'd84} : s = 505;
	{8'd139,8'd85} : s = 84;
	{8'd139,8'd86} : s = 204;
	{8'd139,8'd87} : s = 202;
	{8'd139,8'd88} : s = 346;
	{8'd139,8'd89} : s = 201;
	{8'd139,8'd90} : s = 345;
	{8'd139,8'd91} : s = 342;
	{8'd139,8'd92} : s = 459;
	{8'd139,8'd93} : s = 198;
	{8'd139,8'd94} : s = 341;
	{8'd139,8'd95} : s = 339;
	{8'd139,8'd96} : s = 455;
	{8'd139,8'd97} : s = 334;
	{8'd139,8'd98} : s = 444;
	{8'd139,8'd99} : s = 442;
	{8'd139,8'd100} : s = 502;
	{8'd139,8'd101} : s = 197;
	{8'd139,8'd102} : s = 333;
	{8'd139,8'd103} : s = 331;
	{8'd139,8'd104} : s = 441;
	{8'd139,8'd105} : s = 327;
	{8'd139,8'd106} : s = 438;
	{8'd139,8'd107} : s = 437;
	{8'd139,8'd108} : s = 501;
	{8'd139,8'd109} : s = 316;
	{8'd139,8'd110} : s = 435;
	{8'd139,8'd111} : s = 430;
	{8'd139,8'd112} : s = 499;
	{8'd139,8'd113} : s = 429;
	{8'd139,8'd114} : s = 494;
	{8'd139,8'd115} : s = 493;
	{8'd139,8'd116} : s = 510;
	{8'd139,8'd117} : s = 1;
	{8'd139,8'd118} : s = 18;
	{8'd139,8'd119} : s = 17;
	{8'd139,8'd120} : s = 82;
	{8'd139,8'd121} : s = 12;
	{8'd139,8'd122} : s = 81;
	{8'd139,8'd123} : s = 76;
	{8'd139,8'd124} : s = 195;
	{8'd139,8'd125} : s = 10;
	{8'd139,8'd126} : s = 74;
	{8'd139,8'd127} : s = 73;
	{8'd139,8'd128} : s = 184;
	{8'd139,8'd129} : s = 70;
	{8'd139,8'd130} : s = 180;
	{8'd139,8'd131} : s = 178;
	{8'd139,8'd132} : s = 314;
	{8'd139,8'd133} : s = 9;
	{8'd139,8'd134} : s = 69;
	{8'd139,8'd135} : s = 67;
	{8'd139,8'd136} : s = 177;
	{8'd139,8'd137} : s = 56;
	{8'd139,8'd138} : s = 172;
	{8'd139,8'd139} : s = 170;
	{8'd139,8'd140} : s = 313;
	{8'd139,8'd141} : s = 52;
	{8'd139,8'd142} : s = 169;
	{8'd139,8'd143} : s = 166;
	{8'd139,8'd144} : s = 310;
	{8'd139,8'd145} : s = 165;
	{8'd139,8'd146} : s = 309;
	{8'd139,8'd147} : s = 307;
	{8'd139,8'd148} : s = 427;
	{8'd139,8'd149} : s = 6;
	{8'd139,8'd150} : s = 50;
	{8'd139,8'd151} : s = 49;
	{8'd139,8'd152} : s = 163;
	{8'd139,8'd153} : s = 44;
	{8'd139,8'd154} : s = 156;
	{8'd139,8'd155} : s = 154;
	{8'd139,8'd156} : s = 302;
	{8'd139,8'd157} : s = 42;
	{8'd139,8'd158} : s = 153;
	{8'd139,8'd159} : s = 150;
	{8'd139,8'd160} : s = 301;
	{8'd139,8'd161} : s = 149;
	{8'd139,8'd162} : s = 299;
	{8'd139,8'd163} : s = 295;
	{8'd139,8'd164} : s = 423;
	{8'd139,8'd165} : s = 41;
	{8'd139,8'd166} : s = 147;
	{8'd139,8'd167} : s = 142;
	{8'd139,8'd168} : s = 286;
	{8'd139,8'd169} : s = 141;
	{8'd139,8'd170} : s = 285;
	{8'd139,8'd171} : s = 283;
	{8'd139,8'd172} : s = 414;
	{8'd139,8'd173} : s = 139;
	{8'd139,8'd174} : s = 279;
	{8'd139,8'd175} : s = 271;
	{8'd139,8'd176} : s = 413;
	{8'd139,8'd177} : s = 248;
	{8'd139,8'd178} : s = 411;
	{8'd139,8'd179} : s = 407;
	{8'd139,8'd180} : s = 491;
	{8'd139,8'd181} : s = 5;
	{8'd139,8'd182} : s = 38;
	{8'd139,8'd183} : s = 37;
	{8'd139,8'd184} : s = 135;
	{8'd139,8'd185} : s = 35;
	{8'd139,8'd186} : s = 120;
	{8'd139,8'd187} : s = 116;
	{8'd139,8'd188} : s = 244;
	{8'd139,8'd189} : s = 28;
	{8'd139,8'd190} : s = 114;
	{8'd139,8'd191} : s = 113;
	{8'd139,8'd192} : s = 242;
	{8'd139,8'd193} : s = 108;
	{8'd139,8'd194} : s = 241;
	{8'd139,8'd195} : s = 236;
	{8'd139,8'd196} : s = 399;
	{8'd139,8'd197} : s = 26;
	{8'd139,8'd198} : s = 106;
	{8'd139,8'd199} : s = 105;
	{8'd139,8'd200} : s = 234;
	{8'd139,8'd201} : s = 102;
	{8'd139,8'd202} : s = 233;
	{8'd139,8'd203} : s = 230;
	{8'd139,8'd204} : s = 380;
	{8'd139,8'd205} : s = 101;
	{8'd139,8'd206} : s = 229;
	{8'd139,8'd207} : s = 227;
	{8'd139,8'd208} : s = 378;
	{8'd139,8'd209} : s = 220;
	{8'd139,8'd210} : s = 377;
	{8'd139,8'd211} : s = 374;
	{8'd139,8'd212} : s = 487;
	{8'd139,8'd213} : s = 25;
	{8'd139,8'd214} : s = 99;
	{8'd139,8'd215} : s = 92;
	{8'd139,8'd216} : s = 218;
	{8'd139,8'd217} : s = 90;
	{8'd139,8'd218} : s = 217;
	{8'd139,8'd219} : s = 214;
	{8'd139,8'd220} : s = 373;
	{8'd139,8'd221} : s = 89;
	{8'd139,8'd222} : s = 213;
	{8'd139,8'd223} : s = 211;
	{8'd139,8'd224} : s = 371;
	{8'd139,8'd225} : s = 206;
	{8'd139,8'd226} : s = 366;
	{8'd139,8'd227} : s = 365;
	{8'd139,8'd228} : s = 478;
	{8'd139,8'd229} : s = 86;
	{8'd139,8'd230} : s = 205;
	{8'd139,8'd231} : s = 203;
	{8'd139,8'd232} : s = 363;
	{8'd139,8'd233} : s = 199;
	{8'd139,8'd234} : s = 359;
	{8'd139,8'd235} : s = 350;
	{8'd139,8'd236} : s = 477;
	{8'd139,8'd237} : s = 188;
	{8'd139,8'd238} : s = 349;
	{8'd139,8'd239} : s = 347;
	{8'd139,8'd240} : s = 475;
	{8'd139,8'd241} : s = 343;
	{8'd139,8'd242} : s = 471;
	{8'd139,8'd243} : s = 463;
	{8'd139,8'd244} : s = 509;
	{8'd139,8'd245} : s = 3;
	{8'd139,8'd246} : s = 22;
	{8'd139,8'd247} : s = 21;
	{8'd139,8'd248} : s = 85;
	{8'd139,8'd249} : s = 19;
	{8'd139,8'd250} : s = 83;
	{8'd139,8'd251} : s = 78;
	{8'd139,8'd252} : s = 186;
	{8'd139,8'd253} : s = 14;
	{8'd139,8'd254} : s = 77;
	{8'd139,8'd255} : s = 75;
	{8'd140,8'd0} : s = 148;
	{8'd140,8'd1} : s = 308;
	{8'd140,8'd2} : s = 306;
	{8'd140,8'd3} : s = 425;
	{8'd140,8'd4} : s = 33;
	{8'd140,8'd5} : s = 146;
	{8'd140,8'd6} : s = 145;
	{8'd140,8'd7} : s = 305;
	{8'd140,8'd8} : s = 140;
	{8'd140,8'd9} : s = 300;
	{8'd140,8'd10} : s = 298;
	{8'd140,8'd11} : s = 422;
	{8'd140,8'd12} : s = 138;
	{8'd140,8'd13} : s = 297;
	{8'd140,8'd14} : s = 294;
	{8'd140,8'd15} : s = 421;
	{8'd140,8'd16} : s = 293;
	{8'd140,8'd17} : s = 419;
	{8'd140,8'd18} : s = 412;
	{8'd140,8'd19} : s = 486;
	{8'd140,8'd20} : s = 24;
	{8'd140,8'd21} : s = 137;
	{8'd140,8'd22} : s = 134;
	{8'd140,8'd23} : s = 291;
	{8'd140,8'd24} : s = 133;
	{8'd140,8'd25} : s = 284;
	{8'd140,8'd26} : s = 282;
	{8'd140,8'd27} : s = 410;
	{8'd140,8'd28} : s = 131;
	{8'd140,8'd29} : s = 281;
	{8'd140,8'd30} : s = 278;
	{8'd140,8'd31} : s = 409;
	{8'd140,8'd32} : s = 277;
	{8'd140,8'd33} : s = 406;
	{8'd140,8'd34} : s = 405;
	{8'd140,8'd35} : s = 485;
	{8'd140,8'd36} : s = 112;
	{8'd140,8'd37} : s = 275;
	{8'd140,8'd38} : s = 270;
	{8'd140,8'd39} : s = 403;
	{8'd140,8'd40} : s = 269;
	{8'd140,8'd41} : s = 398;
	{8'd140,8'd42} : s = 397;
	{8'd140,8'd43} : s = 483;
	{8'd140,8'd44} : s = 267;
	{8'd140,8'd45} : s = 395;
	{8'd140,8'd46} : s = 391;
	{8'd140,8'd47} : s = 476;
	{8'd140,8'd48} : s = 376;
	{8'd140,8'd49} : s = 474;
	{8'd140,8'd50} : s = 473;
	{8'd140,8'd51} : s = 506;
	{8'd140,8'd52} : s = 20;
	{8'd140,8'd53} : s = 104;
	{8'd140,8'd54} : s = 100;
	{8'd140,8'd55} : s = 263;
	{8'd140,8'd56} : s = 98;
	{8'd140,8'd57} : s = 240;
	{8'd140,8'd58} : s = 232;
	{8'd140,8'd59} : s = 372;
	{8'd140,8'd60} : s = 97;
	{8'd140,8'd61} : s = 228;
	{8'd140,8'd62} : s = 226;
	{8'd140,8'd63} : s = 370;
	{8'd140,8'd64} : s = 225;
	{8'd140,8'd65} : s = 369;
	{8'd140,8'd66} : s = 364;
	{8'd140,8'd67} : s = 470;
	{8'd140,8'd68} : s = 88;
	{8'd140,8'd69} : s = 216;
	{8'd140,8'd70} : s = 212;
	{8'd140,8'd71} : s = 362;
	{8'd140,8'd72} : s = 210;
	{8'd140,8'd73} : s = 361;
	{8'd140,8'd74} : s = 358;
	{8'd140,8'd75} : s = 469;
	{8'd140,8'd76} : s = 209;
	{8'd140,8'd77} : s = 357;
	{8'd140,8'd78} : s = 355;
	{8'd140,8'd79} : s = 467;
	{8'd140,8'd80} : s = 348;
	{8'd140,8'd81} : s = 462;
	{8'd140,8'd82} : s = 461;
	{8'd140,8'd83} : s = 505;
	{8'd140,8'd84} : s = 84;
	{8'd140,8'd85} : s = 204;
	{8'd140,8'd86} : s = 202;
	{8'd140,8'd87} : s = 346;
	{8'd140,8'd88} : s = 201;
	{8'd140,8'd89} : s = 345;
	{8'd140,8'd90} : s = 342;
	{8'd140,8'd91} : s = 459;
	{8'd140,8'd92} : s = 198;
	{8'd140,8'd93} : s = 341;
	{8'd140,8'd94} : s = 339;
	{8'd140,8'd95} : s = 455;
	{8'd140,8'd96} : s = 334;
	{8'd140,8'd97} : s = 444;
	{8'd140,8'd98} : s = 442;
	{8'd140,8'd99} : s = 502;
	{8'd140,8'd100} : s = 197;
	{8'd140,8'd101} : s = 333;
	{8'd140,8'd102} : s = 331;
	{8'd140,8'd103} : s = 441;
	{8'd140,8'd104} : s = 327;
	{8'd140,8'd105} : s = 438;
	{8'd140,8'd106} : s = 437;
	{8'd140,8'd107} : s = 501;
	{8'd140,8'd108} : s = 316;
	{8'd140,8'd109} : s = 435;
	{8'd140,8'd110} : s = 430;
	{8'd140,8'd111} : s = 499;
	{8'd140,8'd112} : s = 429;
	{8'd140,8'd113} : s = 494;
	{8'd140,8'd114} : s = 493;
	{8'd140,8'd115} : s = 510;
	{8'd140,8'd116} : s = 1;
	{8'd140,8'd117} : s = 18;
	{8'd140,8'd118} : s = 17;
	{8'd140,8'd119} : s = 82;
	{8'd140,8'd120} : s = 12;
	{8'd140,8'd121} : s = 81;
	{8'd140,8'd122} : s = 76;
	{8'd140,8'd123} : s = 195;
	{8'd140,8'd124} : s = 10;
	{8'd140,8'd125} : s = 74;
	{8'd140,8'd126} : s = 73;
	{8'd140,8'd127} : s = 184;
	{8'd140,8'd128} : s = 70;
	{8'd140,8'd129} : s = 180;
	{8'd140,8'd130} : s = 178;
	{8'd140,8'd131} : s = 314;
	{8'd140,8'd132} : s = 9;
	{8'd140,8'd133} : s = 69;
	{8'd140,8'd134} : s = 67;
	{8'd140,8'd135} : s = 177;
	{8'd140,8'd136} : s = 56;
	{8'd140,8'd137} : s = 172;
	{8'd140,8'd138} : s = 170;
	{8'd140,8'd139} : s = 313;
	{8'd140,8'd140} : s = 52;
	{8'd140,8'd141} : s = 169;
	{8'd140,8'd142} : s = 166;
	{8'd140,8'd143} : s = 310;
	{8'd140,8'd144} : s = 165;
	{8'd140,8'd145} : s = 309;
	{8'd140,8'd146} : s = 307;
	{8'd140,8'd147} : s = 427;
	{8'd140,8'd148} : s = 6;
	{8'd140,8'd149} : s = 50;
	{8'd140,8'd150} : s = 49;
	{8'd140,8'd151} : s = 163;
	{8'd140,8'd152} : s = 44;
	{8'd140,8'd153} : s = 156;
	{8'd140,8'd154} : s = 154;
	{8'd140,8'd155} : s = 302;
	{8'd140,8'd156} : s = 42;
	{8'd140,8'd157} : s = 153;
	{8'd140,8'd158} : s = 150;
	{8'd140,8'd159} : s = 301;
	{8'd140,8'd160} : s = 149;
	{8'd140,8'd161} : s = 299;
	{8'd140,8'd162} : s = 295;
	{8'd140,8'd163} : s = 423;
	{8'd140,8'd164} : s = 41;
	{8'd140,8'd165} : s = 147;
	{8'd140,8'd166} : s = 142;
	{8'd140,8'd167} : s = 286;
	{8'd140,8'd168} : s = 141;
	{8'd140,8'd169} : s = 285;
	{8'd140,8'd170} : s = 283;
	{8'd140,8'd171} : s = 414;
	{8'd140,8'd172} : s = 139;
	{8'd140,8'd173} : s = 279;
	{8'd140,8'd174} : s = 271;
	{8'd140,8'd175} : s = 413;
	{8'd140,8'd176} : s = 248;
	{8'd140,8'd177} : s = 411;
	{8'd140,8'd178} : s = 407;
	{8'd140,8'd179} : s = 491;
	{8'd140,8'd180} : s = 5;
	{8'd140,8'd181} : s = 38;
	{8'd140,8'd182} : s = 37;
	{8'd140,8'd183} : s = 135;
	{8'd140,8'd184} : s = 35;
	{8'd140,8'd185} : s = 120;
	{8'd140,8'd186} : s = 116;
	{8'd140,8'd187} : s = 244;
	{8'd140,8'd188} : s = 28;
	{8'd140,8'd189} : s = 114;
	{8'd140,8'd190} : s = 113;
	{8'd140,8'd191} : s = 242;
	{8'd140,8'd192} : s = 108;
	{8'd140,8'd193} : s = 241;
	{8'd140,8'd194} : s = 236;
	{8'd140,8'd195} : s = 399;
	{8'd140,8'd196} : s = 26;
	{8'd140,8'd197} : s = 106;
	{8'd140,8'd198} : s = 105;
	{8'd140,8'd199} : s = 234;
	{8'd140,8'd200} : s = 102;
	{8'd140,8'd201} : s = 233;
	{8'd140,8'd202} : s = 230;
	{8'd140,8'd203} : s = 380;
	{8'd140,8'd204} : s = 101;
	{8'd140,8'd205} : s = 229;
	{8'd140,8'd206} : s = 227;
	{8'd140,8'd207} : s = 378;
	{8'd140,8'd208} : s = 220;
	{8'd140,8'd209} : s = 377;
	{8'd140,8'd210} : s = 374;
	{8'd140,8'd211} : s = 487;
	{8'd140,8'd212} : s = 25;
	{8'd140,8'd213} : s = 99;
	{8'd140,8'd214} : s = 92;
	{8'd140,8'd215} : s = 218;
	{8'd140,8'd216} : s = 90;
	{8'd140,8'd217} : s = 217;
	{8'd140,8'd218} : s = 214;
	{8'd140,8'd219} : s = 373;
	{8'd140,8'd220} : s = 89;
	{8'd140,8'd221} : s = 213;
	{8'd140,8'd222} : s = 211;
	{8'd140,8'd223} : s = 371;
	{8'd140,8'd224} : s = 206;
	{8'd140,8'd225} : s = 366;
	{8'd140,8'd226} : s = 365;
	{8'd140,8'd227} : s = 478;
	{8'd140,8'd228} : s = 86;
	{8'd140,8'd229} : s = 205;
	{8'd140,8'd230} : s = 203;
	{8'd140,8'd231} : s = 363;
	{8'd140,8'd232} : s = 199;
	{8'd140,8'd233} : s = 359;
	{8'd140,8'd234} : s = 350;
	{8'd140,8'd235} : s = 477;
	{8'd140,8'd236} : s = 188;
	{8'd140,8'd237} : s = 349;
	{8'd140,8'd238} : s = 347;
	{8'd140,8'd239} : s = 475;
	{8'd140,8'd240} : s = 343;
	{8'd140,8'd241} : s = 471;
	{8'd140,8'd242} : s = 463;
	{8'd140,8'd243} : s = 509;
	{8'd140,8'd244} : s = 3;
	{8'd140,8'd245} : s = 22;
	{8'd140,8'd246} : s = 21;
	{8'd140,8'd247} : s = 85;
	{8'd140,8'd248} : s = 19;
	{8'd140,8'd249} : s = 83;
	{8'd140,8'd250} : s = 78;
	{8'd140,8'd251} : s = 186;
	{8'd140,8'd252} : s = 14;
	{8'd140,8'd253} : s = 77;
	{8'd140,8'd254} : s = 75;
	{8'd140,8'd255} : s = 185;
	{8'd141,8'd0} : s = 308;
	{8'd141,8'd1} : s = 306;
	{8'd141,8'd2} : s = 425;
	{8'd141,8'd3} : s = 33;
	{8'd141,8'd4} : s = 146;
	{8'd141,8'd5} : s = 145;
	{8'd141,8'd6} : s = 305;
	{8'd141,8'd7} : s = 140;
	{8'd141,8'd8} : s = 300;
	{8'd141,8'd9} : s = 298;
	{8'd141,8'd10} : s = 422;
	{8'd141,8'd11} : s = 138;
	{8'd141,8'd12} : s = 297;
	{8'd141,8'd13} : s = 294;
	{8'd141,8'd14} : s = 421;
	{8'd141,8'd15} : s = 293;
	{8'd141,8'd16} : s = 419;
	{8'd141,8'd17} : s = 412;
	{8'd141,8'd18} : s = 486;
	{8'd141,8'd19} : s = 24;
	{8'd141,8'd20} : s = 137;
	{8'd141,8'd21} : s = 134;
	{8'd141,8'd22} : s = 291;
	{8'd141,8'd23} : s = 133;
	{8'd141,8'd24} : s = 284;
	{8'd141,8'd25} : s = 282;
	{8'd141,8'd26} : s = 410;
	{8'd141,8'd27} : s = 131;
	{8'd141,8'd28} : s = 281;
	{8'd141,8'd29} : s = 278;
	{8'd141,8'd30} : s = 409;
	{8'd141,8'd31} : s = 277;
	{8'd141,8'd32} : s = 406;
	{8'd141,8'd33} : s = 405;
	{8'd141,8'd34} : s = 485;
	{8'd141,8'd35} : s = 112;
	{8'd141,8'd36} : s = 275;
	{8'd141,8'd37} : s = 270;
	{8'd141,8'd38} : s = 403;
	{8'd141,8'd39} : s = 269;
	{8'd141,8'd40} : s = 398;
	{8'd141,8'd41} : s = 397;
	{8'd141,8'd42} : s = 483;
	{8'd141,8'd43} : s = 267;
	{8'd141,8'd44} : s = 395;
	{8'd141,8'd45} : s = 391;
	{8'd141,8'd46} : s = 476;
	{8'd141,8'd47} : s = 376;
	{8'd141,8'd48} : s = 474;
	{8'd141,8'd49} : s = 473;
	{8'd141,8'd50} : s = 506;
	{8'd141,8'd51} : s = 20;
	{8'd141,8'd52} : s = 104;
	{8'd141,8'd53} : s = 100;
	{8'd141,8'd54} : s = 263;
	{8'd141,8'd55} : s = 98;
	{8'd141,8'd56} : s = 240;
	{8'd141,8'd57} : s = 232;
	{8'd141,8'd58} : s = 372;
	{8'd141,8'd59} : s = 97;
	{8'd141,8'd60} : s = 228;
	{8'd141,8'd61} : s = 226;
	{8'd141,8'd62} : s = 370;
	{8'd141,8'd63} : s = 225;
	{8'd141,8'd64} : s = 369;
	{8'd141,8'd65} : s = 364;
	{8'd141,8'd66} : s = 470;
	{8'd141,8'd67} : s = 88;
	{8'd141,8'd68} : s = 216;
	{8'd141,8'd69} : s = 212;
	{8'd141,8'd70} : s = 362;
	{8'd141,8'd71} : s = 210;
	{8'd141,8'd72} : s = 361;
	{8'd141,8'd73} : s = 358;
	{8'd141,8'd74} : s = 469;
	{8'd141,8'd75} : s = 209;
	{8'd141,8'd76} : s = 357;
	{8'd141,8'd77} : s = 355;
	{8'd141,8'd78} : s = 467;
	{8'd141,8'd79} : s = 348;
	{8'd141,8'd80} : s = 462;
	{8'd141,8'd81} : s = 461;
	{8'd141,8'd82} : s = 505;
	{8'd141,8'd83} : s = 84;
	{8'd141,8'd84} : s = 204;
	{8'd141,8'd85} : s = 202;
	{8'd141,8'd86} : s = 346;
	{8'd141,8'd87} : s = 201;
	{8'd141,8'd88} : s = 345;
	{8'd141,8'd89} : s = 342;
	{8'd141,8'd90} : s = 459;
	{8'd141,8'd91} : s = 198;
	{8'd141,8'd92} : s = 341;
	{8'd141,8'd93} : s = 339;
	{8'd141,8'd94} : s = 455;
	{8'd141,8'd95} : s = 334;
	{8'd141,8'd96} : s = 444;
	{8'd141,8'd97} : s = 442;
	{8'd141,8'd98} : s = 502;
	{8'd141,8'd99} : s = 197;
	{8'd141,8'd100} : s = 333;
	{8'd141,8'd101} : s = 331;
	{8'd141,8'd102} : s = 441;
	{8'd141,8'd103} : s = 327;
	{8'd141,8'd104} : s = 438;
	{8'd141,8'd105} : s = 437;
	{8'd141,8'd106} : s = 501;
	{8'd141,8'd107} : s = 316;
	{8'd141,8'd108} : s = 435;
	{8'd141,8'd109} : s = 430;
	{8'd141,8'd110} : s = 499;
	{8'd141,8'd111} : s = 429;
	{8'd141,8'd112} : s = 494;
	{8'd141,8'd113} : s = 493;
	{8'd141,8'd114} : s = 510;
	{8'd141,8'd115} : s = 1;
	{8'd141,8'd116} : s = 18;
	{8'd141,8'd117} : s = 17;
	{8'd141,8'd118} : s = 82;
	{8'd141,8'd119} : s = 12;
	{8'd141,8'd120} : s = 81;
	{8'd141,8'd121} : s = 76;
	{8'd141,8'd122} : s = 195;
	{8'd141,8'd123} : s = 10;
	{8'd141,8'd124} : s = 74;
	{8'd141,8'd125} : s = 73;
	{8'd141,8'd126} : s = 184;
	{8'd141,8'd127} : s = 70;
	{8'd141,8'd128} : s = 180;
	{8'd141,8'd129} : s = 178;
	{8'd141,8'd130} : s = 314;
	{8'd141,8'd131} : s = 9;
	{8'd141,8'd132} : s = 69;
	{8'd141,8'd133} : s = 67;
	{8'd141,8'd134} : s = 177;
	{8'd141,8'd135} : s = 56;
	{8'd141,8'd136} : s = 172;
	{8'd141,8'd137} : s = 170;
	{8'd141,8'd138} : s = 313;
	{8'd141,8'd139} : s = 52;
	{8'd141,8'd140} : s = 169;
	{8'd141,8'd141} : s = 166;
	{8'd141,8'd142} : s = 310;
	{8'd141,8'd143} : s = 165;
	{8'd141,8'd144} : s = 309;
	{8'd141,8'd145} : s = 307;
	{8'd141,8'd146} : s = 427;
	{8'd141,8'd147} : s = 6;
	{8'd141,8'd148} : s = 50;
	{8'd141,8'd149} : s = 49;
	{8'd141,8'd150} : s = 163;
	{8'd141,8'd151} : s = 44;
	{8'd141,8'd152} : s = 156;
	{8'd141,8'd153} : s = 154;
	{8'd141,8'd154} : s = 302;
	{8'd141,8'd155} : s = 42;
	{8'd141,8'd156} : s = 153;
	{8'd141,8'd157} : s = 150;
	{8'd141,8'd158} : s = 301;
	{8'd141,8'd159} : s = 149;
	{8'd141,8'd160} : s = 299;
	{8'd141,8'd161} : s = 295;
	{8'd141,8'd162} : s = 423;
	{8'd141,8'd163} : s = 41;
	{8'd141,8'd164} : s = 147;
	{8'd141,8'd165} : s = 142;
	{8'd141,8'd166} : s = 286;
	{8'd141,8'd167} : s = 141;
	{8'd141,8'd168} : s = 285;
	{8'd141,8'd169} : s = 283;
	{8'd141,8'd170} : s = 414;
	{8'd141,8'd171} : s = 139;
	{8'd141,8'd172} : s = 279;
	{8'd141,8'd173} : s = 271;
	{8'd141,8'd174} : s = 413;
	{8'd141,8'd175} : s = 248;
	{8'd141,8'd176} : s = 411;
	{8'd141,8'd177} : s = 407;
	{8'd141,8'd178} : s = 491;
	{8'd141,8'd179} : s = 5;
	{8'd141,8'd180} : s = 38;
	{8'd141,8'd181} : s = 37;
	{8'd141,8'd182} : s = 135;
	{8'd141,8'd183} : s = 35;
	{8'd141,8'd184} : s = 120;
	{8'd141,8'd185} : s = 116;
	{8'd141,8'd186} : s = 244;
	{8'd141,8'd187} : s = 28;
	{8'd141,8'd188} : s = 114;
	{8'd141,8'd189} : s = 113;
	{8'd141,8'd190} : s = 242;
	{8'd141,8'd191} : s = 108;
	{8'd141,8'd192} : s = 241;
	{8'd141,8'd193} : s = 236;
	{8'd141,8'd194} : s = 399;
	{8'd141,8'd195} : s = 26;
	{8'd141,8'd196} : s = 106;
	{8'd141,8'd197} : s = 105;
	{8'd141,8'd198} : s = 234;
	{8'd141,8'd199} : s = 102;
	{8'd141,8'd200} : s = 233;
	{8'd141,8'd201} : s = 230;
	{8'd141,8'd202} : s = 380;
	{8'd141,8'd203} : s = 101;
	{8'd141,8'd204} : s = 229;
	{8'd141,8'd205} : s = 227;
	{8'd141,8'd206} : s = 378;
	{8'd141,8'd207} : s = 220;
	{8'd141,8'd208} : s = 377;
	{8'd141,8'd209} : s = 374;
	{8'd141,8'd210} : s = 487;
	{8'd141,8'd211} : s = 25;
	{8'd141,8'd212} : s = 99;
	{8'd141,8'd213} : s = 92;
	{8'd141,8'd214} : s = 218;
	{8'd141,8'd215} : s = 90;
	{8'd141,8'd216} : s = 217;
	{8'd141,8'd217} : s = 214;
	{8'd141,8'd218} : s = 373;
	{8'd141,8'd219} : s = 89;
	{8'd141,8'd220} : s = 213;
	{8'd141,8'd221} : s = 211;
	{8'd141,8'd222} : s = 371;
	{8'd141,8'd223} : s = 206;
	{8'd141,8'd224} : s = 366;
	{8'd141,8'd225} : s = 365;
	{8'd141,8'd226} : s = 478;
	{8'd141,8'd227} : s = 86;
	{8'd141,8'd228} : s = 205;
	{8'd141,8'd229} : s = 203;
	{8'd141,8'd230} : s = 363;
	{8'd141,8'd231} : s = 199;
	{8'd141,8'd232} : s = 359;
	{8'd141,8'd233} : s = 350;
	{8'd141,8'd234} : s = 477;
	{8'd141,8'd235} : s = 188;
	{8'd141,8'd236} : s = 349;
	{8'd141,8'd237} : s = 347;
	{8'd141,8'd238} : s = 475;
	{8'd141,8'd239} : s = 343;
	{8'd141,8'd240} : s = 471;
	{8'd141,8'd241} : s = 463;
	{8'd141,8'd242} : s = 509;
	{8'd141,8'd243} : s = 3;
	{8'd141,8'd244} : s = 22;
	{8'd141,8'd245} : s = 21;
	{8'd141,8'd246} : s = 85;
	{8'd141,8'd247} : s = 19;
	{8'd141,8'd248} : s = 83;
	{8'd141,8'd249} : s = 78;
	{8'd141,8'd250} : s = 186;
	{8'd141,8'd251} : s = 14;
	{8'd141,8'd252} : s = 77;
	{8'd141,8'd253} : s = 75;
	{8'd141,8'd254} : s = 185;
	{8'd141,8'd255} : s = 71;
	{8'd142,8'd0} : s = 306;
	{8'd142,8'd1} : s = 425;
	{8'd142,8'd2} : s = 33;
	{8'd142,8'd3} : s = 146;
	{8'd142,8'd4} : s = 145;
	{8'd142,8'd5} : s = 305;
	{8'd142,8'd6} : s = 140;
	{8'd142,8'd7} : s = 300;
	{8'd142,8'd8} : s = 298;
	{8'd142,8'd9} : s = 422;
	{8'd142,8'd10} : s = 138;
	{8'd142,8'd11} : s = 297;
	{8'd142,8'd12} : s = 294;
	{8'd142,8'd13} : s = 421;
	{8'd142,8'd14} : s = 293;
	{8'd142,8'd15} : s = 419;
	{8'd142,8'd16} : s = 412;
	{8'd142,8'd17} : s = 486;
	{8'd142,8'd18} : s = 24;
	{8'd142,8'd19} : s = 137;
	{8'd142,8'd20} : s = 134;
	{8'd142,8'd21} : s = 291;
	{8'd142,8'd22} : s = 133;
	{8'd142,8'd23} : s = 284;
	{8'd142,8'd24} : s = 282;
	{8'd142,8'd25} : s = 410;
	{8'd142,8'd26} : s = 131;
	{8'd142,8'd27} : s = 281;
	{8'd142,8'd28} : s = 278;
	{8'd142,8'd29} : s = 409;
	{8'd142,8'd30} : s = 277;
	{8'd142,8'd31} : s = 406;
	{8'd142,8'd32} : s = 405;
	{8'd142,8'd33} : s = 485;
	{8'd142,8'd34} : s = 112;
	{8'd142,8'd35} : s = 275;
	{8'd142,8'd36} : s = 270;
	{8'd142,8'd37} : s = 403;
	{8'd142,8'd38} : s = 269;
	{8'd142,8'd39} : s = 398;
	{8'd142,8'd40} : s = 397;
	{8'd142,8'd41} : s = 483;
	{8'd142,8'd42} : s = 267;
	{8'd142,8'd43} : s = 395;
	{8'd142,8'd44} : s = 391;
	{8'd142,8'd45} : s = 476;
	{8'd142,8'd46} : s = 376;
	{8'd142,8'd47} : s = 474;
	{8'd142,8'd48} : s = 473;
	{8'd142,8'd49} : s = 506;
	{8'd142,8'd50} : s = 20;
	{8'd142,8'd51} : s = 104;
	{8'd142,8'd52} : s = 100;
	{8'd142,8'd53} : s = 263;
	{8'd142,8'd54} : s = 98;
	{8'd142,8'd55} : s = 240;
	{8'd142,8'd56} : s = 232;
	{8'd142,8'd57} : s = 372;
	{8'd142,8'd58} : s = 97;
	{8'd142,8'd59} : s = 228;
	{8'd142,8'd60} : s = 226;
	{8'd142,8'd61} : s = 370;
	{8'd142,8'd62} : s = 225;
	{8'd142,8'd63} : s = 369;
	{8'd142,8'd64} : s = 364;
	{8'd142,8'd65} : s = 470;
	{8'd142,8'd66} : s = 88;
	{8'd142,8'd67} : s = 216;
	{8'd142,8'd68} : s = 212;
	{8'd142,8'd69} : s = 362;
	{8'd142,8'd70} : s = 210;
	{8'd142,8'd71} : s = 361;
	{8'd142,8'd72} : s = 358;
	{8'd142,8'd73} : s = 469;
	{8'd142,8'd74} : s = 209;
	{8'd142,8'd75} : s = 357;
	{8'd142,8'd76} : s = 355;
	{8'd142,8'd77} : s = 467;
	{8'd142,8'd78} : s = 348;
	{8'd142,8'd79} : s = 462;
	{8'd142,8'd80} : s = 461;
	{8'd142,8'd81} : s = 505;
	{8'd142,8'd82} : s = 84;
	{8'd142,8'd83} : s = 204;
	{8'd142,8'd84} : s = 202;
	{8'd142,8'd85} : s = 346;
	{8'd142,8'd86} : s = 201;
	{8'd142,8'd87} : s = 345;
	{8'd142,8'd88} : s = 342;
	{8'd142,8'd89} : s = 459;
	{8'd142,8'd90} : s = 198;
	{8'd142,8'd91} : s = 341;
	{8'd142,8'd92} : s = 339;
	{8'd142,8'd93} : s = 455;
	{8'd142,8'd94} : s = 334;
	{8'd142,8'd95} : s = 444;
	{8'd142,8'd96} : s = 442;
	{8'd142,8'd97} : s = 502;
	{8'd142,8'd98} : s = 197;
	{8'd142,8'd99} : s = 333;
	{8'd142,8'd100} : s = 331;
	{8'd142,8'd101} : s = 441;
	{8'd142,8'd102} : s = 327;
	{8'd142,8'd103} : s = 438;
	{8'd142,8'd104} : s = 437;
	{8'd142,8'd105} : s = 501;
	{8'd142,8'd106} : s = 316;
	{8'd142,8'd107} : s = 435;
	{8'd142,8'd108} : s = 430;
	{8'd142,8'd109} : s = 499;
	{8'd142,8'd110} : s = 429;
	{8'd142,8'd111} : s = 494;
	{8'd142,8'd112} : s = 493;
	{8'd142,8'd113} : s = 510;
	{8'd142,8'd114} : s = 1;
	{8'd142,8'd115} : s = 18;
	{8'd142,8'd116} : s = 17;
	{8'd142,8'd117} : s = 82;
	{8'd142,8'd118} : s = 12;
	{8'd142,8'd119} : s = 81;
	{8'd142,8'd120} : s = 76;
	{8'd142,8'd121} : s = 195;
	{8'd142,8'd122} : s = 10;
	{8'd142,8'd123} : s = 74;
	{8'd142,8'd124} : s = 73;
	{8'd142,8'd125} : s = 184;
	{8'd142,8'd126} : s = 70;
	{8'd142,8'd127} : s = 180;
	{8'd142,8'd128} : s = 178;
	{8'd142,8'd129} : s = 314;
	{8'd142,8'd130} : s = 9;
	{8'd142,8'd131} : s = 69;
	{8'd142,8'd132} : s = 67;
	{8'd142,8'd133} : s = 177;
	{8'd142,8'd134} : s = 56;
	{8'd142,8'd135} : s = 172;
	{8'd142,8'd136} : s = 170;
	{8'd142,8'd137} : s = 313;
	{8'd142,8'd138} : s = 52;
	{8'd142,8'd139} : s = 169;
	{8'd142,8'd140} : s = 166;
	{8'd142,8'd141} : s = 310;
	{8'd142,8'd142} : s = 165;
	{8'd142,8'd143} : s = 309;
	{8'd142,8'd144} : s = 307;
	{8'd142,8'd145} : s = 427;
	{8'd142,8'd146} : s = 6;
	{8'd142,8'd147} : s = 50;
	{8'd142,8'd148} : s = 49;
	{8'd142,8'd149} : s = 163;
	{8'd142,8'd150} : s = 44;
	{8'd142,8'd151} : s = 156;
	{8'd142,8'd152} : s = 154;
	{8'd142,8'd153} : s = 302;
	{8'd142,8'd154} : s = 42;
	{8'd142,8'd155} : s = 153;
	{8'd142,8'd156} : s = 150;
	{8'd142,8'd157} : s = 301;
	{8'd142,8'd158} : s = 149;
	{8'd142,8'd159} : s = 299;
	{8'd142,8'd160} : s = 295;
	{8'd142,8'd161} : s = 423;
	{8'd142,8'd162} : s = 41;
	{8'd142,8'd163} : s = 147;
	{8'd142,8'd164} : s = 142;
	{8'd142,8'd165} : s = 286;
	{8'd142,8'd166} : s = 141;
	{8'd142,8'd167} : s = 285;
	{8'd142,8'd168} : s = 283;
	{8'd142,8'd169} : s = 414;
	{8'd142,8'd170} : s = 139;
	{8'd142,8'd171} : s = 279;
	{8'd142,8'd172} : s = 271;
	{8'd142,8'd173} : s = 413;
	{8'd142,8'd174} : s = 248;
	{8'd142,8'd175} : s = 411;
	{8'd142,8'd176} : s = 407;
	{8'd142,8'd177} : s = 491;
	{8'd142,8'd178} : s = 5;
	{8'd142,8'd179} : s = 38;
	{8'd142,8'd180} : s = 37;
	{8'd142,8'd181} : s = 135;
	{8'd142,8'd182} : s = 35;
	{8'd142,8'd183} : s = 120;
	{8'd142,8'd184} : s = 116;
	{8'd142,8'd185} : s = 244;
	{8'd142,8'd186} : s = 28;
	{8'd142,8'd187} : s = 114;
	{8'd142,8'd188} : s = 113;
	{8'd142,8'd189} : s = 242;
	{8'd142,8'd190} : s = 108;
	{8'd142,8'd191} : s = 241;
	{8'd142,8'd192} : s = 236;
	{8'd142,8'd193} : s = 399;
	{8'd142,8'd194} : s = 26;
	{8'd142,8'd195} : s = 106;
	{8'd142,8'd196} : s = 105;
	{8'd142,8'd197} : s = 234;
	{8'd142,8'd198} : s = 102;
	{8'd142,8'd199} : s = 233;
	{8'd142,8'd200} : s = 230;
	{8'd142,8'd201} : s = 380;
	{8'd142,8'd202} : s = 101;
	{8'd142,8'd203} : s = 229;
	{8'd142,8'd204} : s = 227;
	{8'd142,8'd205} : s = 378;
	{8'd142,8'd206} : s = 220;
	{8'd142,8'd207} : s = 377;
	{8'd142,8'd208} : s = 374;
	{8'd142,8'd209} : s = 487;
	{8'd142,8'd210} : s = 25;
	{8'd142,8'd211} : s = 99;
	{8'd142,8'd212} : s = 92;
	{8'd142,8'd213} : s = 218;
	{8'd142,8'd214} : s = 90;
	{8'd142,8'd215} : s = 217;
	{8'd142,8'd216} : s = 214;
	{8'd142,8'd217} : s = 373;
	{8'd142,8'd218} : s = 89;
	{8'd142,8'd219} : s = 213;
	{8'd142,8'd220} : s = 211;
	{8'd142,8'd221} : s = 371;
	{8'd142,8'd222} : s = 206;
	{8'd142,8'd223} : s = 366;
	{8'd142,8'd224} : s = 365;
	{8'd142,8'd225} : s = 478;
	{8'd142,8'd226} : s = 86;
	{8'd142,8'd227} : s = 205;
	{8'd142,8'd228} : s = 203;
	{8'd142,8'd229} : s = 363;
	{8'd142,8'd230} : s = 199;
	{8'd142,8'd231} : s = 359;
	{8'd142,8'd232} : s = 350;
	{8'd142,8'd233} : s = 477;
	{8'd142,8'd234} : s = 188;
	{8'd142,8'd235} : s = 349;
	{8'd142,8'd236} : s = 347;
	{8'd142,8'd237} : s = 475;
	{8'd142,8'd238} : s = 343;
	{8'd142,8'd239} : s = 471;
	{8'd142,8'd240} : s = 463;
	{8'd142,8'd241} : s = 509;
	{8'd142,8'd242} : s = 3;
	{8'd142,8'd243} : s = 22;
	{8'd142,8'd244} : s = 21;
	{8'd142,8'd245} : s = 85;
	{8'd142,8'd246} : s = 19;
	{8'd142,8'd247} : s = 83;
	{8'd142,8'd248} : s = 78;
	{8'd142,8'd249} : s = 186;
	{8'd142,8'd250} : s = 14;
	{8'd142,8'd251} : s = 77;
	{8'd142,8'd252} : s = 75;
	{8'd142,8'd253} : s = 185;
	{8'd142,8'd254} : s = 71;
	{8'd142,8'd255} : s = 182;
	{8'd143,8'd0} : s = 425;
	{8'd143,8'd1} : s = 33;
	{8'd143,8'd2} : s = 146;
	{8'd143,8'd3} : s = 145;
	{8'd143,8'd4} : s = 305;
	{8'd143,8'd5} : s = 140;
	{8'd143,8'd6} : s = 300;
	{8'd143,8'd7} : s = 298;
	{8'd143,8'd8} : s = 422;
	{8'd143,8'd9} : s = 138;
	{8'd143,8'd10} : s = 297;
	{8'd143,8'd11} : s = 294;
	{8'd143,8'd12} : s = 421;
	{8'd143,8'd13} : s = 293;
	{8'd143,8'd14} : s = 419;
	{8'd143,8'd15} : s = 412;
	{8'd143,8'd16} : s = 486;
	{8'd143,8'd17} : s = 24;
	{8'd143,8'd18} : s = 137;
	{8'd143,8'd19} : s = 134;
	{8'd143,8'd20} : s = 291;
	{8'd143,8'd21} : s = 133;
	{8'd143,8'd22} : s = 284;
	{8'd143,8'd23} : s = 282;
	{8'd143,8'd24} : s = 410;
	{8'd143,8'd25} : s = 131;
	{8'd143,8'd26} : s = 281;
	{8'd143,8'd27} : s = 278;
	{8'd143,8'd28} : s = 409;
	{8'd143,8'd29} : s = 277;
	{8'd143,8'd30} : s = 406;
	{8'd143,8'd31} : s = 405;
	{8'd143,8'd32} : s = 485;
	{8'd143,8'd33} : s = 112;
	{8'd143,8'd34} : s = 275;
	{8'd143,8'd35} : s = 270;
	{8'd143,8'd36} : s = 403;
	{8'd143,8'd37} : s = 269;
	{8'd143,8'd38} : s = 398;
	{8'd143,8'd39} : s = 397;
	{8'd143,8'd40} : s = 483;
	{8'd143,8'd41} : s = 267;
	{8'd143,8'd42} : s = 395;
	{8'd143,8'd43} : s = 391;
	{8'd143,8'd44} : s = 476;
	{8'd143,8'd45} : s = 376;
	{8'd143,8'd46} : s = 474;
	{8'd143,8'd47} : s = 473;
	{8'd143,8'd48} : s = 506;
	{8'd143,8'd49} : s = 20;
	{8'd143,8'd50} : s = 104;
	{8'd143,8'd51} : s = 100;
	{8'd143,8'd52} : s = 263;
	{8'd143,8'd53} : s = 98;
	{8'd143,8'd54} : s = 240;
	{8'd143,8'd55} : s = 232;
	{8'd143,8'd56} : s = 372;
	{8'd143,8'd57} : s = 97;
	{8'd143,8'd58} : s = 228;
	{8'd143,8'd59} : s = 226;
	{8'd143,8'd60} : s = 370;
	{8'd143,8'd61} : s = 225;
	{8'd143,8'd62} : s = 369;
	{8'd143,8'd63} : s = 364;
	{8'd143,8'd64} : s = 470;
	{8'd143,8'd65} : s = 88;
	{8'd143,8'd66} : s = 216;
	{8'd143,8'd67} : s = 212;
	{8'd143,8'd68} : s = 362;
	{8'd143,8'd69} : s = 210;
	{8'd143,8'd70} : s = 361;
	{8'd143,8'd71} : s = 358;
	{8'd143,8'd72} : s = 469;
	{8'd143,8'd73} : s = 209;
	{8'd143,8'd74} : s = 357;
	{8'd143,8'd75} : s = 355;
	{8'd143,8'd76} : s = 467;
	{8'd143,8'd77} : s = 348;
	{8'd143,8'd78} : s = 462;
	{8'd143,8'd79} : s = 461;
	{8'd143,8'd80} : s = 505;
	{8'd143,8'd81} : s = 84;
	{8'd143,8'd82} : s = 204;
	{8'd143,8'd83} : s = 202;
	{8'd143,8'd84} : s = 346;
	{8'd143,8'd85} : s = 201;
	{8'd143,8'd86} : s = 345;
	{8'd143,8'd87} : s = 342;
	{8'd143,8'd88} : s = 459;
	{8'd143,8'd89} : s = 198;
	{8'd143,8'd90} : s = 341;
	{8'd143,8'd91} : s = 339;
	{8'd143,8'd92} : s = 455;
	{8'd143,8'd93} : s = 334;
	{8'd143,8'd94} : s = 444;
	{8'd143,8'd95} : s = 442;
	{8'd143,8'd96} : s = 502;
	{8'd143,8'd97} : s = 197;
	{8'd143,8'd98} : s = 333;
	{8'd143,8'd99} : s = 331;
	{8'd143,8'd100} : s = 441;
	{8'd143,8'd101} : s = 327;
	{8'd143,8'd102} : s = 438;
	{8'd143,8'd103} : s = 437;
	{8'd143,8'd104} : s = 501;
	{8'd143,8'd105} : s = 316;
	{8'd143,8'd106} : s = 435;
	{8'd143,8'd107} : s = 430;
	{8'd143,8'd108} : s = 499;
	{8'd143,8'd109} : s = 429;
	{8'd143,8'd110} : s = 494;
	{8'd143,8'd111} : s = 493;
	{8'd143,8'd112} : s = 510;
	{8'd143,8'd113} : s = 1;
	{8'd143,8'd114} : s = 18;
	{8'd143,8'd115} : s = 17;
	{8'd143,8'd116} : s = 82;
	{8'd143,8'd117} : s = 12;
	{8'd143,8'd118} : s = 81;
	{8'd143,8'd119} : s = 76;
	{8'd143,8'd120} : s = 195;
	{8'd143,8'd121} : s = 10;
	{8'd143,8'd122} : s = 74;
	{8'd143,8'd123} : s = 73;
	{8'd143,8'd124} : s = 184;
	{8'd143,8'd125} : s = 70;
	{8'd143,8'd126} : s = 180;
	{8'd143,8'd127} : s = 178;
	{8'd143,8'd128} : s = 314;
	{8'd143,8'd129} : s = 9;
	{8'd143,8'd130} : s = 69;
	{8'd143,8'd131} : s = 67;
	{8'd143,8'd132} : s = 177;
	{8'd143,8'd133} : s = 56;
	{8'd143,8'd134} : s = 172;
	{8'd143,8'd135} : s = 170;
	{8'd143,8'd136} : s = 313;
	{8'd143,8'd137} : s = 52;
	{8'd143,8'd138} : s = 169;
	{8'd143,8'd139} : s = 166;
	{8'd143,8'd140} : s = 310;
	{8'd143,8'd141} : s = 165;
	{8'd143,8'd142} : s = 309;
	{8'd143,8'd143} : s = 307;
	{8'd143,8'd144} : s = 427;
	{8'd143,8'd145} : s = 6;
	{8'd143,8'd146} : s = 50;
	{8'd143,8'd147} : s = 49;
	{8'd143,8'd148} : s = 163;
	{8'd143,8'd149} : s = 44;
	{8'd143,8'd150} : s = 156;
	{8'd143,8'd151} : s = 154;
	{8'd143,8'd152} : s = 302;
	{8'd143,8'd153} : s = 42;
	{8'd143,8'd154} : s = 153;
	{8'd143,8'd155} : s = 150;
	{8'd143,8'd156} : s = 301;
	{8'd143,8'd157} : s = 149;
	{8'd143,8'd158} : s = 299;
	{8'd143,8'd159} : s = 295;
	{8'd143,8'd160} : s = 423;
	{8'd143,8'd161} : s = 41;
	{8'd143,8'd162} : s = 147;
	{8'd143,8'd163} : s = 142;
	{8'd143,8'd164} : s = 286;
	{8'd143,8'd165} : s = 141;
	{8'd143,8'd166} : s = 285;
	{8'd143,8'd167} : s = 283;
	{8'd143,8'd168} : s = 414;
	{8'd143,8'd169} : s = 139;
	{8'd143,8'd170} : s = 279;
	{8'd143,8'd171} : s = 271;
	{8'd143,8'd172} : s = 413;
	{8'd143,8'd173} : s = 248;
	{8'd143,8'd174} : s = 411;
	{8'd143,8'd175} : s = 407;
	{8'd143,8'd176} : s = 491;
	{8'd143,8'd177} : s = 5;
	{8'd143,8'd178} : s = 38;
	{8'd143,8'd179} : s = 37;
	{8'd143,8'd180} : s = 135;
	{8'd143,8'd181} : s = 35;
	{8'd143,8'd182} : s = 120;
	{8'd143,8'd183} : s = 116;
	{8'd143,8'd184} : s = 244;
	{8'd143,8'd185} : s = 28;
	{8'd143,8'd186} : s = 114;
	{8'd143,8'd187} : s = 113;
	{8'd143,8'd188} : s = 242;
	{8'd143,8'd189} : s = 108;
	{8'd143,8'd190} : s = 241;
	{8'd143,8'd191} : s = 236;
	{8'd143,8'd192} : s = 399;
	{8'd143,8'd193} : s = 26;
	{8'd143,8'd194} : s = 106;
	{8'd143,8'd195} : s = 105;
	{8'd143,8'd196} : s = 234;
	{8'd143,8'd197} : s = 102;
	{8'd143,8'd198} : s = 233;
	{8'd143,8'd199} : s = 230;
	{8'd143,8'd200} : s = 380;
	{8'd143,8'd201} : s = 101;
	{8'd143,8'd202} : s = 229;
	{8'd143,8'd203} : s = 227;
	{8'd143,8'd204} : s = 378;
	{8'd143,8'd205} : s = 220;
	{8'd143,8'd206} : s = 377;
	{8'd143,8'd207} : s = 374;
	{8'd143,8'd208} : s = 487;
	{8'd143,8'd209} : s = 25;
	{8'd143,8'd210} : s = 99;
	{8'd143,8'd211} : s = 92;
	{8'd143,8'd212} : s = 218;
	{8'd143,8'd213} : s = 90;
	{8'd143,8'd214} : s = 217;
	{8'd143,8'd215} : s = 214;
	{8'd143,8'd216} : s = 373;
	{8'd143,8'd217} : s = 89;
	{8'd143,8'd218} : s = 213;
	{8'd143,8'd219} : s = 211;
	{8'd143,8'd220} : s = 371;
	{8'd143,8'd221} : s = 206;
	{8'd143,8'd222} : s = 366;
	{8'd143,8'd223} : s = 365;
	{8'd143,8'd224} : s = 478;
	{8'd143,8'd225} : s = 86;
	{8'd143,8'd226} : s = 205;
	{8'd143,8'd227} : s = 203;
	{8'd143,8'd228} : s = 363;
	{8'd143,8'd229} : s = 199;
	{8'd143,8'd230} : s = 359;
	{8'd143,8'd231} : s = 350;
	{8'd143,8'd232} : s = 477;
	{8'd143,8'd233} : s = 188;
	{8'd143,8'd234} : s = 349;
	{8'd143,8'd235} : s = 347;
	{8'd143,8'd236} : s = 475;
	{8'd143,8'd237} : s = 343;
	{8'd143,8'd238} : s = 471;
	{8'd143,8'd239} : s = 463;
	{8'd143,8'd240} : s = 509;
	{8'd143,8'd241} : s = 3;
	{8'd143,8'd242} : s = 22;
	{8'd143,8'd243} : s = 21;
	{8'd143,8'd244} : s = 85;
	{8'd143,8'd245} : s = 19;
	{8'd143,8'd246} : s = 83;
	{8'd143,8'd247} : s = 78;
	{8'd143,8'd248} : s = 186;
	{8'd143,8'd249} : s = 14;
	{8'd143,8'd250} : s = 77;
	{8'd143,8'd251} : s = 75;
	{8'd143,8'd252} : s = 185;
	{8'd143,8'd253} : s = 71;
	{8'd143,8'd254} : s = 182;
	{8'd143,8'd255} : s = 181;
	{8'd144,8'd0} : s = 33;
	{8'd144,8'd1} : s = 146;
	{8'd144,8'd2} : s = 145;
	{8'd144,8'd3} : s = 305;
	{8'd144,8'd4} : s = 140;
	{8'd144,8'd5} : s = 300;
	{8'd144,8'd6} : s = 298;
	{8'd144,8'd7} : s = 422;
	{8'd144,8'd8} : s = 138;
	{8'd144,8'd9} : s = 297;
	{8'd144,8'd10} : s = 294;
	{8'd144,8'd11} : s = 421;
	{8'd144,8'd12} : s = 293;
	{8'd144,8'd13} : s = 419;
	{8'd144,8'd14} : s = 412;
	{8'd144,8'd15} : s = 486;
	{8'd144,8'd16} : s = 24;
	{8'd144,8'd17} : s = 137;
	{8'd144,8'd18} : s = 134;
	{8'd144,8'd19} : s = 291;
	{8'd144,8'd20} : s = 133;
	{8'd144,8'd21} : s = 284;
	{8'd144,8'd22} : s = 282;
	{8'd144,8'd23} : s = 410;
	{8'd144,8'd24} : s = 131;
	{8'd144,8'd25} : s = 281;
	{8'd144,8'd26} : s = 278;
	{8'd144,8'd27} : s = 409;
	{8'd144,8'd28} : s = 277;
	{8'd144,8'd29} : s = 406;
	{8'd144,8'd30} : s = 405;
	{8'd144,8'd31} : s = 485;
	{8'd144,8'd32} : s = 112;
	{8'd144,8'd33} : s = 275;
	{8'd144,8'd34} : s = 270;
	{8'd144,8'd35} : s = 403;
	{8'd144,8'd36} : s = 269;
	{8'd144,8'd37} : s = 398;
	{8'd144,8'd38} : s = 397;
	{8'd144,8'd39} : s = 483;
	{8'd144,8'd40} : s = 267;
	{8'd144,8'd41} : s = 395;
	{8'd144,8'd42} : s = 391;
	{8'd144,8'd43} : s = 476;
	{8'd144,8'd44} : s = 376;
	{8'd144,8'd45} : s = 474;
	{8'd144,8'd46} : s = 473;
	{8'd144,8'd47} : s = 506;
	{8'd144,8'd48} : s = 20;
	{8'd144,8'd49} : s = 104;
	{8'd144,8'd50} : s = 100;
	{8'd144,8'd51} : s = 263;
	{8'd144,8'd52} : s = 98;
	{8'd144,8'd53} : s = 240;
	{8'd144,8'd54} : s = 232;
	{8'd144,8'd55} : s = 372;
	{8'd144,8'd56} : s = 97;
	{8'd144,8'd57} : s = 228;
	{8'd144,8'd58} : s = 226;
	{8'd144,8'd59} : s = 370;
	{8'd144,8'd60} : s = 225;
	{8'd144,8'd61} : s = 369;
	{8'd144,8'd62} : s = 364;
	{8'd144,8'd63} : s = 470;
	{8'd144,8'd64} : s = 88;
	{8'd144,8'd65} : s = 216;
	{8'd144,8'd66} : s = 212;
	{8'd144,8'd67} : s = 362;
	{8'd144,8'd68} : s = 210;
	{8'd144,8'd69} : s = 361;
	{8'd144,8'd70} : s = 358;
	{8'd144,8'd71} : s = 469;
	{8'd144,8'd72} : s = 209;
	{8'd144,8'd73} : s = 357;
	{8'd144,8'd74} : s = 355;
	{8'd144,8'd75} : s = 467;
	{8'd144,8'd76} : s = 348;
	{8'd144,8'd77} : s = 462;
	{8'd144,8'd78} : s = 461;
	{8'd144,8'd79} : s = 505;
	{8'd144,8'd80} : s = 84;
	{8'd144,8'd81} : s = 204;
	{8'd144,8'd82} : s = 202;
	{8'd144,8'd83} : s = 346;
	{8'd144,8'd84} : s = 201;
	{8'd144,8'd85} : s = 345;
	{8'd144,8'd86} : s = 342;
	{8'd144,8'd87} : s = 459;
	{8'd144,8'd88} : s = 198;
	{8'd144,8'd89} : s = 341;
	{8'd144,8'd90} : s = 339;
	{8'd144,8'd91} : s = 455;
	{8'd144,8'd92} : s = 334;
	{8'd144,8'd93} : s = 444;
	{8'd144,8'd94} : s = 442;
	{8'd144,8'd95} : s = 502;
	{8'd144,8'd96} : s = 197;
	{8'd144,8'd97} : s = 333;
	{8'd144,8'd98} : s = 331;
	{8'd144,8'd99} : s = 441;
	{8'd144,8'd100} : s = 327;
	{8'd144,8'd101} : s = 438;
	{8'd144,8'd102} : s = 437;
	{8'd144,8'd103} : s = 501;
	{8'd144,8'd104} : s = 316;
	{8'd144,8'd105} : s = 435;
	{8'd144,8'd106} : s = 430;
	{8'd144,8'd107} : s = 499;
	{8'd144,8'd108} : s = 429;
	{8'd144,8'd109} : s = 494;
	{8'd144,8'd110} : s = 493;
	{8'd144,8'd111} : s = 510;
	{8'd144,8'd112} : s = 1;
	{8'd144,8'd113} : s = 18;
	{8'd144,8'd114} : s = 17;
	{8'd144,8'd115} : s = 82;
	{8'd144,8'd116} : s = 12;
	{8'd144,8'd117} : s = 81;
	{8'd144,8'd118} : s = 76;
	{8'd144,8'd119} : s = 195;
	{8'd144,8'd120} : s = 10;
	{8'd144,8'd121} : s = 74;
	{8'd144,8'd122} : s = 73;
	{8'd144,8'd123} : s = 184;
	{8'd144,8'd124} : s = 70;
	{8'd144,8'd125} : s = 180;
	{8'd144,8'd126} : s = 178;
	{8'd144,8'd127} : s = 314;
	{8'd144,8'd128} : s = 9;
	{8'd144,8'd129} : s = 69;
	{8'd144,8'd130} : s = 67;
	{8'd144,8'd131} : s = 177;
	{8'd144,8'd132} : s = 56;
	{8'd144,8'd133} : s = 172;
	{8'd144,8'd134} : s = 170;
	{8'd144,8'd135} : s = 313;
	{8'd144,8'd136} : s = 52;
	{8'd144,8'd137} : s = 169;
	{8'd144,8'd138} : s = 166;
	{8'd144,8'd139} : s = 310;
	{8'd144,8'd140} : s = 165;
	{8'd144,8'd141} : s = 309;
	{8'd144,8'd142} : s = 307;
	{8'd144,8'd143} : s = 427;
	{8'd144,8'd144} : s = 6;
	{8'd144,8'd145} : s = 50;
	{8'd144,8'd146} : s = 49;
	{8'd144,8'd147} : s = 163;
	{8'd144,8'd148} : s = 44;
	{8'd144,8'd149} : s = 156;
	{8'd144,8'd150} : s = 154;
	{8'd144,8'd151} : s = 302;
	{8'd144,8'd152} : s = 42;
	{8'd144,8'd153} : s = 153;
	{8'd144,8'd154} : s = 150;
	{8'd144,8'd155} : s = 301;
	{8'd144,8'd156} : s = 149;
	{8'd144,8'd157} : s = 299;
	{8'd144,8'd158} : s = 295;
	{8'd144,8'd159} : s = 423;
	{8'd144,8'd160} : s = 41;
	{8'd144,8'd161} : s = 147;
	{8'd144,8'd162} : s = 142;
	{8'd144,8'd163} : s = 286;
	{8'd144,8'd164} : s = 141;
	{8'd144,8'd165} : s = 285;
	{8'd144,8'd166} : s = 283;
	{8'd144,8'd167} : s = 414;
	{8'd144,8'd168} : s = 139;
	{8'd144,8'd169} : s = 279;
	{8'd144,8'd170} : s = 271;
	{8'd144,8'd171} : s = 413;
	{8'd144,8'd172} : s = 248;
	{8'd144,8'd173} : s = 411;
	{8'd144,8'd174} : s = 407;
	{8'd144,8'd175} : s = 491;
	{8'd144,8'd176} : s = 5;
	{8'd144,8'd177} : s = 38;
	{8'd144,8'd178} : s = 37;
	{8'd144,8'd179} : s = 135;
	{8'd144,8'd180} : s = 35;
	{8'd144,8'd181} : s = 120;
	{8'd144,8'd182} : s = 116;
	{8'd144,8'd183} : s = 244;
	{8'd144,8'd184} : s = 28;
	{8'd144,8'd185} : s = 114;
	{8'd144,8'd186} : s = 113;
	{8'd144,8'd187} : s = 242;
	{8'd144,8'd188} : s = 108;
	{8'd144,8'd189} : s = 241;
	{8'd144,8'd190} : s = 236;
	{8'd144,8'd191} : s = 399;
	{8'd144,8'd192} : s = 26;
	{8'd144,8'd193} : s = 106;
	{8'd144,8'd194} : s = 105;
	{8'd144,8'd195} : s = 234;
	{8'd144,8'd196} : s = 102;
	{8'd144,8'd197} : s = 233;
	{8'd144,8'd198} : s = 230;
	{8'd144,8'd199} : s = 380;
	{8'd144,8'd200} : s = 101;
	{8'd144,8'd201} : s = 229;
	{8'd144,8'd202} : s = 227;
	{8'd144,8'd203} : s = 378;
	{8'd144,8'd204} : s = 220;
	{8'd144,8'd205} : s = 377;
	{8'd144,8'd206} : s = 374;
	{8'd144,8'd207} : s = 487;
	{8'd144,8'd208} : s = 25;
	{8'd144,8'd209} : s = 99;
	{8'd144,8'd210} : s = 92;
	{8'd144,8'd211} : s = 218;
	{8'd144,8'd212} : s = 90;
	{8'd144,8'd213} : s = 217;
	{8'd144,8'd214} : s = 214;
	{8'd144,8'd215} : s = 373;
	{8'd144,8'd216} : s = 89;
	{8'd144,8'd217} : s = 213;
	{8'd144,8'd218} : s = 211;
	{8'd144,8'd219} : s = 371;
	{8'd144,8'd220} : s = 206;
	{8'd144,8'd221} : s = 366;
	{8'd144,8'd222} : s = 365;
	{8'd144,8'd223} : s = 478;
	{8'd144,8'd224} : s = 86;
	{8'd144,8'd225} : s = 205;
	{8'd144,8'd226} : s = 203;
	{8'd144,8'd227} : s = 363;
	{8'd144,8'd228} : s = 199;
	{8'd144,8'd229} : s = 359;
	{8'd144,8'd230} : s = 350;
	{8'd144,8'd231} : s = 477;
	{8'd144,8'd232} : s = 188;
	{8'd144,8'd233} : s = 349;
	{8'd144,8'd234} : s = 347;
	{8'd144,8'd235} : s = 475;
	{8'd144,8'd236} : s = 343;
	{8'd144,8'd237} : s = 471;
	{8'd144,8'd238} : s = 463;
	{8'd144,8'd239} : s = 509;
	{8'd144,8'd240} : s = 3;
	{8'd144,8'd241} : s = 22;
	{8'd144,8'd242} : s = 21;
	{8'd144,8'd243} : s = 85;
	{8'd144,8'd244} : s = 19;
	{8'd144,8'd245} : s = 83;
	{8'd144,8'd246} : s = 78;
	{8'd144,8'd247} : s = 186;
	{8'd144,8'd248} : s = 14;
	{8'd144,8'd249} : s = 77;
	{8'd144,8'd250} : s = 75;
	{8'd144,8'd251} : s = 185;
	{8'd144,8'd252} : s = 71;
	{8'd144,8'd253} : s = 182;
	{8'd144,8'd254} : s = 181;
	{8'd144,8'd255} : s = 335;
	{8'd145,8'd0} : s = 146;
	{8'd145,8'd1} : s = 145;
	{8'd145,8'd2} : s = 305;
	{8'd145,8'd3} : s = 140;
	{8'd145,8'd4} : s = 300;
	{8'd145,8'd5} : s = 298;
	{8'd145,8'd6} : s = 422;
	{8'd145,8'd7} : s = 138;
	{8'd145,8'd8} : s = 297;
	{8'd145,8'd9} : s = 294;
	{8'd145,8'd10} : s = 421;
	{8'd145,8'd11} : s = 293;
	{8'd145,8'd12} : s = 419;
	{8'd145,8'd13} : s = 412;
	{8'd145,8'd14} : s = 486;
	{8'd145,8'd15} : s = 24;
	{8'd145,8'd16} : s = 137;
	{8'd145,8'd17} : s = 134;
	{8'd145,8'd18} : s = 291;
	{8'd145,8'd19} : s = 133;
	{8'd145,8'd20} : s = 284;
	{8'd145,8'd21} : s = 282;
	{8'd145,8'd22} : s = 410;
	{8'd145,8'd23} : s = 131;
	{8'd145,8'd24} : s = 281;
	{8'd145,8'd25} : s = 278;
	{8'd145,8'd26} : s = 409;
	{8'd145,8'd27} : s = 277;
	{8'd145,8'd28} : s = 406;
	{8'd145,8'd29} : s = 405;
	{8'd145,8'd30} : s = 485;
	{8'd145,8'd31} : s = 112;
	{8'd145,8'd32} : s = 275;
	{8'd145,8'd33} : s = 270;
	{8'd145,8'd34} : s = 403;
	{8'd145,8'd35} : s = 269;
	{8'd145,8'd36} : s = 398;
	{8'd145,8'd37} : s = 397;
	{8'd145,8'd38} : s = 483;
	{8'd145,8'd39} : s = 267;
	{8'd145,8'd40} : s = 395;
	{8'd145,8'd41} : s = 391;
	{8'd145,8'd42} : s = 476;
	{8'd145,8'd43} : s = 376;
	{8'd145,8'd44} : s = 474;
	{8'd145,8'd45} : s = 473;
	{8'd145,8'd46} : s = 506;
	{8'd145,8'd47} : s = 20;
	{8'd145,8'd48} : s = 104;
	{8'd145,8'd49} : s = 100;
	{8'd145,8'd50} : s = 263;
	{8'd145,8'd51} : s = 98;
	{8'd145,8'd52} : s = 240;
	{8'd145,8'd53} : s = 232;
	{8'd145,8'd54} : s = 372;
	{8'd145,8'd55} : s = 97;
	{8'd145,8'd56} : s = 228;
	{8'd145,8'd57} : s = 226;
	{8'd145,8'd58} : s = 370;
	{8'd145,8'd59} : s = 225;
	{8'd145,8'd60} : s = 369;
	{8'd145,8'd61} : s = 364;
	{8'd145,8'd62} : s = 470;
	{8'd145,8'd63} : s = 88;
	{8'd145,8'd64} : s = 216;
	{8'd145,8'd65} : s = 212;
	{8'd145,8'd66} : s = 362;
	{8'd145,8'd67} : s = 210;
	{8'd145,8'd68} : s = 361;
	{8'd145,8'd69} : s = 358;
	{8'd145,8'd70} : s = 469;
	{8'd145,8'd71} : s = 209;
	{8'd145,8'd72} : s = 357;
	{8'd145,8'd73} : s = 355;
	{8'd145,8'd74} : s = 467;
	{8'd145,8'd75} : s = 348;
	{8'd145,8'd76} : s = 462;
	{8'd145,8'd77} : s = 461;
	{8'd145,8'd78} : s = 505;
	{8'd145,8'd79} : s = 84;
	{8'd145,8'd80} : s = 204;
	{8'd145,8'd81} : s = 202;
	{8'd145,8'd82} : s = 346;
	{8'd145,8'd83} : s = 201;
	{8'd145,8'd84} : s = 345;
	{8'd145,8'd85} : s = 342;
	{8'd145,8'd86} : s = 459;
	{8'd145,8'd87} : s = 198;
	{8'd145,8'd88} : s = 341;
	{8'd145,8'd89} : s = 339;
	{8'd145,8'd90} : s = 455;
	{8'd145,8'd91} : s = 334;
	{8'd145,8'd92} : s = 444;
	{8'd145,8'd93} : s = 442;
	{8'd145,8'd94} : s = 502;
	{8'd145,8'd95} : s = 197;
	{8'd145,8'd96} : s = 333;
	{8'd145,8'd97} : s = 331;
	{8'd145,8'd98} : s = 441;
	{8'd145,8'd99} : s = 327;
	{8'd145,8'd100} : s = 438;
	{8'd145,8'd101} : s = 437;
	{8'd145,8'd102} : s = 501;
	{8'd145,8'd103} : s = 316;
	{8'd145,8'd104} : s = 435;
	{8'd145,8'd105} : s = 430;
	{8'd145,8'd106} : s = 499;
	{8'd145,8'd107} : s = 429;
	{8'd145,8'd108} : s = 494;
	{8'd145,8'd109} : s = 493;
	{8'd145,8'd110} : s = 510;
	{8'd145,8'd111} : s = 1;
	{8'd145,8'd112} : s = 18;
	{8'd145,8'd113} : s = 17;
	{8'd145,8'd114} : s = 82;
	{8'd145,8'd115} : s = 12;
	{8'd145,8'd116} : s = 81;
	{8'd145,8'd117} : s = 76;
	{8'd145,8'd118} : s = 195;
	{8'd145,8'd119} : s = 10;
	{8'd145,8'd120} : s = 74;
	{8'd145,8'd121} : s = 73;
	{8'd145,8'd122} : s = 184;
	{8'd145,8'd123} : s = 70;
	{8'd145,8'd124} : s = 180;
	{8'd145,8'd125} : s = 178;
	{8'd145,8'd126} : s = 314;
	{8'd145,8'd127} : s = 9;
	{8'd145,8'd128} : s = 69;
	{8'd145,8'd129} : s = 67;
	{8'd145,8'd130} : s = 177;
	{8'd145,8'd131} : s = 56;
	{8'd145,8'd132} : s = 172;
	{8'd145,8'd133} : s = 170;
	{8'd145,8'd134} : s = 313;
	{8'd145,8'd135} : s = 52;
	{8'd145,8'd136} : s = 169;
	{8'd145,8'd137} : s = 166;
	{8'd145,8'd138} : s = 310;
	{8'd145,8'd139} : s = 165;
	{8'd145,8'd140} : s = 309;
	{8'd145,8'd141} : s = 307;
	{8'd145,8'd142} : s = 427;
	{8'd145,8'd143} : s = 6;
	{8'd145,8'd144} : s = 50;
	{8'd145,8'd145} : s = 49;
	{8'd145,8'd146} : s = 163;
	{8'd145,8'd147} : s = 44;
	{8'd145,8'd148} : s = 156;
	{8'd145,8'd149} : s = 154;
	{8'd145,8'd150} : s = 302;
	{8'd145,8'd151} : s = 42;
	{8'd145,8'd152} : s = 153;
	{8'd145,8'd153} : s = 150;
	{8'd145,8'd154} : s = 301;
	{8'd145,8'd155} : s = 149;
	{8'd145,8'd156} : s = 299;
	{8'd145,8'd157} : s = 295;
	{8'd145,8'd158} : s = 423;
	{8'd145,8'd159} : s = 41;
	{8'd145,8'd160} : s = 147;
	{8'd145,8'd161} : s = 142;
	{8'd145,8'd162} : s = 286;
	{8'd145,8'd163} : s = 141;
	{8'd145,8'd164} : s = 285;
	{8'd145,8'd165} : s = 283;
	{8'd145,8'd166} : s = 414;
	{8'd145,8'd167} : s = 139;
	{8'd145,8'd168} : s = 279;
	{8'd145,8'd169} : s = 271;
	{8'd145,8'd170} : s = 413;
	{8'd145,8'd171} : s = 248;
	{8'd145,8'd172} : s = 411;
	{8'd145,8'd173} : s = 407;
	{8'd145,8'd174} : s = 491;
	{8'd145,8'd175} : s = 5;
	{8'd145,8'd176} : s = 38;
	{8'd145,8'd177} : s = 37;
	{8'd145,8'd178} : s = 135;
	{8'd145,8'd179} : s = 35;
	{8'd145,8'd180} : s = 120;
	{8'd145,8'd181} : s = 116;
	{8'd145,8'd182} : s = 244;
	{8'd145,8'd183} : s = 28;
	{8'd145,8'd184} : s = 114;
	{8'd145,8'd185} : s = 113;
	{8'd145,8'd186} : s = 242;
	{8'd145,8'd187} : s = 108;
	{8'd145,8'd188} : s = 241;
	{8'd145,8'd189} : s = 236;
	{8'd145,8'd190} : s = 399;
	{8'd145,8'd191} : s = 26;
	{8'd145,8'd192} : s = 106;
	{8'd145,8'd193} : s = 105;
	{8'd145,8'd194} : s = 234;
	{8'd145,8'd195} : s = 102;
	{8'd145,8'd196} : s = 233;
	{8'd145,8'd197} : s = 230;
	{8'd145,8'd198} : s = 380;
	{8'd145,8'd199} : s = 101;
	{8'd145,8'd200} : s = 229;
	{8'd145,8'd201} : s = 227;
	{8'd145,8'd202} : s = 378;
	{8'd145,8'd203} : s = 220;
	{8'd145,8'd204} : s = 377;
	{8'd145,8'd205} : s = 374;
	{8'd145,8'd206} : s = 487;
	{8'd145,8'd207} : s = 25;
	{8'd145,8'd208} : s = 99;
	{8'd145,8'd209} : s = 92;
	{8'd145,8'd210} : s = 218;
	{8'd145,8'd211} : s = 90;
	{8'd145,8'd212} : s = 217;
	{8'd145,8'd213} : s = 214;
	{8'd145,8'd214} : s = 373;
	{8'd145,8'd215} : s = 89;
	{8'd145,8'd216} : s = 213;
	{8'd145,8'd217} : s = 211;
	{8'd145,8'd218} : s = 371;
	{8'd145,8'd219} : s = 206;
	{8'd145,8'd220} : s = 366;
	{8'd145,8'd221} : s = 365;
	{8'd145,8'd222} : s = 478;
	{8'd145,8'd223} : s = 86;
	{8'd145,8'd224} : s = 205;
	{8'd145,8'd225} : s = 203;
	{8'd145,8'd226} : s = 363;
	{8'd145,8'd227} : s = 199;
	{8'd145,8'd228} : s = 359;
	{8'd145,8'd229} : s = 350;
	{8'd145,8'd230} : s = 477;
	{8'd145,8'd231} : s = 188;
	{8'd145,8'd232} : s = 349;
	{8'd145,8'd233} : s = 347;
	{8'd145,8'd234} : s = 475;
	{8'd145,8'd235} : s = 343;
	{8'd145,8'd236} : s = 471;
	{8'd145,8'd237} : s = 463;
	{8'd145,8'd238} : s = 509;
	{8'd145,8'd239} : s = 3;
	{8'd145,8'd240} : s = 22;
	{8'd145,8'd241} : s = 21;
	{8'd145,8'd242} : s = 85;
	{8'd145,8'd243} : s = 19;
	{8'd145,8'd244} : s = 83;
	{8'd145,8'd245} : s = 78;
	{8'd145,8'd246} : s = 186;
	{8'd145,8'd247} : s = 14;
	{8'd145,8'd248} : s = 77;
	{8'd145,8'd249} : s = 75;
	{8'd145,8'd250} : s = 185;
	{8'd145,8'd251} : s = 71;
	{8'd145,8'd252} : s = 182;
	{8'd145,8'd253} : s = 181;
	{8'd145,8'd254} : s = 335;
	{8'd145,8'd255} : s = 13;
	{8'd146,8'd0} : s = 145;
	{8'd146,8'd1} : s = 305;
	{8'd146,8'd2} : s = 140;
	{8'd146,8'd3} : s = 300;
	{8'd146,8'd4} : s = 298;
	{8'd146,8'd5} : s = 422;
	{8'd146,8'd6} : s = 138;
	{8'd146,8'd7} : s = 297;
	{8'd146,8'd8} : s = 294;
	{8'd146,8'd9} : s = 421;
	{8'd146,8'd10} : s = 293;
	{8'd146,8'd11} : s = 419;
	{8'd146,8'd12} : s = 412;
	{8'd146,8'd13} : s = 486;
	{8'd146,8'd14} : s = 24;
	{8'd146,8'd15} : s = 137;
	{8'd146,8'd16} : s = 134;
	{8'd146,8'd17} : s = 291;
	{8'd146,8'd18} : s = 133;
	{8'd146,8'd19} : s = 284;
	{8'd146,8'd20} : s = 282;
	{8'd146,8'd21} : s = 410;
	{8'd146,8'd22} : s = 131;
	{8'd146,8'd23} : s = 281;
	{8'd146,8'd24} : s = 278;
	{8'd146,8'd25} : s = 409;
	{8'd146,8'd26} : s = 277;
	{8'd146,8'd27} : s = 406;
	{8'd146,8'd28} : s = 405;
	{8'd146,8'd29} : s = 485;
	{8'd146,8'd30} : s = 112;
	{8'd146,8'd31} : s = 275;
	{8'd146,8'd32} : s = 270;
	{8'd146,8'd33} : s = 403;
	{8'd146,8'd34} : s = 269;
	{8'd146,8'd35} : s = 398;
	{8'd146,8'd36} : s = 397;
	{8'd146,8'd37} : s = 483;
	{8'd146,8'd38} : s = 267;
	{8'd146,8'd39} : s = 395;
	{8'd146,8'd40} : s = 391;
	{8'd146,8'd41} : s = 476;
	{8'd146,8'd42} : s = 376;
	{8'd146,8'd43} : s = 474;
	{8'd146,8'd44} : s = 473;
	{8'd146,8'd45} : s = 506;
	{8'd146,8'd46} : s = 20;
	{8'd146,8'd47} : s = 104;
	{8'd146,8'd48} : s = 100;
	{8'd146,8'd49} : s = 263;
	{8'd146,8'd50} : s = 98;
	{8'd146,8'd51} : s = 240;
	{8'd146,8'd52} : s = 232;
	{8'd146,8'd53} : s = 372;
	{8'd146,8'd54} : s = 97;
	{8'd146,8'd55} : s = 228;
	{8'd146,8'd56} : s = 226;
	{8'd146,8'd57} : s = 370;
	{8'd146,8'd58} : s = 225;
	{8'd146,8'd59} : s = 369;
	{8'd146,8'd60} : s = 364;
	{8'd146,8'd61} : s = 470;
	{8'd146,8'd62} : s = 88;
	{8'd146,8'd63} : s = 216;
	{8'd146,8'd64} : s = 212;
	{8'd146,8'd65} : s = 362;
	{8'd146,8'd66} : s = 210;
	{8'd146,8'd67} : s = 361;
	{8'd146,8'd68} : s = 358;
	{8'd146,8'd69} : s = 469;
	{8'd146,8'd70} : s = 209;
	{8'd146,8'd71} : s = 357;
	{8'd146,8'd72} : s = 355;
	{8'd146,8'd73} : s = 467;
	{8'd146,8'd74} : s = 348;
	{8'd146,8'd75} : s = 462;
	{8'd146,8'd76} : s = 461;
	{8'd146,8'd77} : s = 505;
	{8'd146,8'd78} : s = 84;
	{8'd146,8'd79} : s = 204;
	{8'd146,8'd80} : s = 202;
	{8'd146,8'd81} : s = 346;
	{8'd146,8'd82} : s = 201;
	{8'd146,8'd83} : s = 345;
	{8'd146,8'd84} : s = 342;
	{8'd146,8'd85} : s = 459;
	{8'd146,8'd86} : s = 198;
	{8'd146,8'd87} : s = 341;
	{8'd146,8'd88} : s = 339;
	{8'd146,8'd89} : s = 455;
	{8'd146,8'd90} : s = 334;
	{8'd146,8'd91} : s = 444;
	{8'd146,8'd92} : s = 442;
	{8'd146,8'd93} : s = 502;
	{8'd146,8'd94} : s = 197;
	{8'd146,8'd95} : s = 333;
	{8'd146,8'd96} : s = 331;
	{8'd146,8'd97} : s = 441;
	{8'd146,8'd98} : s = 327;
	{8'd146,8'd99} : s = 438;
	{8'd146,8'd100} : s = 437;
	{8'd146,8'd101} : s = 501;
	{8'd146,8'd102} : s = 316;
	{8'd146,8'd103} : s = 435;
	{8'd146,8'd104} : s = 430;
	{8'd146,8'd105} : s = 499;
	{8'd146,8'd106} : s = 429;
	{8'd146,8'd107} : s = 494;
	{8'd146,8'd108} : s = 493;
	{8'd146,8'd109} : s = 510;
	{8'd146,8'd110} : s = 1;
	{8'd146,8'd111} : s = 18;
	{8'd146,8'd112} : s = 17;
	{8'd146,8'd113} : s = 82;
	{8'd146,8'd114} : s = 12;
	{8'd146,8'd115} : s = 81;
	{8'd146,8'd116} : s = 76;
	{8'd146,8'd117} : s = 195;
	{8'd146,8'd118} : s = 10;
	{8'd146,8'd119} : s = 74;
	{8'd146,8'd120} : s = 73;
	{8'd146,8'd121} : s = 184;
	{8'd146,8'd122} : s = 70;
	{8'd146,8'd123} : s = 180;
	{8'd146,8'd124} : s = 178;
	{8'd146,8'd125} : s = 314;
	{8'd146,8'd126} : s = 9;
	{8'd146,8'd127} : s = 69;
	{8'd146,8'd128} : s = 67;
	{8'd146,8'd129} : s = 177;
	{8'd146,8'd130} : s = 56;
	{8'd146,8'd131} : s = 172;
	{8'd146,8'd132} : s = 170;
	{8'd146,8'd133} : s = 313;
	{8'd146,8'd134} : s = 52;
	{8'd146,8'd135} : s = 169;
	{8'd146,8'd136} : s = 166;
	{8'd146,8'd137} : s = 310;
	{8'd146,8'd138} : s = 165;
	{8'd146,8'd139} : s = 309;
	{8'd146,8'd140} : s = 307;
	{8'd146,8'd141} : s = 427;
	{8'd146,8'd142} : s = 6;
	{8'd146,8'd143} : s = 50;
	{8'd146,8'd144} : s = 49;
	{8'd146,8'd145} : s = 163;
	{8'd146,8'd146} : s = 44;
	{8'd146,8'd147} : s = 156;
	{8'd146,8'd148} : s = 154;
	{8'd146,8'd149} : s = 302;
	{8'd146,8'd150} : s = 42;
	{8'd146,8'd151} : s = 153;
	{8'd146,8'd152} : s = 150;
	{8'd146,8'd153} : s = 301;
	{8'd146,8'd154} : s = 149;
	{8'd146,8'd155} : s = 299;
	{8'd146,8'd156} : s = 295;
	{8'd146,8'd157} : s = 423;
	{8'd146,8'd158} : s = 41;
	{8'd146,8'd159} : s = 147;
	{8'd146,8'd160} : s = 142;
	{8'd146,8'd161} : s = 286;
	{8'd146,8'd162} : s = 141;
	{8'd146,8'd163} : s = 285;
	{8'd146,8'd164} : s = 283;
	{8'd146,8'd165} : s = 414;
	{8'd146,8'd166} : s = 139;
	{8'd146,8'd167} : s = 279;
	{8'd146,8'd168} : s = 271;
	{8'd146,8'd169} : s = 413;
	{8'd146,8'd170} : s = 248;
	{8'd146,8'd171} : s = 411;
	{8'd146,8'd172} : s = 407;
	{8'd146,8'd173} : s = 491;
	{8'd146,8'd174} : s = 5;
	{8'd146,8'd175} : s = 38;
	{8'd146,8'd176} : s = 37;
	{8'd146,8'd177} : s = 135;
	{8'd146,8'd178} : s = 35;
	{8'd146,8'd179} : s = 120;
	{8'd146,8'd180} : s = 116;
	{8'd146,8'd181} : s = 244;
	{8'd146,8'd182} : s = 28;
	{8'd146,8'd183} : s = 114;
	{8'd146,8'd184} : s = 113;
	{8'd146,8'd185} : s = 242;
	{8'd146,8'd186} : s = 108;
	{8'd146,8'd187} : s = 241;
	{8'd146,8'd188} : s = 236;
	{8'd146,8'd189} : s = 399;
	{8'd146,8'd190} : s = 26;
	{8'd146,8'd191} : s = 106;
	{8'd146,8'd192} : s = 105;
	{8'd146,8'd193} : s = 234;
	{8'd146,8'd194} : s = 102;
	{8'd146,8'd195} : s = 233;
	{8'd146,8'd196} : s = 230;
	{8'd146,8'd197} : s = 380;
	{8'd146,8'd198} : s = 101;
	{8'd146,8'd199} : s = 229;
	{8'd146,8'd200} : s = 227;
	{8'd146,8'd201} : s = 378;
	{8'd146,8'd202} : s = 220;
	{8'd146,8'd203} : s = 377;
	{8'd146,8'd204} : s = 374;
	{8'd146,8'd205} : s = 487;
	{8'd146,8'd206} : s = 25;
	{8'd146,8'd207} : s = 99;
	{8'd146,8'd208} : s = 92;
	{8'd146,8'd209} : s = 218;
	{8'd146,8'd210} : s = 90;
	{8'd146,8'd211} : s = 217;
	{8'd146,8'd212} : s = 214;
	{8'd146,8'd213} : s = 373;
	{8'd146,8'd214} : s = 89;
	{8'd146,8'd215} : s = 213;
	{8'd146,8'd216} : s = 211;
	{8'd146,8'd217} : s = 371;
	{8'd146,8'd218} : s = 206;
	{8'd146,8'd219} : s = 366;
	{8'd146,8'd220} : s = 365;
	{8'd146,8'd221} : s = 478;
	{8'd146,8'd222} : s = 86;
	{8'd146,8'd223} : s = 205;
	{8'd146,8'd224} : s = 203;
	{8'd146,8'd225} : s = 363;
	{8'd146,8'd226} : s = 199;
	{8'd146,8'd227} : s = 359;
	{8'd146,8'd228} : s = 350;
	{8'd146,8'd229} : s = 477;
	{8'd146,8'd230} : s = 188;
	{8'd146,8'd231} : s = 349;
	{8'd146,8'd232} : s = 347;
	{8'd146,8'd233} : s = 475;
	{8'd146,8'd234} : s = 343;
	{8'd146,8'd235} : s = 471;
	{8'd146,8'd236} : s = 463;
	{8'd146,8'd237} : s = 509;
	{8'd146,8'd238} : s = 3;
	{8'd146,8'd239} : s = 22;
	{8'd146,8'd240} : s = 21;
	{8'd146,8'd241} : s = 85;
	{8'd146,8'd242} : s = 19;
	{8'd146,8'd243} : s = 83;
	{8'd146,8'd244} : s = 78;
	{8'd146,8'd245} : s = 186;
	{8'd146,8'd246} : s = 14;
	{8'd146,8'd247} : s = 77;
	{8'd146,8'd248} : s = 75;
	{8'd146,8'd249} : s = 185;
	{8'd146,8'd250} : s = 71;
	{8'd146,8'd251} : s = 182;
	{8'd146,8'd252} : s = 181;
	{8'd146,8'd253} : s = 335;
	{8'd146,8'd254} : s = 13;
	{8'd146,8'd255} : s = 60;
	{8'd147,8'd0} : s = 305;
	{8'd147,8'd1} : s = 140;
	{8'd147,8'd2} : s = 300;
	{8'd147,8'd3} : s = 298;
	{8'd147,8'd4} : s = 422;
	{8'd147,8'd5} : s = 138;
	{8'd147,8'd6} : s = 297;
	{8'd147,8'd7} : s = 294;
	{8'd147,8'd8} : s = 421;
	{8'd147,8'd9} : s = 293;
	{8'd147,8'd10} : s = 419;
	{8'd147,8'd11} : s = 412;
	{8'd147,8'd12} : s = 486;
	{8'd147,8'd13} : s = 24;
	{8'd147,8'd14} : s = 137;
	{8'd147,8'd15} : s = 134;
	{8'd147,8'd16} : s = 291;
	{8'd147,8'd17} : s = 133;
	{8'd147,8'd18} : s = 284;
	{8'd147,8'd19} : s = 282;
	{8'd147,8'd20} : s = 410;
	{8'd147,8'd21} : s = 131;
	{8'd147,8'd22} : s = 281;
	{8'd147,8'd23} : s = 278;
	{8'd147,8'd24} : s = 409;
	{8'd147,8'd25} : s = 277;
	{8'd147,8'd26} : s = 406;
	{8'd147,8'd27} : s = 405;
	{8'd147,8'd28} : s = 485;
	{8'd147,8'd29} : s = 112;
	{8'd147,8'd30} : s = 275;
	{8'd147,8'd31} : s = 270;
	{8'd147,8'd32} : s = 403;
	{8'd147,8'd33} : s = 269;
	{8'd147,8'd34} : s = 398;
	{8'd147,8'd35} : s = 397;
	{8'd147,8'd36} : s = 483;
	{8'd147,8'd37} : s = 267;
	{8'd147,8'd38} : s = 395;
	{8'd147,8'd39} : s = 391;
	{8'd147,8'd40} : s = 476;
	{8'd147,8'd41} : s = 376;
	{8'd147,8'd42} : s = 474;
	{8'd147,8'd43} : s = 473;
	{8'd147,8'd44} : s = 506;
	{8'd147,8'd45} : s = 20;
	{8'd147,8'd46} : s = 104;
	{8'd147,8'd47} : s = 100;
	{8'd147,8'd48} : s = 263;
	{8'd147,8'd49} : s = 98;
	{8'd147,8'd50} : s = 240;
	{8'd147,8'd51} : s = 232;
	{8'd147,8'd52} : s = 372;
	{8'd147,8'd53} : s = 97;
	{8'd147,8'd54} : s = 228;
	{8'd147,8'd55} : s = 226;
	{8'd147,8'd56} : s = 370;
	{8'd147,8'd57} : s = 225;
	{8'd147,8'd58} : s = 369;
	{8'd147,8'd59} : s = 364;
	{8'd147,8'd60} : s = 470;
	{8'd147,8'd61} : s = 88;
	{8'd147,8'd62} : s = 216;
	{8'd147,8'd63} : s = 212;
	{8'd147,8'd64} : s = 362;
	{8'd147,8'd65} : s = 210;
	{8'd147,8'd66} : s = 361;
	{8'd147,8'd67} : s = 358;
	{8'd147,8'd68} : s = 469;
	{8'd147,8'd69} : s = 209;
	{8'd147,8'd70} : s = 357;
	{8'd147,8'd71} : s = 355;
	{8'd147,8'd72} : s = 467;
	{8'd147,8'd73} : s = 348;
	{8'd147,8'd74} : s = 462;
	{8'd147,8'd75} : s = 461;
	{8'd147,8'd76} : s = 505;
	{8'd147,8'd77} : s = 84;
	{8'd147,8'd78} : s = 204;
	{8'd147,8'd79} : s = 202;
	{8'd147,8'd80} : s = 346;
	{8'd147,8'd81} : s = 201;
	{8'd147,8'd82} : s = 345;
	{8'd147,8'd83} : s = 342;
	{8'd147,8'd84} : s = 459;
	{8'd147,8'd85} : s = 198;
	{8'd147,8'd86} : s = 341;
	{8'd147,8'd87} : s = 339;
	{8'd147,8'd88} : s = 455;
	{8'd147,8'd89} : s = 334;
	{8'd147,8'd90} : s = 444;
	{8'd147,8'd91} : s = 442;
	{8'd147,8'd92} : s = 502;
	{8'd147,8'd93} : s = 197;
	{8'd147,8'd94} : s = 333;
	{8'd147,8'd95} : s = 331;
	{8'd147,8'd96} : s = 441;
	{8'd147,8'd97} : s = 327;
	{8'd147,8'd98} : s = 438;
	{8'd147,8'd99} : s = 437;
	{8'd147,8'd100} : s = 501;
	{8'd147,8'd101} : s = 316;
	{8'd147,8'd102} : s = 435;
	{8'd147,8'd103} : s = 430;
	{8'd147,8'd104} : s = 499;
	{8'd147,8'd105} : s = 429;
	{8'd147,8'd106} : s = 494;
	{8'd147,8'd107} : s = 493;
	{8'd147,8'd108} : s = 510;
	{8'd147,8'd109} : s = 1;
	{8'd147,8'd110} : s = 18;
	{8'd147,8'd111} : s = 17;
	{8'd147,8'd112} : s = 82;
	{8'd147,8'd113} : s = 12;
	{8'd147,8'd114} : s = 81;
	{8'd147,8'd115} : s = 76;
	{8'd147,8'd116} : s = 195;
	{8'd147,8'd117} : s = 10;
	{8'd147,8'd118} : s = 74;
	{8'd147,8'd119} : s = 73;
	{8'd147,8'd120} : s = 184;
	{8'd147,8'd121} : s = 70;
	{8'd147,8'd122} : s = 180;
	{8'd147,8'd123} : s = 178;
	{8'd147,8'd124} : s = 314;
	{8'd147,8'd125} : s = 9;
	{8'd147,8'd126} : s = 69;
	{8'd147,8'd127} : s = 67;
	{8'd147,8'd128} : s = 177;
	{8'd147,8'd129} : s = 56;
	{8'd147,8'd130} : s = 172;
	{8'd147,8'd131} : s = 170;
	{8'd147,8'd132} : s = 313;
	{8'd147,8'd133} : s = 52;
	{8'd147,8'd134} : s = 169;
	{8'd147,8'd135} : s = 166;
	{8'd147,8'd136} : s = 310;
	{8'd147,8'd137} : s = 165;
	{8'd147,8'd138} : s = 309;
	{8'd147,8'd139} : s = 307;
	{8'd147,8'd140} : s = 427;
	{8'd147,8'd141} : s = 6;
	{8'd147,8'd142} : s = 50;
	{8'd147,8'd143} : s = 49;
	{8'd147,8'd144} : s = 163;
	{8'd147,8'd145} : s = 44;
	{8'd147,8'd146} : s = 156;
	{8'd147,8'd147} : s = 154;
	{8'd147,8'd148} : s = 302;
	{8'd147,8'd149} : s = 42;
	{8'd147,8'd150} : s = 153;
	{8'd147,8'd151} : s = 150;
	{8'd147,8'd152} : s = 301;
	{8'd147,8'd153} : s = 149;
	{8'd147,8'd154} : s = 299;
	{8'd147,8'd155} : s = 295;
	{8'd147,8'd156} : s = 423;
	{8'd147,8'd157} : s = 41;
	{8'd147,8'd158} : s = 147;
	{8'd147,8'd159} : s = 142;
	{8'd147,8'd160} : s = 286;
	{8'd147,8'd161} : s = 141;
	{8'd147,8'd162} : s = 285;
	{8'd147,8'd163} : s = 283;
	{8'd147,8'd164} : s = 414;
	{8'd147,8'd165} : s = 139;
	{8'd147,8'd166} : s = 279;
	{8'd147,8'd167} : s = 271;
	{8'd147,8'd168} : s = 413;
	{8'd147,8'd169} : s = 248;
	{8'd147,8'd170} : s = 411;
	{8'd147,8'd171} : s = 407;
	{8'd147,8'd172} : s = 491;
	{8'd147,8'd173} : s = 5;
	{8'd147,8'd174} : s = 38;
	{8'd147,8'd175} : s = 37;
	{8'd147,8'd176} : s = 135;
	{8'd147,8'd177} : s = 35;
	{8'd147,8'd178} : s = 120;
	{8'd147,8'd179} : s = 116;
	{8'd147,8'd180} : s = 244;
	{8'd147,8'd181} : s = 28;
	{8'd147,8'd182} : s = 114;
	{8'd147,8'd183} : s = 113;
	{8'd147,8'd184} : s = 242;
	{8'd147,8'd185} : s = 108;
	{8'd147,8'd186} : s = 241;
	{8'd147,8'd187} : s = 236;
	{8'd147,8'd188} : s = 399;
	{8'd147,8'd189} : s = 26;
	{8'd147,8'd190} : s = 106;
	{8'd147,8'd191} : s = 105;
	{8'd147,8'd192} : s = 234;
	{8'd147,8'd193} : s = 102;
	{8'd147,8'd194} : s = 233;
	{8'd147,8'd195} : s = 230;
	{8'd147,8'd196} : s = 380;
	{8'd147,8'd197} : s = 101;
	{8'd147,8'd198} : s = 229;
	{8'd147,8'd199} : s = 227;
	{8'd147,8'd200} : s = 378;
	{8'd147,8'd201} : s = 220;
	{8'd147,8'd202} : s = 377;
	{8'd147,8'd203} : s = 374;
	{8'd147,8'd204} : s = 487;
	{8'd147,8'd205} : s = 25;
	{8'd147,8'd206} : s = 99;
	{8'd147,8'd207} : s = 92;
	{8'd147,8'd208} : s = 218;
	{8'd147,8'd209} : s = 90;
	{8'd147,8'd210} : s = 217;
	{8'd147,8'd211} : s = 214;
	{8'd147,8'd212} : s = 373;
	{8'd147,8'd213} : s = 89;
	{8'd147,8'd214} : s = 213;
	{8'd147,8'd215} : s = 211;
	{8'd147,8'd216} : s = 371;
	{8'd147,8'd217} : s = 206;
	{8'd147,8'd218} : s = 366;
	{8'd147,8'd219} : s = 365;
	{8'd147,8'd220} : s = 478;
	{8'd147,8'd221} : s = 86;
	{8'd147,8'd222} : s = 205;
	{8'd147,8'd223} : s = 203;
	{8'd147,8'd224} : s = 363;
	{8'd147,8'd225} : s = 199;
	{8'd147,8'd226} : s = 359;
	{8'd147,8'd227} : s = 350;
	{8'd147,8'd228} : s = 477;
	{8'd147,8'd229} : s = 188;
	{8'd147,8'd230} : s = 349;
	{8'd147,8'd231} : s = 347;
	{8'd147,8'd232} : s = 475;
	{8'd147,8'd233} : s = 343;
	{8'd147,8'd234} : s = 471;
	{8'd147,8'd235} : s = 463;
	{8'd147,8'd236} : s = 509;
	{8'd147,8'd237} : s = 3;
	{8'd147,8'd238} : s = 22;
	{8'd147,8'd239} : s = 21;
	{8'd147,8'd240} : s = 85;
	{8'd147,8'd241} : s = 19;
	{8'd147,8'd242} : s = 83;
	{8'd147,8'd243} : s = 78;
	{8'd147,8'd244} : s = 186;
	{8'd147,8'd245} : s = 14;
	{8'd147,8'd246} : s = 77;
	{8'd147,8'd247} : s = 75;
	{8'd147,8'd248} : s = 185;
	{8'd147,8'd249} : s = 71;
	{8'd147,8'd250} : s = 182;
	{8'd147,8'd251} : s = 181;
	{8'd147,8'd252} : s = 335;
	{8'd147,8'd253} : s = 13;
	{8'd147,8'd254} : s = 60;
	{8'd147,8'd255} : s = 58;
	{8'd148,8'd0} : s = 140;
	{8'd148,8'd1} : s = 300;
	{8'd148,8'd2} : s = 298;
	{8'd148,8'd3} : s = 422;
	{8'd148,8'd4} : s = 138;
	{8'd148,8'd5} : s = 297;
	{8'd148,8'd6} : s = 294;
	{8'd148,8'd7} : s = 421;
	{8'd148,8'd8} : s = 293;
	{8'd148,8'd9} : s = 419;
	{8'd148,8'd10} : s = 412;
	{8'd148,8'd11} : s = 486;
	{8'd148,8'd12} : s = 24;
	{8'd148,8'd13} : s = 137;
	{8'd148,8'd14} : s = 134;
	{8'd148,8'd15} : s = 291;
	{8'd148,8'd16} : s = 133;
	{8'd148,8'd17} : s = 284;
	{8'd148,8'd18} : s = 282;
	{8'd148,8'd19} : s = 410;
	{8'd148,8'd20} : s = 131;
	{8'd148,8'd21} : s = 281;
	{8'd148,8'd22} : s = 278;
	{8'd148,8'd23} : s = 409;
	{8'd148,8'd24} : s = 277;
	{8'd148,8'd25} : s = 406;
	{8'd148,8'd26} : s = 405;
	{8'd148,8'd27} : s = 485;
	{8'd148,8'd28} : s = 112;
	{8'd148,8'd29} : s = 275;
	{8'd148,8'd30} : s = 270;
	{8'd148,8'd31} : s = 403;
	{8'd148,8'd32} : s = 269;
	{8'd148,8'd33} : s = 398;
	{8'd148,8'd34} : s = 397;
	{8'd148,8'd35} : s = 483;
	{8'd148,8'd36} : s = 267;
	{8'd148,8'd37} : s = 395;
	{8'd148,8'd38} : s = 391;
	{8'd148,8'd39} : s = 476;
	{8'd148,8'd40} : s = 376;
	{8'd148,8'd41} : s = 474;
	{8'd148,8'd42} : s = 473;
	{8'd148,8'd43} : s = 506;
	{8'd148,8'd44} : s = 20;
	{8'd148,8'd45} : s = 104;
	{8'd148,8'd46} : s = 100;
	{8'd148,8'd47} : s = 263;
	{8'd148,8'd48} : s = 98;
	{8'd148,8'd49} : s = 240;
	{8'd148,8'd50} : s = 232;
	{8'd148,8'd51} : s = 372;
	{8'd148,8'd52} : s = 97;
	{8'd148,8'd53} : s = 228;
	{8'd148,8'd54} : s = 226;
	{8'd148,8'd55} : s = 370;
	{8'd148,8'd56} : s = 225;
	{8'd148,8'd57} : s = 369;
	{8'd148,8'd58} : s = 364;
	{8'd148,8'd59} : s = 470;
	{8'd148,8'd60} : s = 88;
	{8'd148,8'd61} : s = 216;
	{8'd148,8'd62} : s = 212;
	{8'd148,8'd63} : s = 362;
	{8'd148,8'd64} : s = 210;
	{8'd148,8'd65} : s = 361;
	{8'd148,8'd66} : s = 358;
	{8'd148,8'd67} : s = 469;
	{8'd148,8'd68} : s = 209;
	{8'd148,8'd69} : s = 357;
	{8'd148,8'd70} : s = 355;
	{8'd148,8'd71} : s = 467;
	{8'd148,8'd72} : s = 348;
	{8'd148,8'd73} : s = 462;
	{8'd148,8'd74} : s = 461;
	{8'd148,8'd75} : s = 505;
	{8'd148,8'd76} : s = 84;
	{8'd148,8'd77} : s = 204;
	{8'd148,8'd78} : s = 202;
	{8'd148,8'd79} : s = 346;
	{8'd148,8'd80} : s = 201;
	{8'd148,8'd81} : s = 345;
	{8'd148,8'd82} : s = 342;
	{8'd148,8'd83} : s = 459;
	{8'd148,8'd84} : s = 198;
	{8'd148,8'd85} : s = 341;
	{8'd148,8'd86} : s = 339;
	{8'd148,8'd87} : s = 455;
	{8'd148,8'd88} : s = 334;
	{8'd148,8'd89} : s = 444;
	{8'd148,8'd90} : s = 442;
	{8'd148,8'd91} : s = 502;
	{8'd148,8'd92} : s = 197;
	{8'd148,8'd93} : s = 333;
	{8'd148,8'd94} : s = 331;
	{8'd148,8'd95} : s = 441;
	{8'd148,8'd96} : s = 327;
	{8'd148,8'd97} : s = 438;
	{8'd148,8'd98} : s = 437;
	{8'd148,8'd99} : s = 501;
	{8'd148,8'd100} : s = 316;
	{8'd148,8'd101} : s = 435;
	{8'd148,8'd102} : s = 430;
	{8'd148,8'd103} : s = 499;
	{8'd148,8'd104} : s = 429;
	{8'd148,8'd105} : s = 494;
	{8'd148,8'd106} : s = 493;
	{8'd148,8'd107} : s = 510;
	{8'd148,8'd108} : s = 1;
	{8'd148,8'd109} : s = 18;
	{8'd148,8'd110} : s = 17;
	{8'd148,8'd111} : s = 82;
	{8'd148,8'd112} : s = 12;
	{8'd148,8'd113} : s = 81;
	{8'd148,8'd114} : s = 76;
	{8'd148,8'd115} : s = 195;
	{8'd148,8'd116} : s = 10;
	{8'd148,8'd117} : s = 74;
	{8'd148,8'd118} : s = 73;
	{8'd148,8'd119} : s = 184;
	{8'd148,8'd120} : s = 70;
	{8'd148,8'd121} : s = 180;
	{8'd148,8'd122} : s = 178;
	{8'd148,8'd123} : s = 314;
	{8'd148,8'd124} : s = 9;
	{8'd148,8'd125} : s = 69;
	{8'd148,8'd126} : s = 67;
	{8'd148,8'd127} : s = 177;
	{8'd148,8'd128} : s = 56;
	{8'd148,8'd129} : s = 172;
	{8'd148,8'd130} : s = 170;
	{8'd148,8'd131} : s = 313;
	{8'd148,8'd132} : s = 52;
	{8'd148,8'd133} : s = 169;
	{8'd148,8'd134} : s = 166;
	{8'd148,8'd135} : s = 310;
	{8'd148,8'd136} : s = 165;
	{8'd148,8'd137} : s = 309;
	{8'd148,8'd138} : s = 307;
	{8'd148,8'd139} : s = 427;
	{8'd148,8'd140} : s = 6;
	{8'd148,8'd141} : s = 50;
	{8'd148,8'd142} : s = 49;
	{8'd148,8'd143} : s = 163;
	{8'd148,8'd144} : s = 44;
	{8'd148,8'd145} : s = 156;
	{8'd148,8'd146} : s = 154;
	{8'd148,8'd147} : s = 302;
	{8'd148,8'd148} : s = 42;
	{8'd148,8'd149} : s = 153;
	{8'd148,8'd150} : s = 150;
	{8'd148,8'd151} : s = 301;
	{8'd148,8'd152} : s = 149;
	{8'd148,8'd153} : s = 299;
	{8'd148,8'd154} : s = 295;
	{8'd148,8'd155} : s = 423;
	{8'd148,8'd156} : s = 41;
	{8'd148,8'd157} : s = 147;
	{8'd148,8'd158} : s = 142;
	{8'd148,8'd159} : s = 286;
	{8'd148,8'd160} : s = 141;
	{8'd148,8'd161} : s = 285;
	{8'd148,8'd162} : s = 283;
	{8'd148,8'd163} : s = 414;
	{8'd148,8'd164} : s = 139;
	{8'd148,8'd165} : s = 279;
	{8'd148,8'd166} : s = 271;
	{8'd148,8'd167} : s = 413;
	{8'd148,8'd168} : s = 248;
	{8'd148,8'd169} : s = 411;
	{8'd148,8'd170} : s = 407;
	{8'd148,8'd171} : s = 491;
	{8'd148,8'd172} : s = 5;
	{8'd148,8'd173} : s = 38;
	{8'd148,8'd174} : s = 37;
	{8'd148,8'd175} : s = 135;
	{8'd148,8'd176} : s = 35;
	{8'd148,8'd177} : s = 120;
	{8'd148,8'd178} : s = 116;
	{8'd148,8'd179} : s = 244;
	{8'd148,8'd180} : s = 28;
	{8'd148,8'd181} : s = 114;
	{8'd148,8'd182} : s = 113;
	{8'd148,8'd183} : s = 242;
	{8'd148,8'd184} : s = 108;
	{8'd148,8'd185} : s = 241;
	{8'd148,8'd186} : s = 236;
	{8'd148,8'd187} : s = 399;
	{8'd148,8'd188} : s = 26;
	{8'd148,8'd189} : s = 106;
	{8'd148,8'd190} : s = 105;
	{8'd148,8'd191} : s = 234;
	{8'd148,8'd192} : s = 102;
	{8'd148,8'd193} : s = 233;
	{8'd148,8'd194} : s = 230;
	{8'd148,8'd195} : s = 380;
	{8'd148,8'd196} : s = 101;
	{8'd148,8'd197} : s = 229;
	{8'd148,8'd198} : s = 227;
	{8'd148,8'd199} : s = 378;
	{8'd148,8'd200} : s = 220;
	{8'd148,8'd201} : s = 377;
	{8'd148,8'd202} : s = 374;
	{8'd148,8'd203} : s = 487;
	{8'd148,8'd204} : s = 25;
	{8'd148,8'd205} : s = 99;
	{8'd148,8'd206} : s = 92;
	{8'd148,8'd207} : s = 218;
	{8'd148,8'd208} : s = 90;
	{8'd148,8'd209} : s = 217;
	{8'd148,8'd210} : s = 214;
	{8'd148,8'd211} : s = 373;
	{8'd148,8'd212} : s = 89;
	{8'd148,8'd213} : s = 213;
	{8'd148,8'd214} : s = 211;
	{8'd148,8'd215} : s = 371;
	{8'd148,8'd216} : s = 206;
	{8'd148,8'd217} : s = 366;
	{8'd148,8'd218} : s = 365;
	{8'd148,8'd219} : s = 478;
	{8'd148,8'd220} : s = 86;
	{8'd148,8'd221} : s = 205;
	{8'd148,8'd222} : s = 203;
	{8'd148,8'd223} : s = 363;
	{8'd148,8'd224} : s = 199;
	{8'd148,8'd225} : s = 359;
	{8'd148,8'd226} : s = 350;
	{8'd148,8'd227} : s = 477;
	{8'd148,8'd228} : s = 188;
	{8'd148,8'd229} : s = 349;
	{8'd148,8'd230} : s = 347;
	{8'd148,8'd231} : s = 475;
	{8'd148,8'd232} : s = 343;
	{8'd148,8'd233} : s = 471;
	{8'd148,8'd234} : s = 463;
	{8'd148,8'd235} : s = 509;
	{8'd148,8'd236} : s = 3;
	{8'd148,8'd237} : s = 22;
	{8'd148,8'd238} : s = 21;
	{8'd148,8'd239} : s = 85;
	{8'd148,8'd240} : s = 19;
	{8'd148,8'd241} : s = 83;
	{8'd148,8'd242} : s = 78;
	{8'd148,8'd243} : s = 186;
	{8'd148,8'd244} : s = 14;
	{8'd148,8'd245} : s = 77;
	{8'd148,8'd246} : s = 75;
	{8'd148,8'd247} : s = 185;
	{8'd148,8'd248} : s = 71;
	{8'd148,8'd249} : s = 182;
	{8'd148,8'd250} : s = 181;
	{8'd148,8'd251} : s = 335;
	{8'd148,8'd252} : s = 13;
	{8'd148,8'd253} : s = 60;
	{8'd148,8'd254} : s = 58;
	{8'd148,8'd255} : s = 179;
	{8'd149,8'd0} : s = 300;
	{8'd149,8'd1} : s = 298;
	{8'd149,8'd2} : s = 422;
	{8'd149,8'd3} : s = 138;
	{8'd149,8'd4} : s = 297;
	{8'd149,8'd5} : s = 294;
	{8'd149,8'd6} : s = 421;
	{8'd149,8'd7} : s = 293;
	{8'd149,8'd8} : s = 419;
	{8'd149,8'd9} : s = 412;
	{8'd149,8'd10} : s = 486;
	{8'd149,8'd11} : s = 24;
	{8'd149,8'd12} : s = 137;
	{8'd149,8'd13} : s = 134;
	{8'd149,8'd14} : s = 291;
	{8'd149,8'd15} : s = 133;
	{8'd149,8'd16} : s = 284;
	{8'd149,8'd17} : s = 282;
	{8'd149,8'd18} : s = 410;
	{8'd149,8'd19} : s = 131;
	{8'd149,8'd20} : s = 281;
	{8'd149,8'd21} : s = 278;
	{8'd149,8'd22} : s = 409;
	{8'd149,8'd23} : s = 277;
	{8'd149,8'd24} : s = 406;
	{8'd149,8'd25} : s = 405;
	{8'd149,8'd26} : s = 485;
	{8'd149,8'd27} : s = 112;
	{8'd149,8'd28} : s = 275;
	{8'd149,8'd29} : s = 270;
	{8'd149,8'd30} : s = 403;
	{8'd149,8'd31} : s = 269;
	{8'd149,8'd32} : s = 398;
	{8'd149,8'd33} : s = 397;
	{8'd149,8'd34} : s = 483;
	{8'd149,8'd35} : s = 267;
	{8'd149,8'd36} : s = 395;
	{8'd149,8'd37} : s = 391;
	{8'd149,8'd38} : s = 476;
	{8'd149,8'd39} : s = 376;
	{8'd149,8'd40} : s = 474;
	{8'd149,8'd41} : s = 473;
	{8'd149,8'd42} : s = 506;
	{8'd149,8'd43} : s = 20;
	{8'd149,8'd44} : s = 104;
	{8'd149,8'd45} : s = 100;
	{8'd149,8'd46} : s = 263;
	{8'd149,8'd47} : s = 98;
	{8'd149,8'd48} : s = 240;
	{8'd149,8'd49} : s = 232;
	{8'd149,8'd50} : s = 372;
	{8'd149,8'd51} : s = 97;
	{8'd149,8'd52} : s = 228;
	{8'd149,8'd53} : s = 226;
	{8'd149,8'd54} : s = 370;
	{8'd149,8'd55} : s = 225;
	{8'd149,8'd56} : s = 369;
	{8'd149,8'd57} : s = 364;
	{8'd149,8'd58} : s = 470;
	{8'd149,8'd59} : s = 88;
	{8'd149,8'd60} : s = 216;
	{8'd149,8'd61} : s = 212;
	{8'd149,8'd62} : s = 362;
	{8'd149,8'd63} : s = 210;
	{8'd149,8'd64} : s = 361;
	{8'd149,8'd65} : s = 358;
	{8'd149,8'd66} : s = 469;
	{8'd149,8'd67} : s = 209;
	{8'd149,8'd68} : s = 357;
	{8'd149,8'd69} : s = 355;
	{8'd149,8'd70} : s = 467;
	{8'd149,8'd71} : s = 348;
	{8'd149,8'd72} : s = 462;
	{8'd149,8'd73} : s = 461;
	{8'd149,8'd74} : s = 505;
	{8'd149,8'd75} : s = 84;
	{8'd149,8'd76} : s = 204;
	{8'd149,8'd77} : s = 202;
	{8'd149,8'd78} : s = 346;
	{8'd149,8'd79} : s = 201;
	{8'd149,8'd80} : s = 345;
	{8'd149,8'd81} : s = 342;
	{8'd149,8'd82} : s = 459;
	{8'd149,8'd83} : s = 198;
	{8'd149,8'd84} : s = 341;
	{8'd149,8'd85} : s = 339;
	{8'd149,8'd86} : s = 455;
	{8'd149,8'd87} : s = 334;
	{8'd149,8'd88} : s = 444;
	{8'd149,8'd89} : s = 442;
	{8'd149,8'd90} : s = 502;
	{8'd149,8'd91} : s = 197;
	{8'd149,8'd92} : s = 333;
	{8'd149,8'd93} : s = 331;
	{8'd149,8'd94} : s = 441;
	{8'd149,8'd95} : s = 327;
	{8'd149,8'd96} : s = 438;
	{8'd149,8'd97} : s = 437;
	{8'd149,8'd98} : s = 501;
	{8'd149,8'd99} : s = 316;
	{8'd149,8'd100} : s = 435;
	{8'd149,8'd101} : s = 430;
	{8'd149,8'd102} : s = 499;
	{8'd149,8'd103} : s = 429;
	{8'd149,8'd104} : s = 494;
	{8'd149,8'd105} : s = 493;
	{8'd149,8'd106} : s = 510;
	{8'd149,8'd107} : s = 1;
	{8'd149,8'd108} : s = 18;
	{8'd149,8'd109} : s = 17;
	{8'd149,8'd110} : s = 82;
	{8'd149,8'd111} : s = 12;
	{8'd149,8'd112} : s = 81;
	{8'd149,8'd113} : s = 76;
	{8'd149,8'd114} : s = 195;
	{8'd149,8'd115} : s = 10;
	{8'd149,8'd116} : s = 74;
	{8'd149,8'd117} : s = 73;
	{8'd149,8'd118} : s = 184;
	{8'd149,8'd119} : s = 70;
	{8'd149,8'd120} : s = 180;
	{8'd149,8'd121} : s = 178;
	{8'd149,8'd122} : s = 314;
	{8'd149,8'd123} : s = 9;
	{8'd149,8'd124} : s = 69;
	{8'd149,8'd125} : s = 67;
	{8'd149,8'd126} : s = 177;
	{8'd149,8'd127} : s = 56;
	{8'd149,8'd128} : s = 172;
	{8'd149,8'd129} : s = 170;
	{8'd149,8'd130} : s = 313;
	{8'd149,8'd131} : s = 52;
	{8'd149,8'd132} : s = 169;
	{8'd149,8'd133} : s = 166;
	{8'd149,8'd134} : s = 310;
	{8'd149,8'd135} : s = 165;
	{8'd149,8'd136} : s = 309;
	{8'd149,8'd137} : s = 307;
	{8'd149,8'd138} : s = 427;
	{8'd149,8'd139} : s = 6;
	{8'd149,8'd140} : s = 50;
	{8'd149,8'd141} : s = 49;
	{8'd149,8'd142} : s = 163;
	{8'd149,8'd143} : s = 44;
	{8'd149,8'd144} : s = 156;
	{8'd149,8'd145} : s = 154;
	{8'd149,8'd146} : s = 302;
	{8'd149,8'd147} : s = 42;
	{8'd149,8'd148} : s = 153;
	{8'd149,8'd149} : s = 150;
	{8'd149,8'd150} : s = 301;
	{8'd149,8'd151} : s = 149;
	{8'd149,8'd152} : s = 299;
	{8'd149,8'd153} : s = 295;
	{8'd149,8'd154} : s = 423;
	{8'd149,8'd155} : s = 41;
	{8'd149,8'd156} : s = 147;
	{8'd149,8'd157} : s = 142;
	{8'd149,8'd158} : s = 286;
	{8'd149,8'd159} : s = 141;
	{8'd149,8'd160} : s = 285;
	{8'd149,8'd161} : s = 283;
	{8'd149,8'd162} : s = 414;
	{8'd149,8'd163} : s = 139;
	{8'd149,8'd164} : s = 279;
	{8'd149,8'd165} : s = 271;
	{8'd149,8'd166} : s = 413;
	{8'd149,8'd167} : s = 248;
	{8'd149,8'd168} : s = 411;
	{8'd149,8'd169} : s = 407;
	{8'd149,8'd170} : s = 491;
	{8'd149,8'd171} : s = 5;
	{8'd149,8'd172} : s = 38;
	{8'd149,8'd173} : s = 37;
	{8'd149,8'd174} : s = 135;
	{8'd149,8'd175} : s = 35;
	{8'd149,8'd176} : s = 120;
	{8'd149,8'd177} : s = 116;
	{8'd149,8'd178} : s = 244;
	{8'd149,8'd179} : s = 28;
	{8'd149,8'd180} : s = 114;
	{8'd149,8'd181} : s = 113;
	{8'd149,8'd182} : s = 242;
	{8'd149,8'd183} : s = 108;
	{8'd149,8'd184} : s = 241;
	{8'd149,8'd185} : s = 236;
	{8'd149,8'd186} : s = 399;
	{8'd149,8'd187} : s = 26;
	{8'd149,8'd188} : s = 106;
	{8'd149,8'd189} : s = 105;
	{8'd149,8'd190} : s = 234;
	{8'd149,8'd191} : s = 102;
	{8'd149,8'd192} : s = 233;
	{8'd149,8'd193} : s = 230;
	{8'd149,8'd194} : s = 380;
	{8'd149,8'd195} : s = 101;
	{8'd149,8'd196} : s = 229;
	{8'd149,8'd197} : s = 227;
	{8'd149,8'd198} : s = 378;
	{8'd149,8'd199} : s = 220;
	{8'd149,8'd200} : s = 377;
	{8'd149,8'd201} : s = 374;
	{8'd149,8'd202} : s = 487;
	{8'd149,8'd203} : s = 25;
	{8'd149,8'd204} : s = 99;
	{8'd149,8'd205} : s = 92;
	{8'd149,8'd206} : s = 218;
	{8'd149,8'd207} : s = 90;
	{8'd149,8'd208} : s = 217;
	{8'd149,8'd209} : s = 214;
	{8'd149,8'd210} : s = 373;
	{8'd149,8'd211} : s = 89;
	{8'd149,8'd212} : s = 213;
	{8'd149,8'd213} : s = 211;
	{8'd149,8'd214} : s = 371;
	{8'd149,8'd215} : s = 206;
	{8'd149,8'd216} : s = 366;
	{8'd149,8'd217} : s = 365;
	{8'd149,8'd218} : s = 478;
	{8'd149,8'd219} : s = 86;
	{8'd149,8'd220} : s = 205;
	{8'd149,8'd221} : s = 203;
	{8'd149,8'd222} : s = 363;
	{8'd149,8'd223} : s = 199;
	{8'd149,8'd224} : s = 359;
	{8'd149,8'd225} : s = 350;
	{8'd149,8'd226} : s = 477;
	{8'd149,8'd227} : s = 188;
	{8'd149,8'd228} : s = 349;
	{8'd149,8'd229} : s = 347;
	{8'd149,8'd230} : s = 475;
	{8'd149,8'd231} : s = 343;
	{8'd149,8'd232} : s = 471;
	{8'd149,8'd233} : s = 463;
	{8'd149,8'd234} : s = 509;
	{8'd149,8'd235} : s = 3;
	{8'd149,8'd236} : s = 22;
	{8'd149,8'd237} : s = 21;
	{8'd149,8'd238} : s = 85;
	{8'd149,8'd239} : s = 19;
	{8'd149,8'd240} : s = 83;
	{8'd149,8'd241} : s = 78;
	{8'd149,8'd242} : s = 186;
	{8'd149,8'd243} : s = 14;
	{8'd149,8'd244} : s = 77;
	{8'd149,8'd245} : s = 75;
	{8'd149,8'd246} : s = 185;
	{8'd149,8'd247} : s = 71;
	{8'd149,8'd248} : s = 182;
	{8'd149,8'd249} : s = 181;
	{8'd149,8'd250} : s = 335;
	{8'd149,8'd251} : s = 13;
	{8'd149,8'd252} : s = 60;
	{8'd149,8'd253} : s = 58;
	{8'd149,8'd254} : s = 179;
	{8'd149,8'd255} : s = 57;
	{8'd150,8'd0} : s = 298;
	{8'd150,8'd1} : s = 422;
	{8'd150,8'd2} : s = 138;
	{8'd150,8'd3} : s = 297;
	{8'd150,8'd4} : s = 294;
	{8'd150,8'd5} : s = 421;
	{8'd150,8'd6} : s = 293;
	{8'd150,8'd7} : s = 419;
	{8'd150,8'd8} : s = 412;
	{8'd150,8'd9} : s = 486;
	{8'd150,8'd10} : s = 24;
	{8'd150,8'd11} : s = 137;
	{8'd150,8'd12} : s = 134;
	{8'd150,8'd13} : s = 291;
	{8'd150,8'd14} : s = 133;
	{8'd150,8'd15} : s = 284;
	{8'd150,8'd16} : s = 282;
	{8'd150,8'd17} : s = 410;
	{8'd150,8'd18} : s = 131;
	{8'd150,8'd19} : s = 281;
	{8'd150,8'd20} : s = 278;
	{8'd150,8'd21} : s = 409;
	{8'd150,8'd22} : s = 277;
	{8'd150,8'd23} : s = 406;
	{8'd150,8'd24} : s = 405;
	{8'd150,8'd25} : s = 485;
	{8'd150,8'd26} : s = 112;
	{8'd150,8'd27} : s = 275;
	{8'd150,8'd28} : s = 270;
	{8'd150,8'd29} : s = 403;
	{8'd150,8'd30} : s = 269;
	{8'd150,8'd31} : s = 398;
	{8'd150,8'd32} : s = 397;
	{8'd150,8'd33} : s = 483;
	{8'd150,8'd34} : s = 267;
	{8'd150,8'd35} : s = 395;
	{8'd150,8'd36} : s = 391;
	{8'd150,8'd37} : s = 476;
	{8'd150,8'd38} : s = 376;
	{8'd150,8'd39} : s = 474;
	{8'd150,8'd40} : s = 473;
	{8'd150,8'd41} : s = 506;
	{8'd150,8'd42} : s = 20;
	{8'd150,8'd43} : s = 104;
	{8'd150,8'd44} : s = 100;
	{8'd150,8'd45} : s = 263;
	{8'd150,8'd46} : s = 98;
	{8'd150,8'd47} : s = 240;
	{8'd150,8'd48} : s = 232;
	{8'd150,8'd49} : s = 372;
	{8'd150,8'd50} : s = 97;
	{8'd150,8'd51} : s = 228;
	{8'd150,8'd52} : s = 226;
	{8'd150,8'd53} : s = 370;
	{8'd150,8'd54} : s = 225;
	{8'd150,8'd55} : s = 369;
	{8'd150,8'd56} : s = 364;
	{8'd150,8'd57} : s = 470;
	{8'd150,8'd58} : s = 88;
	{8'd150,8'd59} : s = 216;
	{8'd150,8'd60} : s = 212;
	{8'd150,8'd61} : s = 362;
	{8'd150,8'd62} : s = 210;
	{8'd150,8'd63} : s = 361;
	{8'd150,8'd64} : s = 358;
	{8'd150,8'd65} : s = 469;
	{8'd150,8'd66} : s = 209;
	{8'd150,8'd67} : s = 357;
	{8'd150,8'd68} : s = 355;
	{8'd150,8'd69} : s = 467;
	{8'd150,8'd70} : s = 348;
	{8'd150,8'd71} : s = 462;
	{8'd150,8'd72} : s = 461;
	{8'd150,8'd73} : s = 505;
	{8'd150,8'd74} : s = 84;
	{8'd150,8'd75} : s = 204;
	{8'd150,8'd76} : s = 202;
	{8'd150,8'd77} : s = 346;
	{8'd150,8'd78} : s = 201;
	{8'd150,8'd79} : s = 345;
	{8'd150,8'd80} : s = 342;
	{8'd150,8'd81} : s = 459;
	{8'd150,8'd82} : s = 198;
	{8'd150,8'd83} : s = 341;
	{8'd150,8'd84} : s = 339;
	{8'd150,8'd85} : s = 455;
	{8'd150,8'd86} : s = 334;
	{8'd150,8'd87} : s = 444;
	{8'd150,8'd88} : s = 442;
	{8'd150,8'd89} : s = 502;
	{8'd150,8'd90} : s = 197;
	{8'd150,8'd91} : s = 333;
	{8'd150,8'd92} : s = 331;
	{8'd150,8'd93} : s = 441;
	{8'd150,8'd94} : s = 327;
	{8'd150,8'd95} : s = 438;
	{8'd150,8'd96} : s = 437;
	{8'd150,8'd97} : s = 501;
	{8'd150,8'd98} : s = 316;
	{8'd150,8'd99} : s = 435;
	{8'd150,8'd100} : s = 430;
	{8'd150,8'd101} : s = 499;
	{8'd150,8'd102} : s = 429;
	{8'd150,8'd103} : s = 494;
	{8'd150,8'd104} : s = 493;
	{8'd150,8'd105} : s = 510;
	{8'd150,8'd106} : s = 1;
	{8'd150,8'd107} : s = 18;
	{8'd150,8'd108} : s = 17;
	{8'd150,8'd109} : s = 82;
	{8'd150,8'd110} : s = 12;
	{8'd150,8'd111} : s = 81;
	{8'd150,8'd112} : s = 76;
	{8'd150,8'd113} : s = 195;
	{8'd150,8'd114} : s = 10;
	{8'd150,8'd115} : s = 74;
	{8'd150,8'd116} : s = 73;
	{8'd150,8'd117} : s = 184;
	{8'd150,8'd118} : s = 70;
	{8'd150,8'd119} : s = 180;
	{8'd150,8'd120} : s = 178;
	{8'd150,8'd121} : s = 314;
	{8'd150,8'd122} : s = 9;
	{8'd150,8'd123} : s = 69;
	{8'd150,8'd124} : s = 67;
	{8'd150,8'd125} : s = 177;
	{8'd150,8'd126} : s = 56;
	{8'd150,8'd127} : s = 172;
	{8'd150,8'd128} : s = 170;
	{8'd150,8'd129} : s = 313;
	{8'd150,8'd130} : s = 52;
	{8'd150,8'd131} : s = 169;
	{8'd150,8'd132} : s = 166;
	{8'd150,8'd133} : s = 310;
	{8'd150,8'd134} : s = 165;
	{8'd150,8'd135} : s = 309;
	{8'd150,8'd136} : s = 307;
	{8'd150,8'd137} : s = 427;
	{8'd150,8'd138} : s = 6;
	{8'd150,8'd139} : s = 50;
	{8'd150,8'd140} : s = 49;
	{8'd150,8'd141} : s = 163;
	{8'd150,8'd142} : s = 44;
	{8'd150,8'd143} : s = 156;
	{8'd150,8'd144} : s = 154;
	{8'd150,8'd145} : s = 302;
	{8'd150,8'd146} : s = 42;
	{8'd150,8'd147} : s = 153;
	{8'd150,8'd148} : s = 150;
	{8'd150,8'd149} : s = 301;
	{8'd150,8'd150} : s = 149;
	{8'd150,8'd151} : s = 299;
	{8'd150,8'd152} : s = 295;
	{8'd150,8'd153} : s = 423;
	{8'd150,8'd154} : s = 41;
	{8'd150,8'd155} : s = 147;
	{8'd150,8'd156} : s = 142;
	{8'd150,8'd157} : s = 286;
	{8'd150,8'd158} : s = 141;
	{8'd150,8'd159} : s = 285;
	{8'd150,8'd160} : s = 283;
	{8'd150,8'd161} : s = 414;
	{8'd150,8'd162} : s = 139;
	{8'd150,8'd163} : s = 279;
	{8'd150,8'd164} : s = 271;
	{8'd150,8'd165} : s = 413;
	{8'd150,8'd166} : s = 248;
	{8'd150,8'd167} : s = 411;
	{8'd150,8'd168} : s = 407;
	{8'd150,8'd169} : s = 491;
	{8'd150,8'd170} : s = 5;
	{8'd150,8'd171} : s = 38;
	{8'd150,8'd172} : s = 37;
	{8'd150,8'd173} : s = 135;
	{8'd150,8'd174} : s = 35;
	{8'd150,8'd175} : s = 120;
	{8'd150,8'd176} : s = 116;
	{8'd150,8'd177} : s = 244;
	{8'd150,8'd178} : s = 28;
	{8'd150,8'd179} : s = 114;
	{8'd150,8'd180} : s = 113;
	{8'd150,8'd181} : s = 242;
	{8'd150,8'd182} : s = 108;
	{8'd150,8'd183} : s = 241;
	{8'd150,8'd184} : s = 236;
	{8'd150,8'd185} : s = 399;
	{8'd150,8'd186} : s = 26;
	{8'd150,8'd187} : s = 106;
	{8'd150,8'd188} : s = 105;
	{8'd150,8'd189} : s = 234;
	{8'd150,8'd190} : s = 102;
	{8'd150,8'd191} : s = 233;
	{8'd150,8'd192} : s = 230;
	{8'd150,8'd193} : s = 380;
	{8'd150,8'd194} : s = 101;
	{8'd150,8'd195} : s = 229;
	{8'd150,8'd196} : s = 227;
	{8'd150,8'd197} : s = 378;
	{8'd150,8'd198} : s = 220;
	{8'd150,8'd199} : s = 377;
	{8'd150,8'd200} : s = 374;
	{8'd150,8'd201} : s = 487;
	{8'd150,8'd202} : s = 25;
	{8'd150,8'd203} : s = 99;
	{8'd150,8'd204} : s = 92;
	{8'd150,8'd205} : s = 218;
	{8'd150,8'd206} : s = 90;
	{8'd150,8'd207} : s = 217;
	{8'd150,8'd208} : s = 214;
	{8'd150,8'd209} : s = 373;
	{8'd150,8'd210} : s = 89;
	{8'd150,8'd211} : s = 213;
	{8'd150,8'd212} : s = 211;
	{8'd150,8'd213} : s = 371;
	{8'd150,8'd214} : s = 206;
	{8'd150,8'd215} : s = 366;
	{8'd150,8'd216} : s = 365;
	{8'd150,8'd217} : s = 478;
	{8'd150,8'd218} : s = 86;
	{8'd150,8'd219} : s = 205;
	{8'd150,8'd220} : s = 203;
	{8'd150,8'd221} : s = 363;
	{8'd150,8'd222} : s = 199;
	{8'd150,8'd223} : s = 359;
	{8'd150,8'd224} : s = 350;
	{8'd150,8'd225} : s = 477;
	{8'd150,8'd226} : s = 188;
	{8'd150,8'd227} : s = 349;
	{8'd150,8'd228} : s = 347;
	{8'd150,8'd229} : s = 475;
	{8'd150,8'd230} : s = 343;
	{8'd150,8'd231} : s = 471;
	{8'd150,8'd232} : s = 463;
	{8'd150,8'd233} : s = 509;
	{8'd150,8'd234} : s = 3;
	{8'd150,8'd235} : s = 22;
	{8'd150,8'd236} : s = 21;
	{8'd150,8'd237} : s = 85;
	{8'd150,8'd238} : s = 19;
	{8'd150,8'd239} : s = 83;
	{8'd150,8'd240} : s = 78;
	{8'd150,8'd241} : s = 186;
	{8'd150,8'd242} : s = 14;
	{8'd150,8'd243} : s = 77;
	{8'd150,8'd244} : s = 75;
	{8'd150,8'd245} : s = 185;
	{8'd150,8'd246} : s = 71;
	{8'd150,8'd247} : s = 182;
	{8'd150,8'd248} : s = 181;
	{8'd150,8'd249} : s = 335;
	{8'd150,8'd250} : s = 13;
	{8'd150,8'd251} : s = 60;
	{8'd150,8'd252} : s = 58;
	{8'd150,8'd253} : s = 179;
	{8'd150,8'd254} : s = 57;
	{8'd150,8'd255} : s = 174;
	{8'd151,8'd0} : s = 422;
	{8'd151,8'd1} : s = 138;
	{8'd151,8'd2} : s = 297;
	{8'd151,8'd3} : s = 294;
	{8'd151,8'd4} : s = 421;
	{8'd151,8'd5} : s = 293;
	{8'd151,8'd6} : s = 419;
	{8'd151,8'd7} : s = 412;
	{8'd151,8'd8} : s = 486;
	{8'd151,8'd9} : s = 24;
	{8'd151,8'd10} : s = 137;
	{8'd151,8'd11} : s = 134;
	{8'd151,8'd12} : s = 291;
	{8'd151,8'd13} : s = 133;
	{8'd151,8'd14} : s = 284;
	{8'd151,8'd15} : s = 282;
	{8'd151,8'd16} : s = 410;
	{8'd151,8'd17} : s = 131;
	{8'd151,8'd18} : s = 281;
	{8'd151,8'd19} : s = 278;
	{8'd151,8'd20} : s = 409;
	{8'd151,8'd21} : s = 277;
	{8'd151,8'd22} : s = 406;
	{8'd151,8'd23} : s = 405;
	{8'd151,8'd24} : s = 485;
	{8'd151,8'd25} : s = 112;
	{8'd151,8'd26} : s = 275;
	{8'd151,8'd27} : s = 270;
	{8'd151,8'd28} : s = 403;
	{8'd151,8'd29} : s = 269;
	{8'd151,8'd30} : s = 398;
	{8'd151,8'd31} : s = 397;
	{8'd151,8'd32} : s = 483;
	{8'd151,8'd33} : s = 267;
	{8'd151,8'd34} : s = 395;
	{8'd151,8'd35} : s = 391;
	{8'd151,8'd36} : s = 476;
	{8'd151,8'd37} : s = 376;
	{8'd151,8'd38} : s = 474;
	{8'd151,8'd39} : s = 473;
	{8'd151,8'd40} : s = 506;
	{8'd151,8'd41} : s = 20;
	{8'd151,8'd42} : s = 104;
	{8'd151,8'd43} : s = 100;
	{8'd151,8'd44} : s = 263;
	{8'd151,8'd45} : s = 98;
	{8'd151,8'd46} : s = 240;
	{8'd151,8'd47} : s = 232;
	{8'd151,8'd48} : s = 372;
	{8'd151,8'd49} : s = 97;
	{8'd151,8'd50} : s = 228;
	{8'd151,8'd51} : s = 226;
	{8'd151,8'd52} : s = 370;
	{8'd151,8'd53} : s = 225;
	{8'd151,8'd54} : s = 369;
	{8'd151,8'd55} : s = 364;
	{8'd151,8'd56} : s = 470;
	{8'd151,8'd57} : s = 88;
	{8'd151,8'd58} : s = 216;
	{8'd151,8'd59} : s = 212;
	{8'd151,8'd60} : s = 362;
	{8'd151,8'd61} : s = 210;
	{8'd151,8'd62} : s = 361;
	{8'd151,8'd63} : s = 358;
	{8'd151,8'd64} : s = 469;
	{8'd151,8'd65} : s = 209;
	{8'd151,8'd66} : s = 357;
	{8'd151,8'd67} : s = 355;
	{8'd151,8'd68} : s = 467;
	{8'd151,8'd69} : s = 348;
	{8'd151,8'd70} : s = 462;
	{8'd151,8'd71} : s = 461;
	{8'd151,8'd72} : s = 505;
	{8'd151,8'd73} : s = 84;
	{8'd151,8'd74} : s = 204;
	{8'd151,8'd75} : s = 202;
	{8'd151,8'd76} : s = 346;
	{8'd151,8'd77} : s = 201;
	{8'd151,8'd78} : s = 345;
	{8'd151,8'd79} : s = 342;
	{8'd151,8'd80} : s = 459;
	{8'd151,8'd81} : s = 198;
	{8'd151,8'd82} : s = 341;
	{8'd151,8'd83} : s = 339;
	{8'd151,8'd84} : s = 455;
	{8'd151,8'd85} : s = 334;
	{8'd151,8'd86} : s = 444;
	{8'd151,8'd87} : s = 442;
	{8'd151,8'd88} : s = 502;
	{8'd151,8'd89} : s = 197;
	{8'd151,8'd90} : s = 333;
	{8'd151,8'd91} : s = 331;
	{8'd151,8'd92} : s = 441;
	{8'd151,8'd93} : s = 327;
	{8'd151,8'd94} : s = 438;
	{8'd151,8'd95} : s = 437;
	{8'd151,8'd96} : s = 501;
	{8'd151,8'd97} : s = 316;
	{8'd151,8'd98} : s = 435;
	{8'd151,8'd99} : s = 430;
	{8'd151,8'd100} : s = 499;
	{8'd151,8'd101} : s = 429;
	{8'd151,8'd102} : s = 494;
	{8'd151,8'd103} : s = 493;
	{8'd151,8'd104} : s = 510;
	{8'd151,8'd105} : s = 1;
	{8'd151,8'd106} : s = 18;
	{8'd151,8'd107} : s = 17;
	{8'd151,8'd108} : s = 82;
	{8'd151,8'd109} : s = 12;
	{8'd151,8'd110} : s = 81;
	{8'd151,8'd111} : s = 76;
	{8'd151,8'd112} : s = 195;
	{8'd151,8'd113} : s = 10;
	{8'd151,8'd114} : s = 74;
	{8'd151,8'd115} : s = 73;
	{8'd151,8'd116} : s = 184;
	{8'd151,8'd117} : s = 70;
	{8'd151,8'd118} : s = 180;
	{8'd151,8'd119} : s = 178;
	{8'd151,8'd120} : s = 314;
	{8'd151,8'd121} : s = 9;
	{8'd151,8'd122} : s = 69;
	{8'd151,8'd123} : s = 67;
	{8'd151,8'd124} : s = 177;
	{8'd151,8'd125} : s = 56;
	{8'd151,8'd126} : s = 172;
	{8'd151,8'd127} : s = 170;
	{8'd151,8'd128} : s = 313;
	{8'd151,8'd129} : s = 52;
	{8'd151,8'd130} : s = 169;
	{8'd151,8'd131} : s = 166;
	{8'd151,8'd132} : s = 310;
	{8'd151,8'd133} : s = 165;
	{8'd151,8'd134} : s = 309;
	{8'd151,8'd135} : s = 307;
	{8'd151,8'd136} : s = 427;
	{8'd151,8'd137} : s = 6;
	{8'd151,8'd138} : s = 50;
	{8'd151,8'd139} : s = 49;
	{8'd151,8'd140} : s = 163;
	{8'd151,8'd141} : s = 44;
	{8'd151,8'd142} : s = 156;
	{8'd151,8'd143} : s = 154;
	{8'd151,8'd144} : s = 302;
	{8'd151,8'd145} : s = 42;
	{8'd151,8'd146} : s = 153;
	{8'd151,8'd147} : s = 150;
	{8'd151,8'd148} : s = 301;
	{8'd151,8'd149} : s = 149;
	{8'd151,8'd150} : s = 299;
	{8'd151,8'd151} : s = 295;
	{8'd151,8'd152} : s = 423;
	{8'd151,8'd153} : s = 41;
	{8'd151,8'd154} : s = 147;
	{8'd151,8'd155} : s = 142;
	{8'd151,8'd156} : s = 286;
	{8'd151,8'd157} : s = 141;
	{8'd151,8'd158} : s = 285;
	{8'd151,8'd159} : s = 283;
	{8'd151,8'd160} : s = 414;
	{8'd151,8'd161} : s = 139;
	{8'd151,8'd162} : s = 279;
	{8'd151,8'd163} : s = 271;
	{8'd151,8'd164} : s = 413;
	{8'd151,8'd165} : s = 248;
	{8'd151,8'd166} : s = 411;
	{8'd151,8'd167} : s = 407;
	{8'd151,8'd168} : s = 491;
	{8'd151,8'd169} : s = 5;
	{8'd151,8'd170} : s = 38;
	{8'd151,8'd171} : s = 37;
	{8'd151,8'd172} : s = 135;
	{8'd151,8'd173} : s = 35;
	{8'd151,8'd174} : s = 120;
	{8'd151,8'd175} : s = 116;
	{8'd151,8'd176} : s = 244;
	{8'd151,8'd177} : s = 28;
	{8'd151,8'd178} : s = 114;
	{8'd151,8'd179} : s = 113;
	{8'd151,8'd180} : s = 242;
	{8'd151,8'd181} : s = 108;
	{8'd151,8'd182} : s = 241;
	{8'd151,8'd183} : s = 236;
	{8'd151,8'd184} : s = 399;
	{8'd151,8'd185} : s = 26;
	{8'd151,8'd186} : s = 106;
	{8'd151,8'd187} : s = 105;
	{8'd151,8'd188} : s = 234;
	{8'd151,8'd189} : s = 102;
	{8'd151,8'd190} : s = 233;
	{8'd151,8'd191} : s = 230;
	{8'd151,8'd192} : s = 380;
	{8'd151,8'd193} : s = 101;
	{8'd151,8'd194} : s = 229;
	{8'd151,8'd195} : s = 227;
	{8'd151,8'd196} : s = 378;
	{8'd151,8'd197} : s = 220;
	{8'd151,8'd198} : s = 377;
	{8'd151,8'd199} : s = 374;
	{8'd151,8'd200} : s = 487;
	{8'd151,8'd201} : s = 25;
	{8'd151,8'd202} : s = 99;
	{8'd151,8'd203} : s = 92;
	{8'd151,8'd204} : s = 218;
	{8'd151,8'd205} : s = 90;
	{8'd151,8'd206} : s = 217;
	{8'd151,8'd207} : s = 214;
	{8'd151,8'd208} : s = 373;
	{8'd151,8'd209} : s = 89;
	{8'd151,8'd210} : s = 213;
	{8'd151,8'd211} : s = 211;
	{8'd151,8'd212} : s = 371;
	{8'd151,8'd213} : s = 206;
	{8'd151,8'd214} : s = 366;
	{8'd151,8'd215} : s = 365;
	{8'd151,8'd216} : s = 478;
	{8'd151,8'd217} : s = 86;
	{8'd151,8'd218} : s = 205;
	{8'd151,8'd219} : s = 203;
	{8'd151,8'd220} : s = 363;
	{8'd151,8'd221} : s = 199;
	{8'd151,8'd222} : s = 359;
	{8'd151,8'd223} : s = 350;
	{8'd151,8'd224} : s = 477;
	{8'd151,8'd225} : s = 188;
	{8'd151,8'd226} : s = 349;
	{8'd151,8'd227} : s = 347;
	{8'd151,8'd228} : s = 475;
	{8'd151,8'd229} : s = 343;
	{8'd151,8'd230} : s = 471;
	{8'd151,8'd231} : s = 463;
	{8'd151,8'd232} : s = 509;
	{8'd151,8'd233} : s = 3;
	{8'd151,8'd234} : s = 22;
	{8'd151,8'd235} : s = 21;
	{8'd151,8'd236} : s = 85;
	{8'd151,8'd237} : s = 19;
	{8'd151,8'd238} : s = 83;
	{8'd151,8'd239} : s = 78;
	{8'd151,8'd240} : s = 186;
	{8'd151,8'd241} : s = 14;
	{8'd151,8'd242} : s = 77;
	{8'd151,8'd243} : s = 75;
	{8'd151,8'd244} : s = 185;
	{8'd151,8'd245} : s = 71;
	{8'd151,8'd246} : s = 182;
	{8'd151,8'd247} : s = 181;
	{8'd151,8'd248} : s = 335;
	{8'd151,8'd249} : s = 13;
	{8'd151,8'd250} : s = 60;
	{8'd151,8'd251} : s = 58;
	{8'd151,8'd252} : s = 179;
	{8'd151,8'd253} : s = 57;
	{8'd151,8'd254} : s = 174;
	{8'd151,8'd255} : s = 173;
	{8'd152,8'd0} : s = 138;
	{8'd152,8'd1} : s = 297;
	{8'd152,8'd2} : s = 294;
	{8'd152,8'd3} : s = 421;
	{8'd152,8'd4} : s = 293;
	{8'd152,8'd5} : s = 419;
	{8'd152,8'd6} : s = 412;
	{8'd152,8'd7} : s = 486;
	{8'd152,8'd8} : s = 24;
	{8'd152,8'd9} : s = 137;
	{8'd152,8'd10} : s = 134;
	{8'd152,8'd11} : s = 291;
	{8'd152,8'd12} : s = 133;
	{8'd152,8'd13} : s = 284;
	{8'd152,8'd14} : s = 282;
	{8'd152,8'd15} : s = 410;
	{8'd152,8'd16} : s = 131;
	{8'd152,8'd17} : s = 281;
	{8'd152,8'd18} : s = 278;
	{8'd152,8'd19} : s = 409;
	{8'd152,8'd20} : s = 277;
	{8'd152,8'd21} : s = 406;
	{8'd152,8'd22} : s = 405;
	{8'd152,8'd23} : s = 485;
	{8'd152,8'd24} : s = 112;
	{8'd152,8'd25} : s = 275;
	{8'd152,8'd26} : s = 270;
	{8'd152,8'd27} : s = 403;
	{8'd152,8'd28} : s = 269;
	{8'd152,8'd29} : s = 398;
	{8'd152,8'd30} : s = 397;
	{8'd152,8'd31} : s = 483;
	{8'd152,8'd32} : s = 267;
	{8'd152,8'd33} : s = 395;
	{8'd152,8'd34} : s = 391;
	{8'd152,8'd35} : s = 476;
	{8'd152,8'd36} : s = 376;
	{8'd152,8'd37} : s = 474;
	{8'd152,8'd38} : s = 473;
	{8'd152,8'd39} : s = 506;
	{8'd152,8'd40} : s = 20;
	{8'd152,8'd41} : s = 104;
	{8'd152,8'd42} : s = 100;
	{8'd152,8'd43} : s = 263;
	{8'd152,8'd44} : s = 98;
	{8'd152,8'd45} : s = 240;
	{8'd152,8'd46} : s = 232;
	{8'd152,8'd47} : s = 372;
	{8'd152,8'd48} : s = 97;
	{8'd152,8'd49} : s = 228;
	{8'd152,8'd50} : s = 226;
	{8'd152,8'd51} : s = 370;
	{8'd152,8'd52} : s = 225;
	{8'd152,8'd53} : s = 369;
	{8'd152,8'd54} : s = 364;
	{8'd152,8'd55} : s = 470;
	{8'd152,8'd56} : s = 88;
	{8'd152,8'd57} : s = 216;
	{8'd152,8'd58} : s = 212;
	{8'd152,8'd59} : s = 362;
	{8'd152,8'd60} : s = 210;
	{8'd152,8'd61} : s = 361;
	{8'd152,8'd62} : s = 358;
	{8'd152,8'd63} : s = 469;
	{8'd152,8'd64} : s = 209;
	{8'd152,8'd65} : s = 357;
	{8'd152,8'd66} : s = 355;
	{8'd152,8'd67} : s = 467;
	{8'd152,8'd68} : s = 348;
	{8'd152,8'd69} : s = 462;
	{8'd152,8'd70} : s = 461;
	{8'd152,8'd71} : s = 505;
	{8'd152,8'd72} : s = 84;
	{8'd152,8'd73} : s = 204;
	{8'd152,8'd74} : s = 202;
	{8'd152,8'd75} : s = 346;
	{8'd152,8'd76} : s = 201;
	{8'd152,8'd77} : s = 345;
	{8'd152,8'd78} : s = 342;
	{8'd152,8'd79} : s = 459;
	{8'd152,8'd80} : s = 198;
	{8'd152,8'd81} : s = 341;
	{8'd152,8'd82} : s = 339;
	{8'd152,8'd83} : s = 455;
	{8'd152,8'd84} : s = 334;
	{8'd152,8'd85} : s = 444;
	{8'd152,8'd86} : s = 442;
	{8'd152,8'd87} : s = 502;
	{8'd152,8'd88} : s = 197;
	{8'd152,8'd89} : s = 333;
	{8'd152,8'd90} : s = 331;
	{8'd152,8'd91} : s = 441;
	{8'd152,8'd92} : s = 327;
	{8'd152,8'd93} : s = 438;
	{8'd152,8'd94} : s = 437;
	{8'd152,8'd95} : s = 501;
	{8'd152,8'd96} : s = 316;
	{8'd152,8'd97} : s = 435;
	{8'd152,8'd98} : s = 430;
	{8'd152,8'd99} : s = 499;
	{8'd152,8'd100} : s = 429;
	{8'd152,8'd101} : s = 494;
	{8'd152,8'd102} : s = 493;
	{8'd152,8'd103} : s = 510;
	{8'd152,8'd104} : s = 1;
	{8'd152,8'd105} : s = 18;
	{8'd152,8'd106} : s = 17;
	{8'd152,8'd107} : s = 82;
	{8'd152,8'd108} : s = 12;
	{8'd152,8'd109} : s = 81;
	{8'd152,8'd110} : s = 76;
	{8'd152,8'd111} : s = 195;
	{8'd152,8'd112} : s = 10;
	{8'd152,8'd113} : s = 74;
	{8'd152,8'd114} : s = 73;
	{8'd152,8'd115} : s = 184;
	{8'd152,8'd116} : s = 70;
	{8'd152,8'd117} : s = 180;
	{8'd152,8'd118} : s = 178;
	{8'd152,8'd119} : s = 314;
	{8'd152,8'd120} : s = 9;
	{8'd152,8'd121} : s = 69;
	{8'd152,8'd122} : s = 67;
	{8'd152,8'd123} : s = 177;
	{8'd152,8'd124} : s = 56;
	{8'd152,8'd125} : s = 172;
	{8'd152,8'd126} : s = 170;
	{8'd152,8'd127} : s = 313;
	{8'd152,8'd128} : s = 52;
	{8'd152,8'd129} : s = 169;
	{8'd152,8'd130} : s = 166;
	{8'd152,8'd131} : s = 310;
	{8'd152,8'd132} : s = 165;
	{8'd152,8'd133} : s = 309;
	{8'd152,8'd134} : s = 307;
	{8'd152,8'd135} : s = 427;
	{8'd152,8'd136} : s = 6;
	{8'd152,8'd137} : s = 50;
	{8'd152,8'd138} : s = 49;
	{8'd152,8'd139} : s = 163;
	{8'd152,8'd140} : s = 44;
	{8'd152,8'd141} : s = 156;
	{8'd152,8'd142} : s = 154;
	{8'd152,8'd143} : s = 302;
	{8'd152,8'd144} : s = 42;
	{8'd152,8'd145} : s = 153;
	{8'd152,8'd146} : s = 150;
	{8'd152,8'd147} : s = 301;
	{8'd152,8'd148} : s = 149;
	{8'd152,8'd149} : s = 299;
	{8'd152,8'd150} : s = 295;
	{8'd152,8'd151} : s = 423;
	{8'd152,8'd152} : s = 41;
	{8'd152,8'd153} : s = 147;
	{8'd152,8'd154} : s = 142;
	{8'd152,8'd155} : s = 286;
	{8'd152,8'd156} : s = 141;
	{8'd152,8'd157} : s = 285;
	{8'd152,8'd158} : s = 283;
	{8'd152,8'd159} : s = 414;
	{8'd152,8'd160} : s = 139;
	{8'd152,8'd161} : s = 279;
	{8'd152,8'd162} : s = 271;
	{8'd152,8'd163} : s = 413;
	{8'd152,8'd164} : s = 248;
	{8'd152,8'd165} : s = 411;
	{8'd152,8'd166} : s = 407;
	{8'd152,8'd167} : s = 491;
	{8'd152,8'd168} : s = 5;
	{8'd152,8'd169} : s = 38;
	{8'd152,8'd170} : s = 37;
	{8'd152,8'd171} : s = 135;
	{8'd152,8'd172} : s = 35;
	{8'd152,8'd173} : s = 120;
	{8'd152,8'd174} : s = 116;
	{8'd152,8'd175} : s = 244;
	{8'd152,8'd176} : s = 28;
	{8'd152,8'd177} : s = 114;
	{8'd152,8'd178} : s = 113;
	{8'd152,8'd179} : s = 242;
	{8'd152,8'd180} : s = 108;
	{8'd152,8'd181} : s = 241;
	{8'd152,8'd182} : s = 236;
	{8'd152,8'd183} : s = 399;
	{8'd152,8'd184} : s = 26;
	{8'd152,8'd185} : s = 106;
	{8'd152,8'd186} : s = 105;
	{8'd152,8'd187} : s = 234;
	{8'd152,8'd188} : s = 102;
	{8'd152,8'd189} : s = 233;
	{8'd152,8'd190} : s = 230;
	{8'd152,8'd191} : s = 380;
	{8'd152,8'd192} : s = 101;
	{8'd152,8'd193} : s = 229;
	{8'd152,8'd194} : s = 227;
	{8'd152,8'd195} : s = 378;
	{8'd152,8'd196} : s = 220;
	{8'd152,8'd197} : s = 377;
	{8'd152,8'd198} : s = 374;
	{8'd152,8'd199} : s = 487;
	{8'd152,8'd200} : s = 25;
	{8'd152,8'd201} : s = 99;
	{8'd152,8'd202} : s = 92;
	{8'd152,8'd203} : s = 218;
	{8'd152,8'd204} : s = 90;
	{8'd152,8'd205} : s = 217;
	{8'd152,8'd206} : s = 214;
	{8'd152,8'd207} : s = 373;
	{8'd152,8'd208} : s = 89;
	{8'd152,8'd209} : s = 213;
	{8'd152,8'd210} : s = 211;
	{8'd152,8'd211} : s = 371;
	{8'd152,8'd212} : s = 206;
	{8'd152,8'd213} : s = 366;
	{8'd152,8'd214} : s = 365;
	{8'd152,8'd215} : s = 478;
	{8'd152,8'd216} : s = 86;
	{8'd152,8'd217} : s = 205;
	{8'd152,8'd218} : s = 203;
	{8'd152,8'd219} : s = 363;
	{8'd152,8'd220} : s = 199;
	{8'd152,8'd221} : s = 359;
	{8'd152,8'd222} : s = 350;
	{8'd152,8'd223} : s = 477;
	{8'd152,8'd224} : s = 188;
	{8'd152,8'd225} : s = 349;
	{8'd152,8'd226} : s = 347;
	{8'd152,8'd227} : s = 475;
	{8'd152,8'd228} : s = 343;
	{8'd152,8'd229} : s = 471;
	{8'd152,8'd230} : s = 463;
	{8'd152,8'd231} : s = 509;
	{8'd152,8'd232} : s = 3;
	{8'd152,8'd233} : s = 22;
	{8'd152,8'd234} : s = 21;
	{8'd152,8'd235} : s = 85;
	{8'd152,8'd236} : s = 19;
	{8'd152,8'd237} : s = 83;
	{8'd152,8'd238} : s = 78;
	{8'd152,8'd239} : s = 186;
	{8'd152,8'd240} : s = 14;
	{8'd152,8'd241} : s = 77;
	{8'd152,8'd242} : s = 75;
	{8'd152,8'd243} : s = 185;
	{8'd152,8'd244} : s = 71;
	{8'd152,8'd245} : s = 182;
	{8'd152,8'd246} : s = 181;
	{8'd152,8'd247} : s = 335;
	{8'd152,8'd248} : s = 13;
	{8'd152,8'd249} : s = 60;
	{8'd152,8'd250} : s = 58;
	{8'd152,8'd251} : s = 179;
	{8'd152,8'd252} : s = 57;
	{8'd152,8'd253} : s = 174;
	{8'd152,8'd254} : s = 173;
	{8'd152,8'd255} : s = 318;
	{8'd153,8'd0} : s = 297;
	{8'd153,8'd1} : s = 294;
	{8'd153,8'd2} : s = 421;
	{8'd153,8'd3} : s = 293;
	{8'd153,8'd4} : s = 419;
	{8'd153,8'd5} : s = 412;
	{8'd153,8'd6} : s = 486;
	{8'd153,8'd7} : s = 24;
	{8'd153,8'd8} : s = 137;
	{8'd153,8'd9} : s = 134;
	{8'd153,8'd10} : s = 291;
	{8'd153,8'd11} : s = 133;
	{8'd153,8'd12} : s = 284;
	{8'd153,8'd13} : s = 282;
	{8'd153,8'd14} : s = 410;
	{8'd153,8'd15} : s = 131;
	{8'd153,8'd16} : s = 281;
	{8'd153,8'd17} : s = 278;
	{8'd153,8'd18} : s = 409;
	{8'd153,8'd19} : s = 277;
	{8'd153,8'd20} : s = 406;
	{8'd153,8'd21} : s = 405;
	{8'd153,8'd22} : s = 485;
	{8'd153,8'd23} : s = 112;
	{8'd153,8'd24} : s = 275;
	{8'd153,8'd25} : s = 270;
	{8'd153,8'd26} : s = 403;
	{8'd153,8'd27} : s = 269;
	{8'd153,8'd28} : s = 398;
	{8'd153,8'd29} : s = 397;
	{8'd153,8'd30} : s = 483;
	{8'd153,8'd31} : s = 267;
	{8'd153,8'd32} : s = 395;
	{8'd153,8'd33} : s = 391;
	{8'd153,8'd34} : s = 476;
	{8'd153,8'd35} : s = 376;
	{8'd153,8'd36} : s = 474;
	{8'd153,8'd37} : s = 473;
	{8'd153,8'd38} : s = 506;
	{8'd153,8'd39} : s = 20;
	{8'd153,8'd40} : s = 104;
	{8'd153,8'd41} : s = 100;
	{8'd153,8'd42} : s = 263;
	{8'd153,8'd43} : s = 98;
	{8'd153,8'd44} : s = 240;
	{8'd153,8'd45} : s = 232;
	{8'd153,8'd46} : s = 372;
	{8'd153,8'd47} : s = 97;
	{8'd153,8'd48} : s = 228;
	{8'd153,8'd49} : s = 226;
	{8'd153,8'd50} : s = 370;
	{8'd153,8'd51} : s = 225;
	{8'd153,8'd52} : s = 369;
	{8'd153,8'd53} : s = 364;
	{8'd153,8'd54} : s = 470;
	{8'd153,8'd55} : s = 88;
	{8'd153,8'd56} : s = 216;
	{8'd153,8'd57} : s = 212;
	{8'd153,8'd58} : s = 362;
	{8'd153,8'd59} : s = 210;
	{8'd153,8'd60} : s = 361;
	{8'd153,8'd61} : s = 358;
	{8'd153,8'd62} : s = 469;
	{8'd153,8'd63} : s = 209;
	{8'd153,8'd64} : s = 357;
	{8'd153,8'd65} : s = 355;
	{8'd153,8'd66} : s = 467;
	{8'd153,8'd67} : s = 348;
	{8'd153,8'd68} : s = 462;
	{8'd153,8'd69} : s = 461;
	{8'd153,8'd70} : s = 505;
	{8'd153,8'd71} : s = 84;
	{8'd153,8'd72} : s = 204;
	{8'd153,8'd73} : s = 202;
	{8'd153,8'd74} : s = 346;
	{8'd153,8'd75} : s = 201;
	{8'd153,8'd76} : s = 345;
	{8'd153,8'd77} : s = 342;
	{8'd153,8'd78} : s = 459;
	{8'd153,8'd79} : s = 198;
	{8'd153,8'd80} : s = 341;
	{8'd153,8'd81} : s = 339;
	{8'd153,8'd82} : s = 455;
	{8'd153,8'd83} : s = 334;
	{8'd153,8'd84} : s = 444;
	{8'd153,8'd85} : s = 442;
	{8'd153,8'd86} : s = 502;
	{8'd153,8'd87} : s = 197;
	{8'd153,8'd88} : s = 333;
	{8'd153,8'd89} : s = 331;
	{8'd153,8'd90} : s = 441;
	{8'd153,8'd91} : s = 327;
	{8'd153,8'd92} : s = 438;
	{8'd153,8'd93} : s = 437;
	{8'd153,8'd94} : s = 501;
	{8'd153,8'd95} : s = 316;
	{8'd153,8'd96} : s = 435;
	{8'd153,8'd97} : s = 430;
	{8'd153,8'd98} : s = 499;
	{8'd153,8'd99} : s = 429;
	{8'd153,8'd100} : s = 494;
	{8'd153,8'd101} : s = 493;
	{8'd153,8'd102} : s = 510;
	{8'd153,8'd103} : s = 1;
	{8'd153,8'd104} : s = 18;
	{8'd153,8'd105} : s = 17;
	{8'd153,8'd106} : s = 82;
	{8'd153,8'd107} : s = 12;
	{8'd153,8'd108} : s = 81;
	{8'd153,8'd109} : s = 76;
	{8'd153,8'd110} : s = 195;
	{8'd153,8'd111} : s = 10;
	{8'd153,8'd112} : s = 74;
	{8'd153,8'd113} : s = 73;
	{8'd153,8'd114} : s = 184;
	{8'd153,8'd115} : s = 70;
	{8'd153,8'd116} : s = 180;
	{8'd153,8'd117} : s = 178;
	{8'd153,8'd118} : s = 314;
	{8'd153,8'd119} : s = 9;
	{8'd153,8'd120} : s = 69;
	{8'd153,8'd121} : s = 67;
	{8'd153,8'd122} : s = 177;
	{8'd153,8'd123} : s = 56;
	{8'd153,8'd124} : s = 172;
	{8'd153,8'd125} : s = 170;
	{8'd153,8'd126} : s = 313;
	{8'd153,8'd127} : s = 52;
	{8'd153,8'd128} : s = 169;
	{8'd153,8'd129} : s = 166;
	{8'd153,8'd130} : s = 310;
	{8'd153,8'd131} : s = 165;
	{8'd153,8'd132} : s = 309;
	{8'd153,8'd133} : s = 307;
	{8'd153,8'd134} : s = 427;
	{8'd153,8'd135} : s = 6;
	{8'd153,8'd136} : s = 50;
	{8'd153,8'd137} : s = 49;
	{8'd153,8'd138} : s = 163;
	{8'd153,8'd139} : s = 44;
	{8'd153,8'd140} : s = 156;
	{8'd153,8'd141} : s = 154;
	{8'd153,8'd142} : s = 302;
	{8'd153,8'd143} : s = 42;
	{8'd153,8'd144} : s = 153;
	{8'd153,8'd145} : s = 150;
	{8'd153,8'd146} : s = 301;
	{8'd153,8'd147} : s = 149;
	{8'd153,8'd148} : s = 299;
	{8'd153,8'd149} : s = 295;
	{8'd153,8'd150} : s = 423;
	{8'd153,8'd151} : s = 41;
	{8'd153,8'd152} : s = 147;
	{8'd153,8'd153} : s = 142;
	{8'd153,8'd154} : s = 286;
	{8'd153,8'd155} : s = 141;
	{8'd153,8'd156} : s = 285;
	{8'd153,8'd157} : s = 283;
	{8'd153,8'd158} : s = 414;
	{8'd153,8'd159} : s = 139;
	{8'd153,8'd160} : s = 279;
	{8'd153,8'd161} : s = 271;
	{8'd153,8'd162} : s = 413;
	{8'd153,8'd163} : s = 248;
	{8'd153,8'd164} : s = 411;
	{8'd153,8'd165} : s = 407;
	{8'd153,8'd166} : s = 491;
	{8'd153,8'd167} : s = 5;
	{8'd153,8'd168} : s = 38;
	{8'd153,8'd169} : s = 37;
	{8'd153,8'd170} : s = 135;
	{8'd153,8'd171} : s = 35;
	{8'd153,8'd172} : s = 120;
	{8'd153,8'd173} : s = 116;
	{8'd153,8'd174} : s = 244;
	{8'd153,8'd175} : s = 28;
	{8'd153,8'd176} : s = 114;
	{8'd153,8'd177} : s = 113;
	{8'd153,8'd178} : s = 242;
	{8'd153,8'd179} : s = 108;
	{8'd153,8'd180} : s = 241;
	{8'd153,8'd181} : s = 236;
	{8'd153,8'd182} : s = 399;
	{8'd153,8'd183} : s = 26;
	{8'd153,8'd184} : s = 106;
	{8'd153,8'd185} : s = 105;
	{8'd153,8'd186} : s = 234;
	{8'd153,8'd187} : s = 102;
	{8'd153,8'd188} : s = 233;
	{8'd153,8'd189} : s = 230;
	{8'd153,8'd190} : s = 380;
	{8'd153,8'd191} : s = 101;
	{8'd153,8'd192} : s = 229;
	{8'd153,8'd193} : s = 227;
	{8'd153,8'd194} : s = 378;
	{8'd153,8'd195} : s = 220;
	{8'd153,8'd196} : s = 377;
	{8'd153,8'd197} : s = 374;
	{8'd153,8'd198} : s = 487;
	{8'd153,8'd199} : s = 25;
	{8'd153,8'd200} : s = 99;
	{8'd153,8'd201} : s = 92;
	{8'd153,8'd202} : s = 218;
	{8'd153,8'd203} : s = 90;
	{8'd153,8'd204} : s = 217;
	{8'd153,8'd205} : s = 214;
	{8'd153,8'd206} : s = 373;
	{8'd153,8'd207} : s = 89;
	{8'd153,8'd208} : s = 213;
	{8'd153,8'd209} : s = 211;
	{8'd153,8'd210} : s = 371;
	{8'd153,8'd211} : s = 206;
	{8'd153,8'd212} : s = 366;
	{8'd153,8'd213} : s = 365;
	{8'd153,8'd214} : s = 478;
	{8'd153,8'd215} : s = 86;
	{8'd153,8'd216} : s = 205;
	{8'd153,8'd217} : s = 203;
	{8'd153,8'd218} : s = 363;
	{8'd153,8'd219} : s = 199;
	{8'd153,8'd220} : s = 359;
	{8'd153,8'd221} : s = 350;
	{8'd153,8'd222} : s = 477;
	{8'd153,8'd223} : s = 188;
	{8'd153,8'd224} : s = 349;
	{8'd153,8'd225} : s = 347;
	{8'd153,8'd226} : s = 475;
	{8'd153,8'd227} : s = 343;
	{8'd153,8'd228} : s = 471;
	{8'd153,8'd229} : s = 463;
	{8'd153,8'd230} : s = 509;
	{8'd153,8'd231} : s = 3;
	{8'd153,8'd232} : s = 22;
	{8'd153,8'd233} : s = 21;
	{8'd153,8'd234} : s = 85;
	{8'd153,8'd235} : s = 19;
	{8'd153,8'd236} : s = 83;
	{8'd153,8'd237} : s = 78;
	{8'd153,8'd238} : s = 186;
	{8'd153,8'd239} : s = 14;
	{8'd153,8'd240} : s = 77;
	{8'd153,8'd241} : s = 75;
	{8'd153,8'd242} : s = 185;
	{8'd153,8'd243} : s = 71;
	{8'd153,8'd244} : s = 182;
	{8'd153,8'd245} : s = 181;
	{8'd153,8'd246} : s = 335;
	{8'd153,8'd247} : s = 13;
	{8'd153,8'd248} : s = 60;
	{8'd153,8'd249} : s = 58;
	{8'd153,8'd250} : s = 179;
	{8'd153,8'd251} : s = 57;
	{8'd153,8'd252} : s = 174;
	{8'd153,8'd253} : s = 173;
	{8'd153,8'd254} : s = 318;
	{8'd153,8'd255} : s = 54;
	{8'd154,8'd0} : s = 294;
	{8'd154,8'd1} : s = 421;
	{8'd154,8'd2} : s = 293;
	{8'd154,8'd3} : s = 419;
	{8'd154,8'd4} : s = 412;
	{8'd154,8'd5} : s = 486;
	{8'd154,8'd6} : s = 24;
	{8'd154,8'd7} : s = 137;
	{8'd154,8'd8} : s = 134;
	{8'd154,8'd9} : s = 291;
	{8'd154,8'd10} : s = 133;
	{8'd154,8'd11} : s = 284;
	{8'd154,8'd12} : s = 282;
	{8'd154,8'd13} : s = 410;
	{8'd154,8'd14} : s = 131;
	{8'd154,8'd15} : s = 281;
	{8'd154,8'd16} : s = 278;
	{8'd154,8'd17} : s = 409;
	{8'd154,8'd18} : s = 277;
	{8'd154,8'd19} : s = 406;
	{8'd154,8'd20} : s = 405;
	{8'd154,8'd21} : s = 485;
	{8'd154,8'd22} : s = 112;
	{8'd154,8'd23} : s = 275;
	{8'd154,8'd24} : s = 270;
	{8'd154,8'd25} : s = 403;
	{8'd154,8'd26} : s = 269;
	{8'd154,8'd27} : s = 398;
	{8'd154,8'd28} : s = 397;
	{8'd154,8'd29} : s = 483;
	{8'd154,8'd30} : s = 267;
	{8'd154,8'd31} : s = 395;
	{8'd154,8'd32} : s = 391;
	{8'd154,8'd33} : s = 476;
	{8'd154,8'd34} : s = 376;
	{8'd154,8'd35} : s = 474;
	{8'd154,8'd36} : s = 473;
	{8'd154,8'd37} : s = 506;
	{8'd154,8'd38} : s = 20;
	{8'd154,8'd39} : s = 104;
	{8'd154,8'd40} : s = 100;
	{8'd154,8'd41} : s = 263;
	{8'd154,8'd42} : s = 98;
	{8'd154,8'd43} : s = 240;
	{8'd154,8'd44} : s = 232;
	{8'd154,8'd45} : s = 372;
	{8'd154,8'd46} : s = 97;
	{8'd154,8'd47} : s = 228;
	{8'd154,8'd48} : s = 226;
	{8'd154,8'd49} : s = 370;
	{8'd154,8'd50} : s = 225;
	{8'd154,8'd51} : s = 369;
	{8'd154,8'd52} : s = 364;
	{8'd154,8'd53} : s = 470;
	{8'd154,8'd54} : s = 88;
	{8'd154,8'd55} : s = 216;
	{8'd154,8'd56} : s = 212;
	{8'd154,8'd57} : s = 362;
	{8'd154,8'd58} : s = 210;
	{8'd154,8'd59} : s = 361;
	{8'd154,8'd60} : s = 358;
	{8'd154,8'd61} : s = 469;
	{8'd154,8'd62} : s = 209;
	{8'd154,8'd63} : s = 357;
	{8'd154,8'd64} : s = 355;
	{8'd154,8'd65} : s = 467;
	{8'd154,8'd66} : s = 348;
	{8'd154,8'd67} : s = 462;
	{8'd154,8'd68} : s = 461;
	{8'd154,8'd69} : s = 505;
	{8'd154,8'd70} : s = 84;
	{8'd154,8'd71} : s = 204;
	{8'd154,8'd72} : s = 202;
	{8'd154,8'd73} : s = 346;
	{8'd154,8'd74} : s = 201;
	{8'd154,8'd75} : s = 345;
	{8'd154,8'd76} : s = 342;
	{8'd154,8'd77} : s = 459;
	{8'd154,8'd78} : s = 198;
	{8'd154,8'd79} : s = 341;
	{8'd154,8'd80} : s = 339;
	{8'd154,8'd81} : s = 455;
	{8'd154,8'd82} : s = 334;
	{8'd154,8'd83} : s = 444;
	{8'd154,8'd84} : s = 442;
	{8'd154,8'd85} : s = 502;
	{8'd154,8'd86} : s = 197;
	{8'd154,8'd87} : s = 333;
	{8'd154,8'd88} : s = 331;
	{8'd154,8'd89} : s = 441;
	{8'd154,8'd90} : s = 327;
	{8'd154,8'd91} : s = 438;
	{8'd154,8'd92} : s = 437;
	{8'd154,8'd93} : s = 501;
	{8'd154,8'd94} : s = 316;
	{8'd154,8'd95} : s = 435;
	{8'd154,8'd96} : s = 430;
	{8'd154,8'd97} : s = 499;
	{8'd154,8'd98} : s = 429;
	{8'd154,8'd99} : s = 494;
	{8'd154,8'd100} : s = 493;
	{8'd154,8'd101} : s = 510;
	{8'd154,8'd102} : s = 1;
	{8'd154,8'd103} : s = 18;
	{8'd154,8'd104} : s = 17;
	{8'd154,8'd105} : s = 82;
	{8'd154,8'd106} : s = 12;
	{8'd154,8'd107} : s = 81;
	{8'd154,8'd108} : s = 76;
	{8'd154,8'd109} : s = 195;
	{8'd154,8'd110} : s = 10;
	{8'd154,8'd111} : s = 74;
	{8'd154,8'd112} : s = 73;
	{8'd154,8'd113} : s = 184;
	{8'd154,8'd114} : s = 70;
	{8'd154,8'd115} : s = 180;
	{8'd154,8'd116} : s = 178;
	{8'd154,8'd117} : s = 314;
	{8'd154,8'd118} : s = 9;
	{8'd154,8'd119} : s = 69;
	{8'd154,8'd120} : s = 67;
	{8'd154,8'd121} : s = 177;
	{8'd154,8'd122} : s = 56;
	{8'd154,8'd123} : s = 172;
	{8'd154,8'd124} : s = 170;
	{8'd154,8'd125} : s = 313;
	{8'd154,8'd126} : s = 52;
	{8'd154,8'd127} : s = 169;
	{8'd154,8'd128} : s = 166;
	{8'd154,8'd129} : s = 310;
	{8'd154,8'd130} : s = 165;
	{8'd154,8'd131} : s = 309;
	{8'd154,8'd132} : s = 307;
	{8'd154,8'd133} : s = 427;
	{8'd154,8'd134} : s = 6;
	{8'd154,8'd135} : s = 50;
	{8'd154,8'd136} : s = 49;
	{8'd154,8'd137} : s = 163;
	{8'd154,8'd138} : s = 44;
	{8'd154,8'd139} : s = 156;
	{8'd154,8'd140} : s = 154;
	{8'd154,8'd141} : s = 302;
	{8'd154,8'd142} : s = 42;
	{8'd154,8'd143} : s = 153;
	{8'd154,8'd144} : s = 150;
	{8'd154,8'd145} : s = 301;
	{8'd154,8'd146} : s = 149;
	{8'd154,8'd147} : s = 299;
	{8'd154,8'd148} : s = 295;
	{8'd154,8'd149} : s = 423;
	{8'd154,8'd150} : s = 41;
	{8'd154,8'd151} : s = 147;
	{8'd154,8'd152} : s = 142;
	{8'd154,8'd153} : s = 286;
	{8'd154,8'd154} : s = 141;
	{8'd154,8'd155} : s = 285;
	{8'd154,8'd156} : s = 283;
	{8'd154,8'd157} : s = 414;
	{8'd154,8'd158} : s = 139;
	{8'd154,8'd159} : s = 279;
	{8'd154,8'd160} : s = 271;
	{8'd154,8'd161} : s = 413;
	{8'd154,8'd162} : s = 248;
	{8'd154,8'd163} : s = 411;
	{8'd154,8'd164} : s = 407;
	{8'd154,8'd165} : s = 491;
	{8'd154,8'd166} : s = 5;
	{8'd154,8'd167} : s = 38;
	{8'd154,8'd168} : s = 37;
	{8'd154,8'd169} : s = 135;
	{8'd154,8'd170} : s = 35;
	{8'd154,8'd171} : s = 120;
	{8'd154,8'd172} : s = 116;
	{8'd154,8'd173} : s = 244;
	{8'd154,8'd174} : s = 28;
	{8'd154,8'd175} : s = 114;
	{8'd154,8'd176} : s = 113;
	{8'd154,8'd177} : s = 242;
	{8'd154,8'd178} : s = 108;
	{8'd154,8'd179} : s = 241;
	{8'd154,8'd180} : s = 236;
	{8'd154,8'd181} : s = 399;
	{8'd154,8'd182} : s = 26;
	{8'd154,8'd183} : s = 106;
	{8'd154,8'd184} : s = 105;
	{8'd154,8'd185} : s = 234;
	{8'd154,8'd186} : s = 102;
	{8'd154,8'd187} : s = 233;
	{8'd154,8'd188} : s = 230;
	{8'd154,8'd189} : s = 380;
	{8'd154,8'd190} : s = 101;
	{8'd154,8'd191} : s = 229;
	{8'd154,8'd192} : s = 227;
	{8'd154,8'd193} : s = 378;
	{8'd154,8'd194} : s = 220;
	{8'd154,8'd195} : s = 377;
	{8'd154,8'd196} : s = 374;
	{8'd154,8'd197} : s = 487;
	{8'd154,8'd198} : s = 25;
	{8'd154,8'd199} : s = 99;
	{8'd154,8'd200} : s = 92;
	{8'd154,8'd201} : s = 218;
	{8'd154,8'd202} : s = 90;
	{8'd154,8'd203} : s = 217;
	{8'd154,8'd204} : s = 214;
	{8'd154,8'd205} : s = 373;
	{8'd154,8'd206} : s = 89;
	{8'd154,8'd207} : s = 213;
	{8'd154,8'd208} : s = 211;
	{8'd154,8'd209} : s = 371;
	{8'd154,8'd210} : s = 206;
	{8'd154,8'd211} : s = 366;
	{8'd154,8'd212} : s = 365;
	{8'd154,8'd213} : s = 478;
	{8'd154,8'd214} : s = 86;
	{8'd154,8'd215} : s = 205;
	{8'd154,8'd216} : s = 203;
	{8'd154,8'd217} : s = 363;
	{8'd154,8'd218} : s = 199;
	{8'd154,8'd219} : s = 359;
	{8'd154,8'd220} : s = 350;
	{8'd154,8'd221} : s = 477;
	{8'd154,8'd222} : s = 188;
	{8'd154,8'd223} : s = 349;
	{8'd154,8'd224} : s = 347;
	{8'd154,8'd225} : s = 475;
	{8'd154,8'd226} : s = 343;
	{8'd154,8'd227} : s = 471;
	{8'd154,8'd228} : s = 463;
	{8'd154,8'd229} : s = 509;
	{8'd154,8'd230} : s = 3;
	{8'd154,8'd231} : s = 22;
	{8'd154,8'd232} : s = 21;
	{8'd154,8'd233} : s = 85;
	{8'd154,8'd234} : s = 19;
	{8'd154,8'd235} : s = 83;
	{8'd154,8'd236} : s = 78;
	{8'd154,8'd237} : s = 186;
	{8'd154,8'd238} : s = 14;
	{8'd154,8'd239} : s = 77;
	{8'd154,8'd240} : s = 75;
	{8'd154,8'd241} : s = 185;
	{8'd154,8'd242} : s = 71;
	{8'd154,8'd243} : s = 182;
	{8'd154,8'd244} : s = 181;
	{8'd154,8'd245} : s = 335;
	{8'd154,8'd246} : s = 13;
	{8'd154,8'd247} : s = 60;
	{8'd154,8'd248} : s = 58;
	{8'd154,8'd249} : s = 179;
	{8'd154,8'd250} : s = 57;
	{8'd154,8'd251} : s = 174;
	{8'd154,8'd252} : s = 173;
	{8'd154,8'd253} : s = 318;
	{8'd154,8'd254} : s = 54;
	{8'd154,8'd255} : s = 171;
	{8'd155,8'd0} : s = 421;
	{8'd155,8'd1} : s = 293;
	{8'd155,8'd2} : s = 419;
	{8'd155,8'd3} : s = 412;
	{8'd155,8'd4} : s = 486;
	{8'd155,8'd5} : s = 24;
	{8'd155,8'd6} : s = 137;
	{8'd155,8'd7} : s = 134;
	{8'd155,8'd8} : s = 291;
	{8'd155,8'd9} : s = 133;
	{8'd155,8'd10} : s = 284;
	{8'd155,8'd11} : s = 282;
	{8'd155,8'd12} : s = 410;
	{8'd155,8'd13} : s = 131;
	{8'd155,8'd14} : s = 281;
	{8'd155,8'd15} : s = 278;
	{8'd155,8'd16} : s = 409;
	{8'd155,8'd17} : s = 277;
	{8'd155,8'd18} : s = 406;
	{8'd155,8'd19} : s = 405;
	{8'd155,8'd20} : s = 485;
	{8'd155,8'd21} : s = 112;
	{8'd155,8'd22} : s = 275;
	{8'd155,8'd23} : s = 270;
	{8'd155,8'd24} : s = 403;
	{8'd155,8'd25} : s = 269;
	{8'd155,8'd26} : s = 398;
	{8'd155,8'd27} : s = 397;
	{8'd155,8'd28} : s = 483;
	{8'd155,8'd29} : s = 267;
	{8'd155,8'd30} : s = 395;
	{8'd155,8'd31} : s = 391;
	{8'd155,8'd32} : s = 476;
	{8'd155,8'd33} : s = 376;
	{8'd155,8'd34} : s = 474;
	{8'd155,8'd35} : s = 473;
	{8'd155,8'd36} : s = 506;
	{8'd155,8'd37} : s = 20;
	{8'd155,8'd38} : s = 104;
	{8'd155,8'd39} : s = 100;
	{8'd155,8'd40} : s = 263;
	{8'd155,8'd41} : s = 98;
	{8'd155,8'd42} : s = 240;
	{8'd155,8'd43} : s = 232;
	{8'd155,8'd44} : s = 372;
	{8'd155,8'd45} : s = 97;
	{8'd155,8'd46} : s = 228;
	{8'd155,8'd47} : s = 226;
	{8'd155,8'd48} : s = 370;
	{8'd155,8'd49} : s = 225;
	{8'd155,8'd50} : s = 369;
	{8'd155,8'd51} : s = 364;
	{8'd155,8'd52} : s = 470;
	{8'd155,8'd53} : s = 88;
	{8'd155,8'd54} : s = 216;
	{8'd155,8'd55} : s = 212;
	{8'd155,8'd56} : s = 362;
	{8'd155,8'd57} : s = 210;
	{8'd155,8'd58} : s = 361;
	{8'd155,8'd59} : s = 358;
	{8'd155,8'd60} : s = 469;
	{8'd155,8'd61} : s = 209;
	{8'd155,8'd62} : s = 357;
	{8'd155,8'd63} : s = 355;
	{8'd155,8'd64} : s = 467;
	{8'd155,8'd65} : s = 348;
	{8'd155,8'd66} : s = 462;
	{8'd155,8'd67} : s = 461;
	{8'd155,8'd68} : s = 505;
	{8'd155,8'd69} : s = 84;
	{8'd155,8'd70} : s = 204;
	{8'd155,8'd71} : s = 202;
	{8'd155,8'd72} : s = 346;
	{8'd155,8'd73} : s = 201;
	{8'd155,8'd74} : s = 345;
	{8'd155,8'd75} : s = 342;
	{8'd155,8'd76} : s = 459;
	{8'd155,8'd77} : s = 198;
	{8'd155,8'd78} : s = 341;
	{8'd155,8'd79} : s = 339;
	{8'd155,8'd80} : s = 455;
	{8'd155,8'd81} : s = 334;
	{8'd155,8'd82} : s = 444;
	{8'd155,8'd83} : s = 442;
	{8'd155,8'd84} : s = 502;
	{8'd155,8'd85} : s = 197;
	{8'd155,8'd86} : s = 333;
	{8'd155,8'd87} : s = 331;
	{8'd155,8'd88} : s = 441;
	{8'd155,8'd89} : s = 327;
	{8'd155,8'd90} : s = 438;
	{8'd155,8'd91} : s = 437;
	{8'd155,8'd92} : s = 501;
	{8'd155,8'd93} : s = 316;
	{8'd155,8'd94} : s = 435;
	{8'd155,8'd95} : s = 430;
	{8'd155,8'd96} : s = 499;
	{8'd155,8'd97} : s = 429;
	{8'd155,8'd98} : s = 494;
	{8'd155,8'd99} : s = 493;
	{8'd155,8'd100} : s = 510;
	{8'd155,8'd101} : s = 1;
	{8'd155,8'd102} : s = 18;
	{8'd155,8'd103} : s = 17;
	{8'd155,8'd104} : s = 82;
	{8'd155,8'd105} : s = 12;
	{8'd155,8'd106} : s = 81;
	{8'd155,8'd107} : s = 76;
	{8'd155,8'd108} : s = 195;
	{8'd155,8'd109} : s = 10;
	{8'd155,8'd110} : s = 74;
	{8'd155,8'd111} : s = 73;
	{8'd155,8'd112} : s = 184;
	{8'd155,8'd113} : s = 70;
	{8'd155,8'd114} : s = 180;
	{8'd155,8'd115} : s = 178;
	{8'd155,8'd116} : s = 314;
	{8'd155,8'd117} : s = 9;
	{8'd155,8'd118} : s = 69;
	{8'd155,8'd119} : s = 67;
	{8'd155,8'd120} : s = 177;
	{8'd155,8'd121} : s = 56;
	{8'd155,8'd122} : s = 172;
	{8'd155,8'd123} : s = 170;
	{8'd155,8'd124} : s = 313;
	{8'd155,8'd125} : s = 52;
	{8'd155,8'd126} : s = 169;
	{8'd155,8'd127} : s = 166;
	{8'd155,8'd128} : s = 310;
	{8'd155,8'd129} : s = 165;
	{8'd155,8'd130} : s = 309;
	{8'd155,8'd131} : s = 307;
	{8'd155,8'd132} : s = 427;
	{8'd155,8'd133} : s = 6;
	{8'd155,8'd134} : s = 50;
	{8'd155,8'd135} : s = 49;
	{8'd155,8'd136} : s = 163;
	{8'd155,8'd137} : s = 44;
	{8'd155,8'd138} : s = 156;
	{8'd155,8'd139} : s = 154;
	{8'd155,8'd140} : s = 302;
	{8'd155,8'd141} : s = 42;
	{8'd155,8'd142} : s = 153;
	{8'd155,8'd143} : s = 150;
	{8'd155,8'd144} : s = 301;
	{8'd155,8'd145} : s = 149;
	{8'd155,8'd146} : s = 299;
	{8'd155,8'd147} : s = 295;
	{8'd155,8'd148} : s = 423;
	{8'd155,8'd149} : s = 41;
	{8'd155,8'd150} : s = 147;
	{8'd155,8'd151} : s = 142;
	{8'd155,8'd152} : s = 286;
	{8'd155,8'd153} : s = 141;
	{8'd155,8'd154} : s = 285;
	{8'd155,8'd155} : s = 283;
	{8'd155,8'd156} : s = 414;
	{8'd155,8'd157} : s = 139;
	{8'd155,8'd158} : s = 279;
	{8'd155,8'd159} : s = 271;
	{8'd155,8'd160} : s = 413;
	{8'd155,8'd161} : s = 248;
	{8'd155,8'd162} : s = 411;
	{8'd155,8'd163} : s = 407;
	{8'd155,8'd164} : s = 491;
	{8'd155,8'd165} : s = 5;
	{8'd155,8'd166} : s = 38;
	{8'd155,8'd167} : s = 37;
	{8'd155,8'd168} : s = 135;
	{8'd155,8'd169} : s = 35;
	{8'd155,8'd170} : s = 120;
	{8'd155,8'd171} : s = 116;
	{8'd155,8'd172} : s = 244;
	{8'd155,8'd173} : s = 28;
	{8'd155,8'd174} : s = 114;
	{8'd155,8'd175} : s = 113;
	{8'd155,8'd176} : s = 242;
	{8'd155,8'd177} : s = 108;
	{8'd155,8'd178} : s = 241;
	{8'd155,8'd179} : s = 236;
	{8'd155,8'd180} : s = 399;
	{8'd155,8'd181} : s = 26;
	{8'd155,8'd182} : s = 106;
	{8'd155,8'd183} : s = 105;
	{8'd155,8'd184} : s = 234;
	{8'd155,8'd185} : s = 102;
	{8'd155,8'd186} : s = 233;
	{8'd155,8'd187} : s = 230;
	{8'd155,8'd188} : s = 380;
	{8'd155,8'd189} : s = 101;
	{8'd155,8'd190} : s = 229;
	{8'd155,8'd191} : s = 227;
	{8'd155,8'd192} : s = 378;
	{8'd155,8'd193} : s = 220;
	{8'd155,8'd194} : s = 377;
	{8'd155,8'd195} : s = 374;
	{8'd155,8'd196} : s = 487;
	{8'd155,8'd197} : s = 25;
	{8'd155,8'd198} : s = 99;
	{8'd155,8'd199} : s = 92;
	{8'd155,8'd200} : s = 218;
	{8'd155,8'd201} : s = 90;
	{8'd155,8'd202} : s = 217;
	{8'd155,8'd203} : s = 214;
	{8'd155,8'd204} : s = 373;
	{8'd155,8'd205} : s = 89;
	{8'd155,8'd206} : s = 213;
	{8'd155,8'd207} : s = 211;
	{8'd155,8'd208} : s = 371;
	{8'd155,8'd209} : s = 206;
	{8'd155,8'd210} : s = 366;
	{8'd155,8'd211} : s = 365;
	{8'd155,8'd212} : s = 478;
	{8'd155,8'd213} : s = 86;
	{8'd155,8'd214} : s = 205;
	{8'd155,8'd215} : s = 203;
	{8'd155,8'd216} : s = 363;
	{8'd155,8'd217} : s = 199;
	{8'd155,8'd218} : s = 359;
	{8'd155,8'd219} : s = 350;
	{8'd155,8'd220} : s = 477;
	{8'd155,8'd221} : s = 188;
	{8'd155,8'd222} : s = 349;
	{8'd155,8'd223} : s = 347;
	{8'd155,8'd224} : s = 475;
	{8'd155,8'd225} : s = 343;
	{8'd155,8'd226} : s = 471;
	{8'd155,8'd227} : s = 463;
	{8'd155,8'd228} : s = 509;
	{8'd155,8'd229} : s = 3;
	{8'd155,8'd230} : s = 22;
	{8'd155,8'd231} : s = 21;
	{8'd155,8'd232} : s = 85;
	{8'd155,8'd233} : s = 19;
	{8'd155,8'd234} : s = 83;
	{8'd155,8'd235} : s = 78;
	{8'd155,8'd236} : s = 186;
	{8'd155,8'd237} : s = 14;
	{8'd155,8'd238} : s = 77;
	{8'd155,8'd239} : s = 75;
	{8'd155,8'd240} : s = 185;
	{8'd155,8'd241} : s = 71;
	{8'd155,8'd242} : s = 182;
	{8'd155,8'd243} : s = 181;
	{8'd155,8'd244} : s = 335;
	{8'd155,8'd245} : s = 13;
	{8'd155,8'd246} : s = 60;
	{8'd155,8'd247} : s = 58;
	{8'd155,8'd248} : s = 179;
	{8'd155,8'd249} : s = 57;
	{8'd155,8'd250} : s = 174;
	{8'd155,8'd251} : s = 173;
	{8'd155,8'd252} : s = 318;
	{8'd155,8'd253} : s = 54;
	{8'd155,8'd254} : s = 171;
	{8'd155,8'd255} : s = 167;
	{8'd156,8'd0} : s = 293;
	{8'd156,8'd1} : s = 419;
	{8'd156,8'd2} : s = 412;
	{8'd156,8'd3} : s = 486;
	{8'd156,8'd4} : s = 24;
	{8'd156,8'd5} : s = 137;
	{8'd156,8'd6} : s = 134;
	{8'd156,8'd7} : s = 291;
	{8'd156,8'd8} : s = 133;
	{8'd156,8'd9} : s = 284;
	{8'd156,8'd10} : s = 282;
	{8'd156,8'd11} : s = 410;
	{8'd156,8'd12} : s = 131;
	{8'd156,8'd13} : s = 281;
	{8'd156,8'd14} : s = 278;
	{8'd156,8'd15} : s = 409;
	{8'd156,8'd16} : s = 277;
	{8'd156,8'd17} : s = 406;
	{8'd156,8'd18} : s = 405;
	{8'd156,8'd19} : s = 485;
	{8'd156,8'd20} : s = 112;
	{8'd156,8'd21} : s = 275;
	{8'd156,8'd22} : s = 270;
	{8'd156,8'd23} : s = 403;
	{8'd156,8'd24} : s = 269;
	{8'd156,8'd25} : s = 398;
	{8'd156,8'd26} : s = 397;
	{8'd156,8'd27} : s = 483;
	{8'd156,8'd28} : s = 267;
	{8'd156,8'd29} : s = 395;
	{8'd156,8'd30} : s = 391;
	{8'd156,8'd31} : s = 476;
	{8'd156,8'd32} : s = 376;
	{8'd156,8'd33} : s = 474;
	{8'd156,8'd34} : s = 473;
	{8'd156,8'd35} : s = 506;
	{8'd156,8'd36} : s = 20;
	{8'd156,8'd37} : s = 104;
	{8'd156,8'd38} : s = 100;
	{8'd156,8'd39} : s = 263;
	{8'd156,8'd40} : s = 98;
	{8'd156,8'd41} : s = 240;
	{8'd156,8'd42} : s = 232;
	{8'd156,8'd43} : s = 372;
	{8'd156,8'd44} : s = 97;
	{8'd156,8'd45} : s = 228;
	{8'd156,8'd46} : s = 226;
	{8'd156,8'd47} : s = 370;
	{8'd156,8'd48} : s = 225;
	{8'd156,8'd49} : s = 369;
	{8'd156,8'd50} : s = 364;
	{8'd156,8'd51} : s = 470;
	{8'd156,8'd52} : s = 88;
	{8'd156,8'd53} : s = 216;
	{8'd156,8'd54} : s = 212;
	{8'd156,8'd55} : s = 362;
	{8'd156,8'd56} : s = 210;
	{8'd156,8'd57} : s = 361;
	{8'd156,8'd58} : s = 358;
	{8'd156,8'd59} : s = 469;
	{8'd156,8'd60} : s = 209;
	{8'd156,8'd61} : s = 357;
	{8'd156,8'd62} : s = 355;
	{8'd156,8'd63} : s = 467;
	{8'd156,8'd64} : s = 348;
	{8'd156,8'd65} : s = 462;
	{8'd156,8'd66} : s = 461;
	{8'd156,8'd67} : s = 505;
	{8'd156,8'd68} : s = 84;
	{8'd156,8'd69} : s = 204;
	{8'd156,8'd70} : s = 202;
	{8'd156,8'd71} : s = 346;
	{8'd156,8'd72} : s = 201;
	{8'd156,8'd73} : s = 345;
	{8'd156,8'd74} : s = 342;
	{8'd156,8'd75} : s = 459;
	{8'd156,8'd76} : s = 198;
	{8'd156,8'd77} : s = 341;
	{8'd156,8'd78} : s = 339;
	{8'd156,8'd79} : s = 455;
	{8'd156,8'd80} : s = 334;
	{8'd156,8'd81} : s = 444;
	{8'd156,8'd82} : s = 442;
	{8'd156,8'd83} : s = 502;
	{8'd156,8'd84} : s = 197;
	{8'd156,8'd85} : s = 333;
	{8'd156,8'd86} : s = 331;
	{8'd156,8'd87} : s = 441;
	{8'd156,8'd88} : s = 327;
	{8'd156,8'd89} : s = 438;
	{8'd156,8'd90} : s = 437;
	{8'd156,8'd91} : s = 501;
	{8'd156,8'd92} : s = 316;
	{8'd156,8'd93} : s = 435;
	{8'd156,8'd94} : s = 430;
	{8'd156,8'd95} : s = 499;
	{8'd156,8'd96} : s = 429;
	{8'd156,8'd97} : s = 494;
	{8'd156,8'd98} : s = 493;
	{8'd156,8'd99} : s = 510;
	{8'd156,8'd100} : s = 1;
	{8'd156,8'd101} : s = 18;
	{8'd156,8'd102} : s = 17;
	{8'd156,8'd103} : s = 82;
	{8'd156,8'd104} : s = 12;
	{8'd156,8'd105} : s = 81;
	{8'd156,8'd106} : s = 76;
	{8'd156,8'd107} : s = 195;
	{8'd156,8'd108} : s = 10;
	{8'd156,8'd109} : s = 74;
	{8'd156,8'd110} : s = 73;
	{8'd156,8'd111} : s = 184;
	{8'd156,8'd112} : s = 70;
	{8'd156,8'd113} : s = 180;
	{8'd156,8'd114} : s = 178;
	{8'd156,8'd115} : s = 314;
	{8'd156,8'd116} : s = 9;
	{8'd156,8'd117} : s = 69;
	{8'd156,8'd118} : s = 67;
	{8'd156,8'd119} : s = 177;
	{8'd156,8'd120} : s = 56;
	{8'd156,8'd121} : s = 172;
	{8'd156,8'd122} : s = 170;
	{8'd156,8'd123} : s = 313;
	{8'd156,8'd124} : s = 52;
	{8'd156,8'd125} : s = 169;
	{8'd156,8'd126} : s = 166;
	{8'd156,8'd127} : s = 310;
	{8'd156,8'd128} : s = 165;
	{8'd156,8'd129} : s = 309;
	{8'd156,8'd130} : s = 307;
	{8'd156,8'd131} : s = 427;
	{8'd156,8'd132} : s = 6;
	{8'd156,8'd133} : s = 50;
	{8'd156,8'd134} : s = 49;
	{8'd156,8'd135} : s = 163;
	{8'd156,8'd136} : s = 44;
	{8'd156,8'd137} : s = 156;
	{8'd156,8'd138} : s = 154;
	{8'd156,8'd139} : s = 302;
	{8'd156,8'd140} : s = 42;
	{8'd156,8'd141} : s = 153;
	{8'd156,8'd142} : s = 150;
	{8'd156,8'd143} : s = 301;
	{8'd156,8'd144} : s = 149;
	{8'd156,8'd145} : s = 299;
	{8'd156,8'd146} : s = 295;
	{8'd156,8'd147} : s = 423;
	{8'd156,8'd148} : s = 41;
	{8'd156,8'd149} : s = 147;
	{8'd156,8'd150} : s = 142;
	{8'd156,8'd151} : s = 286;
	{8'd156,8'd152} : s = 141;
	{8'd156,8'd153} : s = 285;
	{8'd156,8'd154} : s = 283;
	{8'd156,8'd155} : s = 414;
	{8'd156,8'd156} : s = 139;
	{8'd156,8'd157} : s = 279;
	{8'd156,8'd158} : s = 271;
	{8'd156,8'd159} : s = 413;
	{8'd156,8'd160} : s = 248;
	{8'd156,8'd161} : s = 411;
	{8'd156,8'd162} : s = 407;
	{8'd156,8'd163} : s = 491;
	{8'd156,8'd164} : s = 5;
	{8'd156,8'd165} : s = 38;
	{8'd156,8'd166} : s = 37;
	{8'd156,8'd167} : s = 135;
	{8'd156,8'd168} : s = 35;
	{8'd156,8'd169} : s = 120;
	{8'd156,8'd170} : s = 116;
	{8'd156,8'd171} : s = 244;
	{8'd156,8'd172} : s = 28;
	{8'd156,8'd173} : s = 114;
	{8'd156,8'd174} : s = 113;
	{8'd156,8'd175} : s = 242;
	{8'd156,8'd176} : s = 108;
	{8'd156,8'd177} : s = 241;
	{8'd156,8'd178} : s = 236;
	{8'd156,8'd179} : s = 399;
	{8'd156,8'd180} : s = 26;
	{8'd156,8'd181} : s = 106;
	{8'd156,8'd182} : s = 105;
	{8'd156,8'd183} : s = 234;
	{8'd156,8'd184} : s = 102;
	{8'd156,8'd185} : s = 233;
	{8'd156,8'd186} : s = 230;
	{8'd156,8'd187} : s = 380;
	{8'd156,8'd188} : s = 101;
	{8'd156,8'd189} : s = 229;
	{8'd156,8'd190} : s = 227;
	{8'd156,8'd191} : s = 378;
	{8'd156,8'd192} : s = 220;
	{8'd156,8'd193} : s = 377;
	{8'd156,8'd194} : s = 374;
	{8'd156,8'd195} : s = 487;
	{8'd156,8'd196} : s = 25;
	{8'd156,8'd197} : s = 99;
	{8'd156,8'd198} : s = 92;
	{8'd156,8'd199} : s = 218;
	{8'd156,8'd200} : s = 90;
	{8'd156,8'd201} : s = 217;
	{8'd156,8'd202} : s = 214;
	{8'd156,8'd203} : s = 373;
	{8'd156,8'd204} : s = 89;
	{8'd156,8'd205} : s = 213;
	{8'd156,8'd206} : s = 211;
	{8'd156,8'd207} : s = 371;
	{8'd156,8'd208} : s = 206;
	{8'd156,8'd209} : s = 366;
	{8'd156,8'd210} : s = 365;
	{8'd156,8'd211} : s = 478;
	{8'd156,8'd212} : s = 86;
	{8'd156,8'd213} : s = 205;
	{8'd156,8'd214} : s = 203;
	{8'd156,8'd215} : s = 363;
	{8'd156,8'd216} : s = 199;
	{8'd156,8'd217} : s = 359;
	{8'd156,8'd218} : s = 350;
	{8'd156,8'd219} : s = 477;
	{8'd156,8'd220} : s = 188;
	{8'd156,8'd221} : s = 349;
	{8'd156,8'd222} : s = 347;
	{8'd156,8'd223} : s = 475;
	{8'd156,8'd224} : s = 343;
	{8'd156,8'd225} : s = 471;
	{8'd156,8'd226} : s = 463;
	{8'd156,8'd227} : s = 509;
	{8'd156,8'd228} : s = 3;
	{8'd156,8'd229} : s = 22;
	{8'd156,8'd230} : s = 21;
	{8'd156,8'd231} : s = 85;
	{8'd156,8'd232} : s = 19;
	{8'd156,8'd233} : s = 83;
	{8'd156,8'd234} : s = 78;
	{8'd156,8'd235} : s = 186;
	{8'd156,8'd236} : s = 14;
	{8'd156,8'd237} : s = 77;
	{8'd156,8'd238} : s = 75;
	{8'd156,8'd239} : s = 185;
	{8'd156,8'd240} : s = 71;
	{8'd156,8'd241} : s = 182;
	{8'd156,8'd242} : s = 181;
	{8'd156,8'd243} : s = 335;
	{8'd156,8'd244} : s = 13;
	{8'd156,8'd245} : s = 60;
	{8'd156,8'd246} : s = 58;
	{8'd156,8'd247} : s = 179;
	{8'd156,8'd248} : s = 57;
	{8'd156,8'd249} : s = 174;
	{8'd156,8'd250} : s = 173;
	{8'd156,8'd251} : s = 318;
	{8'd156,8'd252} : s = 54;
	{8'd156,8'd253} : s = 171;
	{8'd156,8'd254} : s = 167;
	{8'd156,8'd255} : s = 317;
	{8'd157,8'd0} : s = 419;
	{8'd157,8'd1} : s = 412;
	{8'd157,8'd2} : s = 486;
	{8'd157,8'd3} : s = 24;
	{8'd157,8'd4} : s = 137;
	{8'd157,8'd5} : s = 134;
	{8'd157,8'd6} : s = 291;
	{8'd157,8'd7} : s = 133;
	{8'd157,8'd8} : s = 284;
	{8'd157,8'd9} : s = 282;
	{8'd157,8'd10} : s = 410;
	{8'd157,8'd11} : s = 131;
	{8'd157,8'd12} : s = 281;
	{8'd157,8'd13} : s = 278;
	{8'd157,8'd14} : s = 409;
	{8'd157,8'd15} : s = 277;
	{8'd157,8'd16} : s = 406;
	{8'd157,8'd17} : s = 405;
	{8'd157,8'd18} : s = 485;
	{8'd157,8'd19} : s = 112;
	{8'd157,8'd20} : s = 275;
	{8'd157,8'd21} : s = 270;
	{8'd157,8'd22} : s = 403;
	{8'd157,8'd23} : s = 269;
	{8'd157,8'd24} : s = 398;
	{8'd157,8'd25} : s = 397;
	{8'd157,8'd26} : s = 483;
	{8'd157,8'd27} : s = 267;
	{8'd157,8'd28} : s = 395;
	{8'd157,8'd29} : s = 391;
	{8'd157,8'd30} : s = 476;
	{8'd157,8'd31} : s = 376;
	{8'd157,8'd32} : s = 474;
	{8'd157,8'd33} : s = 473;
	{8'd157,8'd34} : s = 506;
	{8'd157,8'd35} : s = 20;
	{8'd157,8'd36} : s = 104;
	{8'd157,8'd37} : s = 100;
	{8'd157,8'd38} : s = 263;
	{8'd157,8'd39} : s = 98;
	{8'd157,8'd40} : s = 240;
	{8'd157,8'd41} : s = 232;
	{8'd157,8'd42} : s = 372;
	{8'd157,8'd43} : s = 97;
	{8'd157,8'd44} : s = 228;
	{8'd157,8'd45} : s = 226;
	{8'd157,8'd46} : s = 370;
	{8'd157,8'd47} : s = 225;
	{8'd157,8'd48} : s = 369;
	{8'd157,8'd49} : s = 364;
	{8'd157,8'd50} : s = 470;
	{8'd157,8'd51} : s = 88;
	{8'd157,8'd52} : s = 216;
	{8'd157,8'd53} : s = 212;
	{8'd157,8'd54} : s = 362;
	{8'd157,8'd55} : s = 210;
	{8'd157,8'd56} : s = 361;
	{8'd157,8'd57} : s = 358;
	{8'd157,8'd58} : s = 469;
	{8'd157,8'd59} : s = 209;
	{8'd157,8'd60} : s = 357;
	{8'd157,8'd61} : s = 355;
	{8'd157,8'd62} : s = 467;
	{8'd157,8'd63} : s = 348;
	{8'd157,8'd64} : s = 462;
	{8'd157,8'd65} : s = 461;
	{8'd157,8'd66} : s = 505;
	{8'd157,8'd67} : s = 84;
	{8'd157,8'd68} : s = 204;
	{8'd157,8'd69} : s = 202;
	{8'd157,8'd70} : s = 346;
	{8'd157,8'd71} : s = 201;
	{8'd157,8'd72} : s = 345;
	{8'd157,8'd73} : s = 342;
	{8'd157,8'd74} : s = 459;
	{8'd157,8'd75} : s = 198;
	{8'd157,8'd76} : s = 341;
	{8'd157,8'd77} : s = 339;
	{8'd157,8'd78} : s = 455;
	{8'd157,8'd79} : s = 334;
	{8'd157,8'd80} : s = 444;
	{8'd157,8'd81} : s = 442;
	{8'd157,8'd82} : s = 502;
	{8'd157,8'd83} : s = 197;
	{8'd157,8'd84} : s = 333;
	{8'd157,8'd85} : s = 331;
	{8'd157,8'd86} : s = 441;
	{8'd157,8'd87} : s = 327;
	{8'd157,8'd88} : s = 438;
	{8'd157,8'd89} : s = 437;
	{8'd157,8'd90} : s = 501;
	{8'd157,8'd91} : s = 316;
	{8'd157,8'd92} : s = 435;
	{8'd157,8'd93} : s = 430;
	{8'd157,8'd94} : s = 499;
	{8'd157,8'd95} : s = 429;
	{8'd157,8'd96} : s = 494;
	{8'd157,8'd97} : s = 493;
	{8'd157,8'd98} : s = 510;
	{8'd157,8'd99} : s = 1;
	{8'd157,8'd100} : s = 18;
	{8'd157,8'd101} : s = 17;
	{8'd157,8'd102} : s = 82;
	{8'd157,8'd103} : s = 12;
	{8'd157,8'd104} : s = 81;
	{8'd157,8'd105} : s = 76;
	{8'd157,8'd106} : s = 195;
	{8'd157,8'd107} : s = 10;
	{8'd157,8'd108} : s = 74;
	{8'd157,8'd109} : s = 73;
	{8'd157,8'd110} : s = 184;
	{8'd157,8'd111} : s = 70;
	{8'd157,8'd112} : s = 180;
	{8'd157,8'd113} : s = 178;
	{8'd157,8'd114} : s = 314;
	{8'd157,8'd115} : s = 9;
	{8'd157,8'd116} : s = 69;
	{8'd157,8'd117} : s = 67;
	{8'd157,8'd118} : s = 177;
	{8'd157,8'd119} : s = 56;
	{8'd157,8'd120} : s = 172;
	{8'd157,8'd121} : s = 170;
	{8'd157,8'd122} : s = 313;
	{8'd157,8'd123} : s = 52;
	{8'd157,8'd124} : s = 169;
	{8'd157,8'd125} : s = 166;
	{8'd157,8'd126} : s = 310;
	{8'd157,8'd127} : s = 165;
	{8'd157,8'd128} : s = 309;
	{8'd157,8'd129} : s = 307;
	{8'd157,8'd130} : s = 427;
	{8'd157,8'd131} : s = 6;
	{8'd157,8'd132} : s = 50;
	{8'd157,8'd133} : s = 49;
	{8'd157,8'd134} : s = 163;
	{8'd157,8'd135} : s = 44;
	{8'd157,8'd136} : s = 156;
	{8'd157,8'd137} : s = 154;
	{8'd157,8'd138} : s = 302;
	{8'd157,8'd139} : s = 42;
	{8'd157,8'd140} : s = 153;
	{8'd157,8'd141} : s = 150;
	{8'd157,8'd142} : s = 301;
	{8'd157,8'd143} : s = 149;
	{8'd157,8'd144} : s = 299;
	{8'd157,8'd145} : s = 295;
	{8'd157,8'd146} : s = 423;
	{8'd157,8'd147} : s = 41;
	{8'd157,8'd148} : s = 147;
	{8'd157,8'd149} : s = 142;
	{8'd157,8'd150} : s = 286;
	{8'd157,8'd151} : s = 141;
	{8'd157,8'd152} : s = 285;
	{8'd157,8'd153} : s = 283;
	{8'd157,8'd154} : s = 414;
	{8'd157,8'd155} : s = 139;
	{8'd157,8'd156} : s = 279;
	{8'd157,8'd157} : s = 271;
	{8'd157,8'd158} : s = 413;
	{8'd157,8'd159} : s = 248;
	{8'd157,8'd160} : s = 411;
	{8'd157,8'd161} : s = 407;
	{8'd157,8'd162} : s = 491;
	{8'd157,8'd163} : s = 5;
	{8'd157,8'd164} : s = 38;
	{8'd157,8'd165} : s = 37;
	{8'd157,8'd166} : s = 135;
	{8'd157,8'd167} : s = 35;
	{8'd157,8'd168} : s = 120;
	{8'd157,8'd169} : s = 116;
	{8'd157,8'd170} : s = 244;
	{8'd157,8'd171} : s = 28;
	{8'd157,8'd172} : s = 114;
	{8'd157,8'd173} : s = 113;
	{8'd157,8'd174} : s = 242;
	{8'd157,8'd175} : s = 108;
	{8'd157,8'd176} : s = 241;
	{8'd157,8'd177} : s = 236;
	{8'd157,8'd178} : s = 399;
	{8'd157,8'd179} : s = 26;
	{8'd157,8'd180} : s = 106;
	{8'd157,8'd181} : s = 105;
	{8'd157,8'd182} : s = 234;
	{8'd157,8'd183} : s = 102;
	{8'd157,8'd184} : s = 233;
	{8'd157,8'd185} : s = 230;
	{8'd157,8'd186} : s = 380;
	{8'd157,8'd187} : s = 101;
	{8'd157,8'd188} : s = 229;
	{8'd157,8'd189} : s = 227;
	{8'd157,8'd190} : s = 378;
	{8'd157,8'd191} : s = 220;
	{8'd157,8'd192} : s = 377;
	{8'd157,8'd193} : s = 374;
	{8'd157,8'd194} : s = 487;
	{8'd157,8'd195} : s = 25;
	{8'd157,8'd196} : s = 99;
	{8'd157,8'd197} : s = 92;
	{8'd157,8'd198} : s = 218;
	{8'd157,8'd199} : s = 90;
	{8'd157,8'd200} : s = 217;
	{8'd157,8'd201} : s = 214;
	{8'd157,8'd202} : s = 373;
	{8'd157,8'd203} : s = 89;
	{8'd157,8'd204} : s = 213;
	{8'd157,8'd205} : s = 211;
	{8'd157,8'd206} : s = 371;
	{8'd157,8'd207} : s = 206;
	{8'd157,8'd208} : s = 366;
	{8'd157,8'd209} : s = 365;
	{8'd157,8'd210} : s = 478;
	{8'd157,8'd211} : s = 86;
	{8'd157,8'd212} : s = 205;
	{8'd157,8'd213} : s = 203;
	{8'd157,8'd214} : s = 363;
	{8'd157,8'd215} : s = 199;
	{8'd157,8'd216} : s = 359;
	{8'd157,8'd217} : s = 350;
	{8'd157,8'd218} : s = 477;
	{8'd157,8'd219} : s = 188;
	{8'd157,8'd220} : s = 349;
	{8'd157,8'd221} : s = 347;
	{8'd157,8'd222} : s = 475;
	{8'd157,8'd223} : s = 343;
	{8'd157,8'd224} : s = 471;
	{8'd157,8'd225} : s = 463;
	{8'd157,8'd226} : s = 509;
	{8'd157,8'd227} : s = 3;
	{8'd157,8'd228} : s = 22;
	{8'd157,8'd229} : s = 21;
	{8'd157,8'd230} : s = 85;
	{8'd157,8'd231} : s = 19;
	{8'd157,8'd232} : s = 83;
	{8'd157,8'd233} : s = 78;
	{8'd157,8'd234} : s = 186;
	{8'd157,8'd235} : s = 14;
	{8'd157,8'd236} : s = 77;
	{8'd157,8'd237} : s = 75;
	{8'd157,8'd238} : s = 185;
	{8'd157,8'd239} : s = 71;
	{8'd157,8'd240} : s = 182;
	{8'd157,8'd241} : s = 181;
	{8'd157,8'd242} : s = 335;
	{8'd157,8'd243} : s = 13;
	{8'd157,8'd244} : s = 60;
	{8'd157,8'd245} : s = 58;
	{8'd157,8'd246} : s = 179;
	{8'd157,8'd247} : s = 57;
	{8'd157,8'd248} : s = 174;
	{8'd157,8'd249} : s = 173;
	{8'd157,8'd250} : s = 318;
	{8'd157,8'd251} : s = 54;
	{8'd157,8'd252} : s = 171;
	{8'd157,8'd253} : s = 167;
	{8'd157,8'd254} : s = 317;
	{8'd157,8'd255} : s = 158;
	{8'd158,8'd0} : s = 412;
	{8'd158,8'd1} : s = 486;
	{8'd158,8'd2} : s = 24;
	{8'd158,8'd3} : s = 137;
	{8'd158,8'd4} : s = 134;
	{8'd158,8'd5} : s = 291;
	{8'd158,8'd6} : s = 133;
	{8'd158,8'd7} : s = 284;
	{8'd158,8'd8} : s = 282;
	{8'd158,8'd9} : s = 410;
	{8'd158,8'd10} : s = 131;
	{8'd158,8'd11} : s = 281;
	{8'd158,8'd12} : s = 278;
	{8'd158,8'd13} : s = 409;
	{8'd158,8'd14} : s = 277;
	{8'd158,8'd15} : s = 406;
	{8'd158,8'd16} : s = 405;
	{8'd158,8'd17} : s = 485;
	{8'd158,8'd18} : s = 112;
	{8'd158,8'd19} : s = 275;
	{8'd158,8'd20} : s = 270;
	{8'd158,8'd21} : s = 403;
	{8'd158,8'd22} : s = 269;
	{8'd158,8'd23} : s = 398;
	{8'd158,8'd24} : s = 397;
	{8'd158,8'd25} : s = 483;
	{8'd158,8'd26} : s = 267;
	{8'd158,8'd27} : s = 395;
	{8'd158,8'd28} : s = 391;
	{8'd158,8'd29} : s = 476;
	{8'd158,8'd30} : s = 376;
	{8'd158,8'd31} : s = 474;
	{8'd158,8'd32} : s = 473;
	{8'd158,8'd33} : s = 506;
	{8'd158,8'd34} : s = 20;
	{8'd158,8'd35} : s = 104;
	{8'd158,8'd36} : s = 100;
	{8'd158,8'd37} : s = 263;
	{8'd158,8'd38} : s = 98;
	{8'd158,8'd39} : s = 240;
	{8'd158,8'd40} : s = 232;
	{8'd158,8'd41} : s = 372;
	{8'd158,8'd42} : s = 97;
	{8'd158,8'd43} : s = 228;
	{8'd158,8'd44} : s = 226;
	{8'd158,8'd45} : s = 370;
	{8'd158,8'd46} : s = 225;
	{8'd158,8'd47} : s = 369;
	{8'd158,8'd48} : s = 364;
	{8'd158,8'd49} : s = 470;
	{8'd158,8'd50} : s = 88;
	{8'd158,8'd51} : s = 216;
	{8'd158,8'd52} : s = 212;
	{8'd158,8'd53} : s = 362;
	{8'd158,8'd54} : s = 210;
	{8'd158,8'd55} : s = 361;
	{8'd158,8'd56} : s = 358;
	{8'd158,8'd57} : s = 469;
	{8'd158,8'd58} : s = 209;
	{8'd158,8'd59} : s = 357;
	{8'd158,8'd60} : s = 355;
	{8'd158,8'd61} : s = 467;
	{8'd158,8'd62} : s = 348;
	{8'd158,8'd63} : s = 462;
	{8'd158,8'd64} : s = 461;
	{8'd158,8'd65} : s = 505;
	{8'd158,8'd66} : s = 84;
	{8'd158,8'd67} : s = 204;
	{8'd158,8'd68} : s = 202;
	{8'd158,8'd69} : s = 346;
	{8'd158,8'd70} : s = 201;
	{8'd158,8'd71} : s = 345;
	{8'd158,8'd72} : s = 342;
	{8'd158,8'd73} : s = 459;
	{8'd158,8'd74} : s = 198;
	{8'd158,8'd75} : s = 341;
	{8'd158,8'd76} : s = 339;
	{8'd158,8'd77} : s = 455;
	{8'd158,8'd78} : s = 334;
	{8'd158,8'd79} : s = 444;
	{8'd158,8'd80} : s = 442;
	{8'd158,8'd81} : s = 502;
	{8'd158,8'd82} : s = 197;
	{8'd158,8'd83} : s = 333;
	{8'd158,8'd84} : s = 331;
	{8'd158,8'd85} : s = 441;
	{8'd158,8'd86} : s = 327;
	{8'd158,8'd87} : s = 438;
	{8'd158,8'd88} : s = 437;
	{8'd158,8'd89} : s = 501;
	{8'd158,8'd90} : s = 316;
	{8'd158,8'd91} : s = 435;
	{8'd158,8'd92} : s = 430;
	{8'd158,8'd93} : s = 499;
	{8'd158,8'd94} : s = 429;
	{8'd158,8'd95} : s = 494;
	{8'd158,8'd96} : s = 493;
	{8'd158,8'd97} : s = 510;
	{8'd158,8'd98} : s = 1;
	{8'd158,8'd99} : s = 18;
	{8'd158,8'd100} : s = 17;
	{8'd158,8'd101} : s = 82;
	{8'd158,8'd102} : s = 12;
	{8'd158,8'd103} : s = 81;
	{8'd158,8'd104} : s = 76;
	{8'd158,8'd105} : s = 195;
	{8'd158,8'd106} : s = 10;
	{8'd158,8'd107} : s = 74;
	{8'd158,8'd108} : s = 73;
	{8'd158,8'd109} : s = 184;
	{8'd158,8'd110} : s = 70;
	{8'd158,8'd111} : s = 180;
	{8'd158,8'd112} : s = 178;
	{8'd158,8'd113} : s = 314;
	{8'd158,8'd114} : s = 9;
	{8'd158,8'd115} : s = 69;
	{8'd158,8'd116} : s = 67;
	{8'd158,8'd117} : s = 177;
	{8'd158,8'd118} : s = 56;
	{8'd158,8'd119} : s = 172;
	{8'd158,8'd120} : s = 170;
	{8'd158,8'd121} : s = 313;
	{8'd158,8'd122} : s = 52;
	{8'd158,8'd123} : s = 169;
	{8'd158,8'd124} : s = 166;
	{8'd158,8'd125} : s = 310;
	{8'd158,8'd126} : s = 165;
	{8'd158,8'd127} : s = 309;
	{8'd158,8'd128} : s = 307;
	{8'd158,8'd129} : s = 427;
	{8'd158,8'd130} : s = 6;
	{8'd158,8'd131} : s = 50;
	{8'd158,8'd132} : s = 49;
	{8'd158,8'd133} : s = 163;
	{8'd158,8'd134} : s = 44;
	{8'd158,8'd135} : s = 156;
	{8'd158,8'd136} : s = 154;
	{8'd158,8'd137} : s = 302;
	{8'd158,8'd138} : s = 42;
	{8'd158,8'd139} : s = 153;
	{8'd158,8'd140} : s = 150;
	{8'd158,8'd141} : s = 301;
	{8'd158,8'd142} : s = 149;
	{8'd158,8'd143} : s = 299;
	{8'd158,8'd144} : s = 295;
	{8'd158,8'd145} : s = 423;
	{8'd158,8'd146} : s = 41;
	{8'd158,8'd147} : s = 147;
	{8'd158,8'd148} : s = 142;
	{8'd158,8'd149} : s = 286;
	{8'd158,8'd150} : s = 141;
	{8'd158,8'd151} : s = 285;
	{8'd158,8'd152} : s = 283;
	{8'd158,8'd153} : s = 414;
	{8'd158,8'd154} : s = 139;
	{8'd158,8'd155} : s = 279;
	{8'd158,8'd156} : s = 271;
	{8'd158,8'd157} : s = 413;
	{8'd158,8'd158} : s = 248;
	{8'd158,8'd159} : s = 411;
	{8'd158,8'd160} : s = 407;
	{8'd158,8'd161} : s = 491;
	{8'd158,8'd162} : s = 5;
	{8'd158,8'd163} : s = 38;
	{8'd158,8'd164} : s = 37;
	{8'd158,8'd165} : s = 135;
	{8'd158,8'd166} : s = 35;
	{8'd158,8'd167} : s = 120;
	{8'd158,8'd168} : s = 116;
	{8'd158,8'd169} : s = 244;
	{8'd158,8'd170} : s = 28;
	{8'd158,8'd171} : s = 114;
	{8'd158,8'd172} : s = 113;
	{8'd158,8'd173} : s = 242;
	{8'd158,8'd174} : s = 108;
	{8'd158,8'd175} : s = 241;
	{8'd158,8'd176} : s = 236;
	{8'd158,8'd177} : s = 399;
	{8'd158,8'd178} : s = 26;
	{8'd158,8'd179} : s = 106;
	{8'd158,8'd180} : s = 105;
	{8'd158,8'd181} : s = 234;
	{8'd158,8'd182} : s = 102;
	{8'd158,8'd183} : s = 233;
	{8'd158,8'd184} : s = 230;
	{8'd158,8'd185} : s = 380;
	{8'd158,8'd186} : s = 101;
	{8'd158,8'd187} : s = 229;
	{8'd158,8'd188} : s = 227;
	{8'd158,8'd189} : s = 378;
	{8'd158,8'd190} : s = 220;
	{8'd158,8'd191} : s = 377;
	{8'd158,8'd192} : s = 374;
	{8'd158,8'd193} : s = 487;
	{8'd158,8'd194} : s = 25;
	{8'd158,8'd195} : s = 99;
	{8'd158,8'd196} : s = 92;
	{8'd158,8'd197} : s = 218;
	{8'd158,8'd198} : s = 90;
	{8'd158,8'd199} : s = 217;
	{8'd158,8'd200} : s = 214;
	{8'd158,8'd201} : s = 373;
	{8'd158,8'd202} : s = 89;
	{8'd158,8'd203} : s = 213;
	{8'd158,8'd204} : s = 211;
	{8'd158,8'd205} : s = 371;
	{8'd158,8'd206} : s = 206;
	{8'd158,8'd207} : s = 366;
	{8'd158,8'd208} : s = 365;
	{8'd158,8'd209} : s = 478;
	{8'd158,8'd210} : s = 86;
	{8'd158,8'd211} : s = 205;
	{8'd158,8'd212} : s = 203;
	{8'd158,8'd213} : s = 363;
	{8'd158,8'd214} : s = 199;
	{8'd158,8'd215} : s = 359;
	{8'd158,8'd216} : s = 350;
	{8'd158,8'd217} : s = 477;
	{8'd158,8'd218} : s = 188;
	{8'd158,8'd219} : s = 349;
	{8'd158,8'd220} : s = 347;
	{8'd158,8'd221} : s = 475;
	{8'd158,8'd222} : s = 343;
	{8'd158,8'd223} : s = 471;
	{8'd158,8'd224} : s = 463;
	{8'd158,8'd225} : s = 509;
	{8'd158,8'd226} : s = 3;
	{8'd158,8'd227} : s = 22;
	{8'd158,8'd228} : s = 21;
	{8'd158,8'd229} : s = 85;
	{8'd158,8'd230} : s = 19;
	{8'd158,8'd231} : s = 83;
	{8'd158,8'd232} : s = 78;
	{8'd158,8'd233} : s = 186;
	{8'd158,8'd234} : s = 14;
	{8'd158,8'd235} : s = 77;
	{8'd158,8'd236} : s = 75;
	{8'd158,8'd237} : s = 185;
	{8'd158,8'd238} : s = 71;
	{8'd158,8'd239} : s = 182;
	{8'd158,8'd240} : s = 181;
	{8'd158,8'd241} : s = 335;
	{8'd158,8'd242} : s = 13;
	{8'd158,8'd243} : s = 60;
	{8'd158,8'd244} : s = 58;
	{8'd158,8'd245} : s = 179;
	{8'd158,8'd246} : s = 57;
	{8'd158,8'd247} : s = 174;
	{8'd158,8'd248} : s = 173;
	{8'd158,8'd249} : s = 318;
	{8'd158,8'd250} : s = 54;
	{8'd158,8'd251} : s = 171;
	{8'd158,8'd252} : s = 167;
	{8'd158,8'd253} : s = 317;
	{8'd158,8'd254} : s = 158;
	{8'd158,8'd255} : s = 315;
	{8'd159,8'd0} : s = 486;
	{8'd159,8'd1} : s = 24;
	{8'd159,8'd2} : s = 137;
	{8'd159,8'd3} : s = 134;
	{8'd159,8'd4} : s = 291;
	{8'd159,8'd5} : s = 133;
	{8'd159,8'd6} : s = 284;
	{8'd159,8'd7} : s = 282;
	{8'd159,8'd8} : s = 410;
	{8'd159,8'd9} : s = 131;
	{8'd159,8'd10} : s = 281;
	{8'd159,8'd11} : s = 278;
	{8'd159,8'd12} : s = 409;
	{8'd159,8'd13} : s = 277;
	{8'd159,8'd14} : s = 406;
	{8'd159,8'd15} : s = 405;
	{8'd159,8'd16} : s = 485;
	{8'd159,8'd17} : s = 112;
	{8'd159,8'd18} : s = 275;
	{8'd159,8'd19} : s = 270;
	{8'd159,8'd20} : s = 403;
	{8'd159,8'd21} : s = 269;
	{8'd159,8'd22} : s = 398;
	{8'd159,8'd23} : s = 397;
	{8'd159,8'd24} : s = 483;
	{8'd159,8'd25} : s = 267;
	{8'd159,8'd26} : s = 395;
	{8'd159,8'd27} : s = 391;
	{8'd159,8'd28} : s = 476;
	{8'd159,8'd29} : s = 376;
	{8'd159,8'd30} : s = 474;
	{8'd159,8'd31} : s = 473;
	{8'd159,8'd32} : s = 506;
	{8'd159,8'd33} : s = 20;
	{8'd159,8'd34} : s = 104;
	{8'd159,8'd35} : s = 100;
	{8'd159,8'd36} : s = 263;
	{8'd159,8'd37} : s = 98;
	{8'd159,8'd38} : s = 240;
	{8'd159,8'd39} : s = 232;
	{8'd159,8'd40} : s = 372;
	{8'd159,8'd41} : s = 97;
	{8'd159,8'd42} : s = 228;
	{8'd159,8'd43} : s = 226;
	{8'd159,8'd44} : s = 370;
	{8'd159,8'd45} : s = 225;
	{8'd159,8'd46} : s = 369;
	{8'd159,8'd47} : s = 364;
	{8'd159,8'd48} : s = 470;
	{8'd159,8'd49} : s = 88;
	{8'd159,8'd50} : s = 216;
	{8'd159,8'd51} : s = 212;
	{8'd159,8'd52} : s = 362;
	{8'd159,8'd53} : s = 210;
	{8'd159,8'd54} : s = 361;
	{8'd159,8'd55} : s = 358;
	{8'd159,8'd56} : s = 469;
	{8'd159,8'd57} : s = 209;
	{8'd159,8'd58} : s = 357;
	{8'd159,8'd59} : s = 355;
	{8'd159,8'd60} : s = 467;
	{8'd159,8'd61} : s = 348;
	{8'd159,8'd62} : s = 462;
	{8'd159,8'd63} : s = 461;
	{8'd159,8'd64} : s = 505;
	{8'd159,8'd65} : s = 84;
	{8'd159,8'd66} : s = 204;
	{8'd159,8'd67} : s = 202;
	{8'd159,8'd68} : s = 346;
	{8'd159,8'd69} : s = 201;
	{8'd159,8'd70} : s = 345;
	{8'd159,8'd71} : s = 342;
	{8'd159,8'd72} : s = 459;
	{8'd159,8'd73} : s = 198;
	{8'd159,8'd74} : s = 341;
	{8'd159,8'd75} : s = 339;
	{8'd159,8'd76} : s = 455;
	{8'd159,8'd77} : s = 334;
	{8'd159,8'd78} : s = 444;
	{8'd159,8'd79} : s = 442;
	{8'd159,8'd80} : s = 502;
	{8'd159,8'd81} : s = 197;
	{8'd159,8'd82} : s = 333;
	{8'd159,8'd83} : s = 331;
	{8'd159,8'd84} : s = 441;
	{8'd159,8'd85} : s = 327;
	{8'd159,8'd86} : s = 438;
	{8'd159,8'd87} : s = 437;
	{8'd159,8'd88} : s = 501;
	{8'd159,8'd89} : s = 316;
	{8'd159,8'd90} : s = 435;
	{8'd159,8'd91} : s = 430;
	{8'd159,8'd92} : s = 499;
	{8'd159,8'd93} : s = 429;
	{8'd159,8'd94} : s = 494;
	{8'd159,8'd95} : s = 493;
	{8'd159,8'd96} : s = 510;
	{8'd159,8'd97} : s = 1;
	{8'd159,8'd98} : s = 18;
	{8'd159,8'd99} : s = 17;
	{8'd159,8'd100} : s = 82;
	{8'd159,8'd101} : s = 12;
	{8'd159,8'd102} : s = 81;
	{8'd159,8'd103} : s = 76;
	{8'd159,8'd104} : s = 195;
	{8'd159,8'd105} : s = 10;
	{8'd159,8'd106} : s = 74;
	{8'd159,8'd107} : s = 73;
	{8'd159,8'd108} : s = 184;
	{8'd159,8'd109} : s = 70;
	{8'd159,8'd110} : s = 180;
	{8'd159,8'd111} : s = 178;
	{8'd159,8'd112} : s = 314;
	{8'd159,8'd113} : s = 9;
	{8'd159,8'd114} : s = 69;
	{8'd159,8'd115} : s = 67;
	{8'd159,8'd116} : s = 177;
	{8'd159,8'd117} : s = 56;
	{8'd159,8'd118} : s = 172;
	{8'd159,8'd119} : s = 170;
	{8'd159,8'd120} : s = 313;
	{8'd159,8'd121} : s = 52;
	{8'd159,8'd122} : s = 169;
	{8'd159,8'd123} : s = 166;
	{8'd159,8'd124} : s = 310;
	{8'd159,8'd125} : s = 165;
	{8'd159,8'd126} : s = 309;
	{8'd159,8'd127} : s = 307;
	{8'd159,8'd128} : s = 427;
	{8'd159,8'd129} : s = 6;
	{8'd159,8'd130} : s = 50;
	{8'd159,8'd131} : s = 49;
	{8'd159,8'd132} : s = 163;
	{8'd159,8'd133} : s = 44;
	{8'd159,8'd134} : s = 156;
	{8'd159,8'd135} : s = 154;
	{8'd159,8'd136} : s = 302;
	{8'd159,8'd137} : s = 42;
	{8'd159,8'd138} : s = 153;
	{8'd159,8'd139} : s = 150;
	{8'd159,8'd140} : s = 301;
	{8'd159,8'd141} : s = 149;
	{8'd159,8'd142} : s = 299;
	{8'd159,8'd143} : s = 295;
	{8'd159,8'd144} : s = 423;
	{8'd159,8'd145} : s = 41;
	{8'd159,8'd146} : s = 147;
	{8'd159,8'd147} : s = 142;
	{8'd159,8'd148} : s = 286;
	{8'd159,8'd149} : s = 141;
	{8'd159,8'd150} : s = 285;
	{8'd159,8'd151} : s = 283;
	{8'd159,8'd152} : s = 414;
	{8'd159,8'd153} : s = 139;
	{8'd159,8'd154} : s = 279;
	{8'd159,8'd155} : s = 271;
	{8'd159,8'd156} : s = 413;
	{8'd159,8'd157} : s = 248;
	{8'd159,8'd158} : s = 411;
	{8'd159,8'd159} : s = 407;
	{8'd159,8'd160} : s = 491;
	{8'd159,8'd161} : s = 5;
	{8'd159,8'd162} : s = 38;
	{8'd159,8'd163} : s = 37;
	{8'd159,8'd164} : s = 135;
	{8'd159,8'd165} : s = 35;
	{8'd159,8'd166} : s = 120;
	{8'd159,8'd167} : s = 116;
	{8'd159,8'd168} : s = 244;
	{8'd159,8'd169} : s = 28;
	{8'd159,8'd170} : s = 114;
	{8'd159,8'd171} : s = 113;
	{8'd159,8'd172} : s = 242;
	{8'd159,8'd173} : s = 108;
	{8'd159,8'd174} : s = 241;
	{8'd159,8'd175} : s = 236;
	{8'd159,8'd176} : s = 399;
	{8'd159,8'd177} : s = 26;
	{8'd159,8'd178} : s = 106;
	{8'd159,8'd179} : s = 105;
	{8'd159,8'd180} : s = 234;
	{8'd159,8'd181} : s = 102;
	{8'd159,8'd182} : s = 233;
	{8'd159,8'd183} : s = 230;
	{8'd159,8'd184} : s = 380;
	{8'd159,8'd185} : s = 101;
	{8'd159,8'd186} : s = 229;
	{8'd159,8'd187} : s = 227;
	{8'd159,8'd188} : s = 378;
	{8'd159,8'd189} : s = 220;
	{8'd159,8'd190} : s = 377;
	{8'd159,8'd191} : s = 374;
	{8'd159,8'd192} : s = 487;
	{8'd159,8'd193} : s = 25;
	{8'd159,8'd194} : s = 99;
	{8'd159,8'd195} : s = 92;
	{8'd159,8'd196} : s = 218;
	{8'd159,8'd197} : s = 90;
	{8'd159,8'd198} : s = 217;
	{8'd159,8'd199} : s = 214;
	{8'd159,8'd200} : s = 373;
	{8'd159,8'd201} : s = 89;
	{8'd159,8'd202} : s = 213;
	{8'd159,8'd203} : s = 211;
	{8'd159,8'd204} : s = 371;
	{8'd159,8'd205} : s = 206;
	{8'd159,8'd206} : s = 366;
	{8'd159,8'd207} : s = 365;
	{8'd159,8'd208} : s = 478;
	{8'd159,8'd209} : s = 86;
	{8'd159,8'd210} : s = 205;
	{8'd159,8'd211} : s = 203;
	{8'd159,8'd212} : s = 363;
	{8'd159,8'd213} : s = 199;
	{8'd159,8'd214} : s = 359;
	{8'd159,8'd215} : s = 350;
	{8'd159,8'd216} : s = 477;
	{8'd159,8'd217} : s = 188;
	{8'd159,8'd218} : s = 349;
	{8'd159,8'd219} : s = 347;
	{8'd159,8'd220} : s = 475;
	{8'd159,8'd221} : s = 343;
	{8'd159,8'd222} : s = 471;
	{8'd159,8'd223} : s = 463;
	{8'd159,8'd224} : s = 509;
	{8'd159,8'd225} : s = 3;
	{8'd159,8'd226} : s = 22;
	{8'd159,8'd227} : s = 21;
	{8'd159,8'd228} : s = 85;
	{8'd159,8'd229} : s = 19;
	{8'd159,8'd230} : s = 83;
	{8'd159,8'd231} : s = 78;
	{8'd159,8'd232} : s = 186;
	{8'd159,8'd233} : s = 14;
	{8'd159,8'd234} : s = 77;
	{8'd159,8'd235} : s = 75;
	{8'd159,8'd236} : s = 185;
	{8'd159,8'd237} : s = 71;
	{8'd159,8'd238} : s = 182;
	{8'd159,8'd239} : s = 181;
	{8'd159,8'd240} : s = 335;
	{8'd159,8'd241} : s = 13;
	{8'd159,8'd242} : s = 60;
	{8'd159,8'd243} : s = 58;
	{8'd159,8'd244} : s = 179;
	{8'd159,8'd245} : s = 57;
	{8'd159,8'd246} : s = 174;
	{8'd159,8'd247} : s = 173;
	{8'd159,8'd248} : s = 318;
	{8'd159,8'd249} : s = 54;
	{8'd159,8'd250} : s = 171;
	{8'd159,8'd251} : s = 167;
	{8'd159,8'd252} : s = 317;
	{8'd159,8'd253} : s = 158;
	{8'd159,8'd254} : s = 315;
	{8'd159,8'd255} : s = 311;
	{8'd160,8'd0} : s = 24;
	{8'd160,8'd1} : s = 137;
	{8'd160,8'd2} : s = 134;
	{8'd160,8'd3} : s = 291;
	{8'd160,8'd4} : s = 133;
	{8'd160,8'd5} : s = 284;
	{8'd160,8'd6} : s = 282;
	{8'd160,8'd7} : s = 410;
	{8'd160,8'd8} : s = 131;
	{8'd160,8'd9} : s = 281;
	{8'd160,8'd10} : s = 278;
	{8'd160,8'd11} : s = 409;
	{8'd160,8'd12} : s = 277;
	{8'd160,8'd13} : s = 406;
	{8'd160,8'd14} : s = 405;
	{8'd160,8'd15} : s = 485;
	{8'd160,8'd16} : s = 112;
	{8'd160,8'd17} : s = 275;
	{8'd160,8'd18} : s = 270;
	{8'd160,8'd19} : s = 403;
	{8'd160,8'd20} : s = 269;
	{8'd160,8'd21} : s = 398;
	{8'd160,8'd22} : s = 397;
	{8'd160,8'd23} : s = 483;
	{8'd160,8'd24} : s = 267;
	{8'd160,8'd25} : s = 395;
	{8'd160,8'd26} : s = 391;
	{8'd160,8'd27} : s = 476;
	{8'd160,8'd28} : s = 376;
	{8'd160,8'd29} : s = 474;
	{8'd160,8'd30} : s = 473;
	{8'd160,8'd31} : s = 506;
	{8'd160,8'd32} : s = 20;
	{8'd160,8'd33} : s = 104;
	{8'd160,8'd34} : s = 100;
	{8'd160,8'd35} : s = 263;
	{8'd160,8'd36} : s = 98;
	{8'd160,8'd37} : s = 240;
	{8'd160,8'd38} : s = 232;
	{8'd160,8'd39} : s = 372;
	{8'd160,8'd40} : s = 97;
	{8'd160,8'd41} : s = 228;
	{8'd160,8'd42} : s = 226;
	{8'd160,8'd43} : s = 370;
	{8'd160,8'd44} : s = 225;
	{8'd160,8'd45} : s = 369;
	{8'd160,8'd46} : s = 364;
	{8'd160,8'd47} : s = 470;
	{8'd160,8'd48} : s = 88;
	{8'd160,8'd49} : s = 216;
	{8'd160,8'd50} : s = 212;
	{8'd160,8'd51} : s = 362;
	{8'd160,8'd52} : s = 210;
	{8'd160,8'd53} : s = 361;
	{8'd160,8'd54} : s = 358;
	{8'd160,8'd55} : s = 469;
	{8'd160,8'd56} : s = 209;
	{8'd160,8'd57} : s = 357;
	{8'd160,8'd58} : s = 355;
	{8'd160,8'd59} : s = 467;
	{8'd160,8'd60} : s = 348;
	{8'd160,8'd61} : s = 462;
	{8'd160,8'd62} : s = 461;
	{8'd160,8'd63} : s = 505;
	{8'd160,8'd64} : s = 84;
	{8'd160,8'd65} : s = 204;
	{8'd160,8'd66} : s = 202;
	{8'd160,8'd67} : s = 346;
	{8'd160,8'd68} : s = 201;
	{8'd160,8'd69} : s = 345;
	{8'd160,8'd70} : s = 342;
	{8'd160,8'd71} : s = 459;
	{8'd160,8'd72} : s = 198;
	{8'd160,8'd73} : s = 341;
	{8'd160,8'd74} : s = 339;
	{8'd160,8'd75} : s = 455;
	{8'd160,8'd76} : s = 334;
	{8'd160,8'd77} : s = 444;
	{8'd160,8'd78} : s = 442;
	{8'd160,8'd79} : s = 502;
	{8'd160,8'd80} : s = 197;
	{8'd160,8'd81} : s = 333;
	{8'd160,8'd82} : s = 331;
	{8'd160,8'd83} : s = 441;
	{8'd160,8'd84} : s = 327;
	{8'd160,8'd85} : s = 438;
	{8'd160,8'd86} : s = 437;
	{8'd160,8'd87} : s = 501;
	{8'd160,8'd88} : s = 316;
	{8'd160,8'd89} : s = 435;
	{8'd160,8'd90} : s = 430;
	{8'd160,8'd91} : s = 499;
	{8'd160,8'd92} : s = 429;
	{8'd160,8'd93} : s = 494;
	{8'd160,8'd94} : s = 493;
	{8'd160,8'd95} : s = 510;
	{8'd160,8'd96} : s = 1;
	{8'd160,8'd97} : s = 18;
	{8'd160,8'd98} : s = 17;
	{8'd160,8'd99} : s = 82;
	{8'd160,8'd100} : s = 12;
	{8'd160,8'd101} : s = 81;
	{8'd160,8'd102} : s = 76;
	{8'd160,8'd103} : s = 195;
	{8'd160,8'd104} : s = 10;
	{8'd160,8'd105} : s = 74;
	{8'd160,8'd106} : s = 73;
	{8'd160,8'd107} : s = 184;
	{8'd160,8'd108} : s = 70;
	{8'd160,8'd109} : s = 180;
	{8'd160,8'd110} : s = 178;
	{8'd160,8'd111} : s = 314;
	{8'd160,8'd112} : s = 9;
	{8'd160,8'd113} : s = 69;
	{8'd160,8'd114} : s = 67;
	{8'd160,8'd115} : s = 177;
	{8'd160,8'd116} : s = 56;
	{8'd160,8'd117} : s = 172;
	{8'd160,8'd118} : s = 170;
	{8'd160,8'd119} : s = 313;
	{8'd160,8'd120} : s = 52;
	{8'd160,8'd121} : s = 169;
	{8'd160,8'd122} : s = 166;
	{8'd160,8'd123} : s = 310;
	{8'd160,8'd124} : s = 165;
	{8'd160,8'd125} : s = 309;
	{8'd160,8'd126} : s = 307;
	{8'd160,8'd127} : s = 427;
	{8'd160,8'd128} : s = 6;
	{8'd160,8'd129} : s = 50;
	{8'd160,8'd130} : s = 49;
	{8'd160,8'd131} : s = 163;
	{8'd160,8'd132} : s = 44;
	{8'd160,8'd133} : s = 156;
	{8'd160,8'd134} : s = 154;
	{8'd160,8'd135} : s = 302;
	{8'd160,8'd136} : s = 42;
	{8'd160,8'd137} : s = 153;
	{8'd160,8'd138} : s = 150;
	{8'd160,8'd139} : s = 301;
	{8'd160,8'd140} : s = 149;
	{8'd160,8'd141} : s = 299;
	{8'd160,8'd142} : s = 295;
	{8'd160,8'd143} : s = 423;
	{8'd160,8'd144} : s = 41;
	{8'd160,8'd145} : s = 147;
	{8'd160,8'd146} : s = 142;
	{8'd160,8'd147} : s = 286;
	{8'd160,8'd148} : s = 141;
	{8'd160,8'd149} : s = 285;
	{8'd160,8'd150} : s = 283;
	{8'd160,8'd151} : s = 414;
	{8'd160,8'd152} : s = 139;
	{8'd160,8'd153} : s = 279;
	{8'd160,8'd154} : s = 271;
	{8'd160,8'd155} : s = 413;
	{8'd160,8'd156} : s = 248;
	{8'd160,8'd157} : s = 411;
	{8'd160,8'd158} : s = 407;
	{8'd160,8'd159} : s = 491;
	{8'd160,8'd160} : s = 5;
	{8'd160,8'd161} : s = 38;
	{8'd160,8'd162} : s = 37;
	{8'd160,8'd163} : s = 135;
	{8'd160,8'd164} : s = 35;
	{8'd160,8'd165} : s = 120;
	{8'd160,8'd166} : s = 116;
	{8'd160,8'd167} : s = 244;
	{8'd160,8'd168} : s = 28;
	{8'd160,8'd169} : s = 114;
	{8'd160,8'd170} : s = 113;
	{8'd160,8'd171} : s = 242;
	{8'd160,8'd172} : s = 108;
	{8'd160,8'd173} : s = 241;
	{8'd160,8'd174} : s = 236;
	{8'd160,8'd175} : s = 399;
	{8'd160,8'd176} : s = 26;
	{8'd160,8'd177} : s = 106;
	{8'd160,8'd178} : s = 105;
	{8'd160,8'd179} : s = 234;
	{8'd160,8'd180} : s = 102;
	{8'd160,8'd181} : s = 233;
	{8'd160,8'd182} : s = 230;
	{8'd160,8'd183} : s = 380;
	{8'd160,8'd184} : s = 101;
	{8'd160,8'd185} : s = 229;
	{8'd160,8'd186} : s = 227;
	{8'd160,8'd187} : s = 378;
	{8'd160,8'd188} : s = 220;
	{8'd160,8'd189} : s = 377;
	{8'd160,8'd190} : s = 374;
	{8'd160,8'd191} : s = 487;
	{8'd160,8'd192} : s = 25;
	{8'd160,8'd193} : s = 99;
	{8'd160,8'd194} : s = 92;
	{8'd160,8'd195} : s = 218;
	{8'd160,8'd196} : s = 90;
	{8'd160,8'd197} : s = 217;
	{8'd160,8'd198} : s = 214;
	{8'd160,8'd199} : s = 373;
	{8'd160,8'd200} : s = 89;
	{8'd160,8'd201} : s = 213;
	{8'd160,8'd202} : s = 211;
	{8'd160,8'd203} : s = 371;
	{8'd160,8'd204} : s = 206;
	{8'd160,8'd205} : s = 366;
	{8'd160,8'd206} : s = 365;
	{8'd160,8'd207} : s = 478;
	{8'd160,8'd208} : s = 86;
	{8'd160,8'd209} : s = 205;
	{8'd160,8'd210} : s = 203;
	{8'd160,8'd211} : s = 363;
	{8'd160,8'd212} : s = 199;
	{8'd160,8'd213} : s = 359;
	{8'd160,8'd214} : s = 350;
	{8'd160,8'd215} : s = 477;
	{8'd160,8'd216} : s = 188;
	{8'd160,8'd217} : s = 349;
	{8'd160,8'd218} : s = 347;
	{8'd160,8'd219} : s = 475;
	{8'd160,8'd220} : s = 343;
	{8'd160,8'd221} : s = 471;
	{8'd160,8'd222} : s = 463;
	{8'd160,8'd223} : s = 509;
	{8'd160,8'd224} : s = 3;
	{8'd160,8'd225} : s = 22;
	{8'd160,8'd226} : s = 21;
	{8'd160,8'd227} : s = 85;
	{8'd160,8'd228} : s = 19;
	{8'd160,8'd229} : s = 83;
	{8'd160,8'd230} : s = 78;
	{8'd160,8'd231} : s = 186;
	{8'd160,8'd232} : s = 14;
	{8'd160,8'd233} : s = 77;
	{8'd160,8'd234} : s = 75;
	{8'd160,8'd235} : s = 185;
	{8'd160,8'd236} : s = 71;
	{8'd160,8'd237} : s = 182;
	{8'd160,8'd238} : s = 181;
	{8'd160,8'd239} : s = 335;
	{8'd160,8'd240} : s = 13;
	{8'd160,8'd241} : s = 60;
	{8'd160,8'd242} : s = 58;
	{8'd160,8'd243} : s = 179;
	{8'd160,8'd244} : s = 57;
	{8'd160,8'd245} : s = 174;
	{8'd160,8'd246} : s = 173;
	{8'd160,8'd247} : s = 318;
	{8'd160,8'd248} : s = 54;
	{8'd160,8'd249} : s = 171;
	{8'd160,8'd250} : s = 167;
	{8'd160,8'd251} : s = 317;
	{8'd160,8'd252} : s = 158;
	{8'd160,8'd253} : s = 315;
	{8'd160,8'd254} : s = 311;
	{8'd160,8'd255} : s = 446;
	{8'd161,8'd0} : s = 137;
	{8'd161,8'd1} : s = 134;
	{8'd161,8'd2} : s = 291;
	{8'd161,8'd3} : s = 133;
	{8'd161,8'd4} : s = 284;
	{8'd161,8'd5} : s = 282;
	{8'd161,8'd6} : s = 410;
	{8'd161,8'd7} : s = 131;
	{8'd161,8'd8} : s = 281;
	{8'd161,8'd9} : s = 278;
	{8'd161,8'd10} : s = 409;
	{8'd161,8'd11} : s = 277;
	{8'd161,8'd12} : s = 406;
	{8'd161,8'd13} : s = 405;
	{8'd161,8'd14} : s = 485;
	{8'd161,8'd15} : s = 112;
	{8'd161,8'd16} : s = 275;
	{8'd161,8'd17} : s = 270;
	{8'd161,8'd18} : s = 403;
	{8'd161,8'd19} : s = 269;
	{8'd161,8'd20} : s = 398;
	{8'd161,8'd21} : s = 397;
	{8'd161,8'd22} : s = 483;
	{8'd161,8'd23} : s = 267;
	{8'd161,8'd24} : s = 395;
	{8'd161,8'd25} : s = 391;
	{8'd161,8'd26} : s = 476;
	{8'd161,8'd27} : s = 376;
	{8'd161,8'd28} : s = 474;
	{8'd161,8'd29} : s = 473;
	{8'd161,8'd30} : s = 506;
	{8'd161,8'd31} : s = 20;
	{8'd161,8'd32} : s = 104;
	{8'd161,8'd33} : s = 100;
	{8'd161,8'd34} : s = 263;
	{8'd161,8'd35} : s = 98;
	{8'd161,8'd36} : s = 240;
	{8'd161,8'd37} : s = 232;
	{8'd161,8'd38} : s = 372;
	{8'd161,8'd39} : s = 97;
	{8'd161,8'd40} : s = 228;
	{8'd161,8'd41} : s = 226;
	{8'd161,8'd42} : s = 370;
	{8'd161,8'd43} : s = 225;
	{8'd161,8'd44} : s = 369;
	{8'd161,8'd45} : s = 364;
	{8'd161,8'd46} : s = 470;
	{8'd161,8'd47} : s = 88;
	{8'd161,8'd48} : s = 216;
	{8'd161,8'd49} : s = 212;
	{8'd161,8'd50} : s = 362;
	{8'd161,8'd51} : s = 210;
	{8'd161,8'd52} : s = 361;
	{8'd161,8'd53} : s = 358;
	{8'd161,8'd54} : s = 469;
	{8'd161,8'd55} : s = 209;
	{8'd161,8'd56} : s = 357;
	{8'd161,8'd57} : s = 355;
	{8'd161,8'd58} : s = 467;
	{8'd161,8'd59} : s = 348;
	{8'd161,8'd60} : s = 462;
	{8'd161,8'd61} : s = 461;
	{8'd161,8'd62} : s = 505;
	{8'd161,8'd63} : s = 84;
	{8'd161,8'd64} : s = 204;
	{8'd161,8'd65} : s = 202;
	{8'd161,8'd66} : s = 346;
	{8'd161,8'd67} : s = 201;
	{8'd161,8'd68} : s = 345;
	{8'd161,8'd69} : s = 342;
	{8'd161,8'd70} : s = 459;
	{8'd161,8'd71} : s = 198;
	{8'd161,8'd72} : s = 341;
	{8'd161,8'd73} : s = 339;
	{8'd161,8'd74} : s = 455;
	{8'd161,8'd75} : s = 334;
	{8'd161,8'd76} : s = 444;
	{8'd161,8'd77} : s = 442;
	{8'd161,8'd78} : s = 502;
	{8'd161,8'd79} : s = 197;
	{8'd161,8'd80} : s = 333;
	{8'd161,8'd81} : s = 331;
	{8'd161,8'd82} : s = 441;
	{8'd161,8'd83} : s = 327;
	{8'd161,8'd84} : s = 438;
	{8'd161,8'd85} : s = 437;
	{8'd161,8'd86} : s = 501;
	{8'd161,8'd87} : s = 316;
	{8'd161,8'd88} : s = 435;
	{8'd161,8'd89} : s = 430;
	{8'd161,8'd90} : s = 499;
	{8'd161,8'd91} : s = 429;
	{8'd161,8'd92} : s = 494;
	{8'd161,8'd93} : s = 493;
	{8'd161,8'd94} : s = 510;
	{8'd161,8'd95} : s = 1;
	{8'd161,8'd96} : s = 18;
	{8'd161,8'd97} : s = 17;
	{8'd161,8'd98} : s = 82;
	{8'd161,8'd99} : s = 12;
	{8'd161,8'd100} : s = 81;
	{8'd161,8'd101} : s = 76;
	{8'd161,8'd102} : s = 195;
	{8'd161,8'd103} : s = 10;
	{8'd161,8'd104} : s = 74;
	{8'd161,8'd105} : s = 73;
	{8'd161,8'd106} : s = 184;
	{8'd161,8'd107} : s = 70;
	{8'd161,8'd108} : s = 180;
	{8'd161,8'd109} : s = 178;
	{8'd161,8'd110} : s = 314;
	{8'd161,8'd111} : s = 9;
	{8'd161,8'd112} : s = 69;
	{8'd161,8'd113} : s = 67;
	{8'd161,8'd114} : s = 177;
	{8'd161,8'd115} : s = 56;
	{8'd161,8'd116} : s = 172;
	{8'd161,8'd117} : s = 170;
	{8'd161,8'd118} : s = 313;
	{8'd161,8'd119} : s = 52;
	{8'd161,8'd120} : s = 169;
	{8'd161,8'd121} : s = 166;
	{8'd161,8'd122} : s = 310;
	{8'd161,8'd123} : s = 165;
	{8'd161,8'd124} : s = 309;
	{8'd161,8'd125} : s = 307;
	{8'd161,8'd126} : s = 427;
	{8'd161,8'd127} : s = 6;
	{8'd161,8'd128} : s = 50;
	{8'd161,8'd129} : s = 49;
	{8'd161,8'd130} : s = 163;
	{8'd161,8'd131} : s = 44;
	{8'd161,8'd132} : s = 156;
	{8'd161,8'd133} : s = 154;
	{8'd161,8'd134} : s = 302;
	{8'd161,8'd135} : s = 42;
	{8'd161,8'd136} : s = 153;
	{8'd161,8'd137} : s = 150;
	{8'd161,8'd138} : s = 301;
	{8'd161,8'd139} : s = 149;
	{8'd161,8'd140} : s = 299;
	{8'd161,8'd141} : s = 295;
	{8'd161,8'd142} : s = 423;
	{8'd161,8'd143} : s = 41;
	{8'd161,8'd144} : s = 147;
	{8'd161,8'd145} : s = 142;
	{8'd161,8'd146} : s = 286;
	{8'd161,8'd147} : s = 141;
	{8'd161,8'd148} : s = 285;
	{8'd161,8'd149} : s = 283;
	{8'd161,8'd150} : s = 414;
	{8'd161,8'd151} : s = 139;
	{8'd161,8'd152} : s = 279;
	{8'd161,8'd153} : s = 271;
	{8'd161,8'd154} : s = 413;
	{8'd161,8'd155} : s = 248;
	{8'd161,8'd156} : s = 411;
	{8'd161,8'd157} : s = 407;
	{8'd161,8'd158} : s = 491;
	{8'd161,8'd159} : s = 5;
	{8'd161,8'd160} : s = 38;
	{8'd161,8'd161} : s = 37;
	{8'd161,8'd162} : s = 135;
	{8'd161,8'd163} : s = 35;
	{8'd161,8'd164} : s = 120;
	{8'd161,8'd165} : s = 116;
	{8'd161,8'd166} : s = 244;
	{8'd161,8'd167} : s = 28;
	{8'd161,8'd168} : s = 114;
	{8'd161,8'd169} : s = 113;
	{8'd161,8'd170} : s = 242;
	{8'd161,8'd171} : s = 108;
	{8'd161,8'd172} : s = 241;
	{8'd161,8'd173} : s = 236;
	{8'd161,8'd174} : s = 399;
	{8'd161,8'd175} : s = 26;
	{8'd161,8'd176} : s = 106;
	{8'd161,8'd177} : s = 105;
	{8'd161,8'd178} : s = 234;
	{8'd161,8'd179} : s = 102;
	{8'd161,8'd180} : s = 233;
	{8'd161,8'd181} : s = 230;
	{8'd161,8'd182} : s = 380;
	{8'd161,8'd183} : s = 101;
	{8'd161,8'd184} : s = 229;
	{8'd161,8'd185} : s = 227;
	{8'd161,8'd186} : s = 378;
	{8'd161,8'd187} : s = 220;
	{8'd161,8'd188} : s = 377;
	{8'd161,8'd189} : s = 374;
	{8'd161,8'd190} : s = 487;
	{8'd161,8'd191} : s = 25;
	{8'd161,8'd192} : s = 99;
	{8'd161,8'd193} : s = 92;
	{8'd161,8'd194} : s = 218;
	{8'd161,8'd195} : s = 90;
	{8'd161,8'd196} : s = 217;
	{8'd161,8'd197} : s = 214;
	{8'd161,8'd198} : s = 373;
	{8'd161,8'd199} : s = 89;
	{8'd161,8'd200} : s = 213;
	{8'd161,8'd201} : s = 211;
	{8'd161,8'd202} : s = 371;
	{8'd161,8'd203} : s = 206;
	{8'd161,8'd204} : s = 366;
	{8'd161,8'd205} : s = 365;
	{8'd161,8'd206} : s = 478;
	{8'd161,8'd207} : s = 86;
	{8'd161,8'd208} : s = 205;
	{8'd161,8'd209} : s = 203;
	{8'd161,8'd210} : s = 363;
	{8'd161,8'd211} : s = 199;
	{8'd161,8'd212} : s = 359;
	{8'd161,8'd213} : s = 350;
	{8'd161,8'd214} : s = 477;
	{8'd161,8'd215} : s = 188;
	{8'd161,8'd216} : s = 349;
	{8'd161,8'd217} : s = 347;
	{8'd161,8'd218} : s = 475;
	{8'd161,8'd219} : s = 343;
	{8'd161,8'd220} : s = 471;
	{8'd161,8'd221} : s = 463;
	{8'd161,8'd222} : s = 509;
	{8'd161,8'd223} : s = 3;
	{8'd161,8'd224} : s = 22;
	{8'd161,8'd225} : s = 21;
	{8'd161,8'd226} : s = 85;
	{8'd161,8'd227} : s = 19;
	{8'd161,8'd228} : s = 83;
	{8'd161,8'd229} : s = 78;
	{8'd161,8'd230} : s = 186;
	{8'd161,8'd231} : s = 14;
	{8'd161,8'd232} : s = 77;
	{8'd161,8'd233} : s = 75;
	{8'd161,8'd234} : s = 185;
	{8'd161,8'd235} : s = 71;
	{8'd161,8'd236} : s = 182;
	{8'd161,8'd237} : s = 181;
	{8'd161,8'd238} : s = 335;
	{8'd161,8'd239} : s = 13;
	{8'd161,8'd240} : s = 60;
	{8'd161,8'd241} : s = 58;
	{8'd161,8'd242} : s = 179;
	{8'd161,8'd243} : s = 57;
	{8'd161,8'd244} : s = 174;
	{8'd161,8'd245} : s = 173;
	{8'd161,8'd246} : s = 318;
	{8'd161,8'd247} : s = 54;
	{8'd161,8'd248} : s = 171;
	{8'd161,8'd249} : s = 167;
	{8'd161,8'd250} : s = 317;
	{8'd161,8'd251} : s = 158;
	{8'd161,8'd252} : s = 315;
	{8'd161,8'd253} : s = 311;
	{8'd161,8'd254} : s = 446;
	{8'd161,8'd255} : s = 11;
	{8'd162,8'd0} : s = 134;
	{8'd162,8'd1} : s = 291;
	{8'd162,8'd2} : s = 133;
	{8'd162,8'd3} : s = 284;
	{8'd162,8'd4} : s = 282;
	{8'd162,8'd5} : s = 410;
	{8'd162,8'd6} : s = 131;
	{8'd162,8'd7} : s = 281;
	{8'd162,8'd8} : s = 278;
	{8'd162,8'd9} : s = 409;
	{8'd162,8'd10} : s = 277;
	{8'd162,8'd11} : s = 406;
	{8'd162,8'd12} : s = 405;
	{8'd162,8'd13} : s = 485;
	{8'd162,8'd14} : s = 112;
	{8'd162,8'd15} : s = 275;
	{8'd162,8'd16} : s = 270;
	{8'd162,8'd17} : s = 403;
	{8'd162,8'd18} : s = 269;
	{8'd162,8'd19} : s = 398;
	{8'd162,8'd20} : s = 397;
	{8'd162,8'd21} : s = 483;
	{8'd162,8'd22} : s = 267;
	{8'd162,8'd23} : s = 395;
	{8'd162,8'd24} : s = 391;
	{8'd162,8'd25} : s = 476;
	{8'd162,8'd26} : s = 376;
	{8'd162,8'd27} : s = 474;
	{8'd162,8'd28} : s = 473;
	{8'd162,8'd29} : s = 506;
	{8'd162,8'd30} : s = 20;
	{8'd162,8'd31} : s = 104;
	{8'd162,8'd32} : s = 100;
	{8'd162,8'd33} : s = 263;
	{8'd162,8'd34} : s = 98;
	{8'd162,8'd35} : s = 240;
	{8'd162,8'd36} : s = 232;
	{8'd162,8'd37} : s = 372;
	{8'd162,8'd38} : s = 97;
	{8'd162,8'd39} : s = 228;
	{8'd162,8'd40} : s = 226;
	{8'd162,8'd41} : s = 370;
	{8'd162,8'd42} : s = 225;
	{8'd162,8'd43} : s = 369;
	{8'd162,8'd44} : s = 364;
	{8'd162,8'd45} : s = 470;
	{8'd162,8'd46} : s = 88;
	{8'd162,8'd47} : s = 216;
	{8'd162,8'd48} : s = 212;
	{8'd162,8'd49} : s = 362;
	{8'd162,8'd50} : s = 210;
	{8'd162,8'd51} : s = 361;
	{8'd162,8'd52} : s = 358;
	{8'd162,8'd53} : s = 469;
	{8'd162,8'd54} : s = 209;
	{8'd162,8'd55} : s = 357;
	{8'd162,8'd56} : s = 355;
	{8'd162,8'd57} : s = 467;
	{8'd162,8'd58} : s = 348;
	{8'd162,8'd59} : s = 462;
	{8'd162,8'd60} : s = 461;
	{8'd162,8'd61} : s = 505;
	{8'd162,8'd62} : s = 84;
	{8'd162,8'd63} : s = 204;
	{8'd162,8'd64} : s = 202;
	{8'd162,8'd65} : s = 346;
	{8'd162,8'd66} : s = 201;
	{8'd162,8'd67} : s = 345;
	{8'd162,8'd68} : s = 342;
	{8'd162,8'd69} : s = 459;
	{8'd162,8'd70} : s = 198;
	{8'd162,8'd71} : s = 341;
	{8'd162,8'd72} : s = 339;
	{8'd162,8'd73} : s = 455;
	{8'd162,8'd74} : s = 334;
	{8'd162,8'd75} : s = 444;
	{8'd162,8'd76} : s = 442;
	{8'd162,8'd77} : s = 502;
	{8'd162,8'd78} : s = 197;
	{8'd162,8'd79} : s = 333;
	{8'd162,8'd80} : s = 331;
	{8'd162,8'd81} : s = 441;
	{8'd162,8'd82} : s = 327;
	{8'd162,8'd83} : s = 438;
	{8'd162,8'd84} : s = 437;
	{8'd162,8'd85} : s = 501;
	{8'd162,8'd86} : s = 316;
	{8'd162,8'd87} : s = 435;
	{8'd162,8'd88} : s = 430;
	{8'd162,8'd89} : s = 499;
	{8'd162,8'd90} : s = 429;
	{8'd162,8'd91} : s = 494;
	{8'd162,8'd92} : s = 493;
	{8'd162,8'd93} : s = 510;
	{8'd162,8'd94} : s = 1;
	{8'd162,8'd95} : s = 18;
	{8'd162,8'd96} : s = 17;
	{8'd162,8'd97} : s = 82;
	{8'd162,8'd98} : s = 12;
	{8'd162,8'd99} : s = 81;
	{8'd162,8'd100} : s = 76;
	{8'd162,8'd101} : s = 195;
	{8'd162,8'd102} : s = 10;
	{8'd162,8'd103} : s = 74;
	{8'd162,8'd104} : s = 73;
	{8'd162,8'd105} : s = 184;
	{8'd162,8'd106} : s = 70;
	{8'd162,8'd107} : s = 180;
	{8'd162,8'd108} : s = 178;
	{8'd162,8'd109} : s = 314;
	{8'd162,8'd110} : s = 9;
	{8'd162,8'd111} : s = 69;
	{8'd162,8'd112} : s = 67;
	{8'd162,8'd113} : s = 177;
	{8'd162,8'd114} : s = 56;
	{8'd162,8'd115} : s = 172;
	{8'd162,8'd116} : s = 170;
	{8'd162,8'd117} : s = 313;
	{8'd162,8'd118} : s = 52;
	{8'd162,8'd119} : s = 169;
	{8'd162,8'd120} : s = 166;
	{8'd162,8'd121} : s = 310;
	{8'd162,8'd122} : s = 165;
	{8'd162,8'd123} : s = 309;
	{8'd162,8'd124} : s = 307;
	{8'd162,8'd125} : s = 427;
	{8'd162,8'd126} : s = 6;
	{8'd162,8'd127} : s = 50;
	{8'd162,8'd128} : s = 49;
	{8'd162,8'd129} : s = 163;
	{8'd162,8'd130} : s = 44;
	{8'd162,8'd131} : s = 156;
	{8'd162,8'd132} : s = 154;
	{8'd162,8'd133} : s = 302;
	{8'd162,8'd134} : s = 42;
	{8'd162,8'd135} : s = 153;
	{8'd162,8'd136} : s = 150;
	{8'd162,8'd137} : s = 301;
	{8'd162,8'd138} : s = 149;
	{8'd162,8'd139} : s = 299;
	{8'd162,8'd140} : s = 295;
	{8'd162,8'd141} : s = 423;
	{8'd162,8'd142} : s = 41;
	{8'd162,8'd143} : s = 147;
	{8'd162,8'd144} : s = 142;
	{8'd162,8'd145} : s = 286;
	{8'd162,8'd146} : s = 141;
	{8'd162,8'd147} : s = 285;
	{8'd162,8'd148} : s = 283;
	{8'd162,8'd149} : s = 414;
	{8'd162,8'd150} : s = 139;
	{8'd162,8'd151} : s = 279;
	{8'd162,8'd152} : s = 271;
	{8'd162,8'd153} : s = 413;
	{8'd162,8'd154} : s = 248;
	{8'd162,8'd155} : s = 411;
	{8'd162,8'd156} : s = 407;
	{8'd162,8'd157} : s = 491;
	{8'd162,8'd158} : s = 5;
	{8'd162,8'd159} : s = 38;
	{8'd162,8'd160} : s = 37;
	{8'd162,8'd161} : s = 135;
	{8'd162,8'd162} : s = 35;
	{8'd162,8'd163} : s = 120;
	{8'd162,8'd164} : s = 116;
	{8'd162,8'd165} : s = 244;
	{8'd162,8'd166} : s = 28;
	{8'd162,8'd167} : s = 114;
	{8'd162,8'd168} : s = 113;
	{8'd162,8'd169} : s = 242;
	{8'd162,8'd170} : s = 108;
	{8'd162,8'd171} : s = 241;
	{8'd162,8'd172} : s = 236;
	{8'd162,8'd173} : s = 399;
	{8'd162,8'd174} : s = 26;
	{8'd162,8'd175} : s = 106;
	{8'd162,8'd176} : s = 105;
	{8'd162,8'd177} : s = 234;
	{8'd162,8'd178} : s = 102;
	{8'd162,8'd179} : s = 233;
	{8'd162,8'd180} : s = 230;
	{8'd162,8'd181} : s = 380;
	{8'd162,8'd182} : s = 101;
	{8'd162,8'd183} : s = 229;
	{8'd162,8'd184} : s = 227;
	{8'd162,8'd185} : s = 378;
	{8'd162,8'd186} : s = 220;
	{8'd162,8'd187} : s = 377;
	{8'd162,8'd188} : s = 374;
	{8'd162,8'd189} : s = 487;
	{8'd162,8'd190} : s = 25;
	{8'd162,8'd191} : s = 99;
	{8'd162,8'd192} : s = 92;
	{8'd162,8'd193} : s = 218;
	{8'd162,8'd194} : s = 90;
	{8'd162,8'd195} : s = 217;
	{8'd162,8'd196} : s = 214;
	{8'd162,8'd197} : s = 373;
	{8'd162,8'd198} : s = 89;
	{8'd162,8'd199} : s = 213;
	{8'd162,8'd200} : s = 211;
	{8'd162,8'd201} : s = 371;
	{8'd162,8'd202} : s = 206;
	{8'd162,8'd203} : s = 366;
	{8'd162,8'd204} : s = 365;
	{8'd162,8'd205} : s = 478;
	{8'd162,8'd206} : s = 86;
	{8'd162,8'd207} : s = 205;
	{8'd162,8'd208} : s = 203;
	{8'd162,8'd209} : s = 363;
	{8'd162,8'd210} : s = 199;
	{8'd162,8'd211} : s = 359;
	{8'd162,8'd212} : s = 350;
	{8'd162,8'd213} : s = 477;
	{8'd162,8'd214} : s = 188;
	{8'd162,8'd215} : s = 349;
	{8'd162,8'd216} : s = 347;
	{8'd162,8'd217} : s = 475;
	{8'd162,8'd218} : s = 343;
	{8'd162,8'd219} : s = 471;
	{8'd162,8'd220} : s = 463;
	{8'd162,8'd221} : s = 509;
	{8'd162,8'd222} : s = 3;
	{8'd162,8'd223} : s = 22;
	{8'd162,8'd224} : s = 21;
	{8'd162,8'd225} : s = 85;
	{8'd162,8'd226} : s = 19;
	{8'd162,8'd227} : s = 83;
	{8'd162,8'd228} : s = 78;
	{8'd162,8'd229} : s = 186;
	{8'd162,8'd230} : s = 14;
	{8'd162,8'd231} : s = 77;
	{8'd162,8'd232} : s = 75;
	{8'd162,8'd233} : s = 185;
	{8'd162,8'd234} : s = 71;
	{8'd162,8'd235} : s = 182;
	{8'd162,8'd236} : s = 181;
	{8'd162,8'd237} : s = 335;
	{8'd162,8'd238} : s = 13;
	{8'd162,8'd239} : s = 60;
	{8'd162,8'd240} : s = 58;
	{8'd162,8'd241} : s = 179;
	{8'd162,8'd242} : s = 57;
	{8'd162,8'd243} : s = 174;
	{8'd162,8'd244} : s = 173;
	{8'd162,8'd245} : s = 318;
	{8'd162,8'd246} : s = 54;
	{8'd162,8'd247} : s = 171;
	{8'd162,8'd248} : s = 167;
	{8'd162,8'd249} : s = 317;
	{8'd162,8'd250} : s = 158;
	{8'd162,8'd251} : s = 315;
	{8'd162,8'd252} : s = 311;
	{8'd162,8'd253} : s = 446;
	{8'd162,8'd254} : s = 11;
	{8'd162,8'd255} : s = 53;
	{8'd163,8'd0} : s = 291;
	{8'd163,8'd1} : s = 133;
	{8'd163,8'd2} : s = 284;
	{8'd163,8'd3} : s = 282;
	{8'd163,8'd4} : s = 410;
	{8'd163,8'd5} : s = 131;
	{8'd163,8'd6} : s = 281;
	{8'd163,8'd7} : s = 278;
	{8'd163,8'd8} : s = 409;
	{8'd163,8'd9} : s = 277;
	{8'd163,8'd10} : s = 406;
	{8'd163,8'd11} : s = 405;
	{8'd163,8'd12} : s = 485;
	{8'd163,8'd13} : s = 112;
	{8'd163,8'd14} : s = 275;
	{8'd163,8'd15} : s = 270;
	{8'd163,8'd16} : s = 403;
	{8'd163,8'd17} : s = 269;
	{8'd163,8'd18} : s = 398;
	{8'd163,8'd19} : s = 397;
	{8'd163,8'd20} : s = 483;
	{8'd163,8'd21} : s = 267;
	{8'd163,8'd22} : s = 395;
	{8'd163,8'd23} : s = 391;
	{8'd163,8'd24} : s = 476;
	{8'd163,8'd25} : s = 376;
	{8'd163,8'd26} : s = 474;
	{8'd163,8'd27} : s = 473;
	{8'd163,8'd28} : s = 506;
	{8'd163,8'd29} : s = 20;
	{8'd163,8'd30} : s = 104;
	{8'd163,8'd31} : s = 100;
	{8'd163,8'd32} : s = 263;
	{8'd163,8'd33} : s = 98;
	{8'd163,8'd34} : s = 240;
	{8'd163,8'd35} : s = 232;
	{8'd163,8'd36} : s = 372;
	{8'd163,8'd37} : s = 97;
	{8'd163,8'd38} : s = 228;
	{8'd163,8'd39} : s = 226;
	{8'd163,8'd40} : s = 370;
	{8'd163,8'd41} : s = 225;
	{8'd163,8'd42} : s = 369;
	{8'd163,8'd43} : s = 364;
	{8'd163,8'd44} : s = 470;
	{8'd163,8'd45} : s = 88;
	{8'd163,8'd46} : s = 216;
	{8'd163,8'd47} : s = 212;
	{8'd163,8'd48} : s = 362;
	{8'd163,8'd49} : s = 210;
	{8'd163,8'd50} : s = 361;
	{8'd163,8'd51} : s = 358;
	{8'd163,8'd52} : s = 469;
	{8'd163,8'd53} : s = 209;
	{8'd163,8'd54} : s = 357;
	{8'd163,8'd55} : s = 355;
	{8'd163,8'd56} : s = 467;
	{8'd163,8'd57} : s = 348;
	{8'd163,8'd58} : s = 462;
	{8'd163,8'd59} : s = 461;
	{8'd163,8'd60} : s = 505;
	{8'd163,8'd61} : s = 84;
	{8'd163,8'd62} : s = 204;
	{8'd163,8'd63} : s = 202;
	{8'd163,8'd64} : s = 346;
	{8'd163,8'd65} : s = 201;
	{8'd163,8'd66} : s = 345;
	{8'd163,8'd67} : s = 342;
	{8'd163,8'd68} : s = 459;
	{8'd163,8'd69} : s = 198;
	{8'd163,8'd70} : s = 341;
	{8'd163,8'd71} : s = 339;
	{8'd163,8'd72} : s = 455;
	{8'd163,8'd73} : s = 334;
	{8'd163,8'd74} : s = 444;
	{8'd163,8'd75} : s = 442;
	{8'd163,8'd76} : s = 502;
	{8'd163,8'd77} : s = 197;
	{8'd163,8'd78} : s = 333;
	{8'd163,8'd79} : s = 331;
	{8'd163,8'd80} : s = 441;
	{8'd163,8'd81} : s = 327;
	{8'd163,8'd82} : s = 438;
	{8'd163,8'd83} : s = 437;
	{8'd163,8'd84} : s = 501;
	{8'd163,8'd85} : s = 316;
	{8'd163,8'd86} : s = 435;
	{8'd163,8'd87} : s = 430;
	{8'd163,8'd88} : s = 499;
	{8'd163,8'd89} : s = 429;
	{8'd163,8'd90} : s = 494;
	{8'd163,8'd91} : s = 493;
	{8'd163,8'd92} : s = 510;
	{8'd163,8'd93} : s = 1;
	{8'd163,8'd94} : s = 18;
	{8'd163,8'd95} : s = 17;
	{8'd163,8'd96} : s = 82;
	{8'd163,8'd97} : s = 12;
	{8'd163,8'd98} : s = 81;
	{8'd163,8'd99} : s = 76;
	{8'd163,8'd100} : s = 195;
	{8'd163,8'd101} : s = 10;
	{8'd163,8'd102} : s = 74;
	{8'd163,8'd103} : s = 73;
	{8'd163,8'd104} : s = 184;
	{8'd163,8'd105} : s = 70;
	{8'd163,8'd106} : s = 180;
	{8'd163,8'd107} : s = 178;
	{8'd163,8'd108} : s = 314;
	{8'd163,8'd109} : s = 9;
	{8'd163,8'd110} : s = 69;
	{8'd163,8'd111} : s = 67;
	{8'd163,8'd112} : s = 177;
	{8'd163,8'd113} : s = 56;
	{8'd163,8'd114} : s = 172;
	{8'd163,8'd115} : s = 170;
	{8'd163,8'd116} : s = 313;
	{8'd163,8'd117} : s = 52;
	{8'd163,8'd118} : s = 169;
	{8'd163,8'd119} : s = 166;
	{8'd163,8'd120} : s = 310;
	{8'd163,8'd121} : s = 165;
	{8'd163,8'd122} : s = 309;
	{8'd163,8'd123} : s = 307;
	{8'd163,8'd124} : s = 427;
	{8'd163,8'd125} : s = 6;
	{8'd163,8'd126} : s = 50;
	{8'd163,8'd127} : s = 49;
	{8'd163,8'd128} : s = 163;
	{8'd163,8'd129} : s = 44;
	{8'd163,8'd130} : s = 156;
	{8'd163,8'd131} : s = 154;
	{8'd163,8'd132} : s = 302;
	{8'd163,8'd133} : s = 42;
	{8'd163,8'd134} : s = 153;
	{8'd163,8'd135} : s = 150;
	{8'd163,8'd136} : s = 301;
	{8'd163,8'd137} : s = 149;
	{8'd163,8'd138} : s = 299;
	{8'd163,8'd139} : s = 295;
	{8'd163,8'd140} : s = 423;
	{8'd163,8'd141} : s = 41;
	{8'd163,8'd142} : s = 147;
	{8'd163,8'd143} : s = 142;
	{8'd163,8'd144} : s = 286;
	{8'd163,8'd145} : s = 141;
	{8'd163,8'd146} : s = 285;
	{8'd163,8'd147} : s = 283;
	{8'd163,8'd148} : s = 414;
	{8'd163,8'd149} : s = 139;
	{8'd163,8'd150} : s = 279;
	{8'd163,8'd151} : s = 271;
	{8'd163,8'd152} : s = 413;
	{8'd163,8'd153} : s = 248;
	{8'd163,8'd154} : s = 411;
	{8'd163,8'd155} : s = 407;
	{8'd163,8'd156} : s = 491;
	{8'd163,8'd157} : s = 5;
	{8'd163,8'd158} : s = 38;
	{8'd163,8'd159} : s = 37;
	{8'd163,8'd160} : s = 135;
	{8'd163,8'd161} : s = 35;
	{8'd163,8'd162} : s = 120;
	{8'd163,8'd163} : s = 116;
	{8'd163,8'd164} : s = 244;
	{8'd163,8'd165} : s = 28;
	{8'd163,8'd166} : s = 114;
	{8'd163,8'd167} : s = 113;
	{8'd163,8'd168} : s = 242;
	{8'd163,8'd169} : s = 108;
	{8'd163,8'd170} : s = 241;
	{8'd163,8'd171} : s = 236;
	{8'd163,8'd172} : s = 399;
	{8'd163,8'd173} : s = 26;
	{8'd163,8'd174} : s = 106;
	{8'd163,8'd175} : s = 105;
	{8'd163,8'd176} : s = 234;
	{8'd163,8'd177} : s = 102;
	{8'd163,8'd178} : s = 233;
	{8'd163,8'd179} : s = 230;
	{8'd163,8'd180} : s = 380;
	{8'd163,8'd181} : s = 101;
	{8'd163,8'd182} : s = 229;
	{8'd163,8'd183} : s = 227;
	{8'd163,8'd184} : s = 378;
	{8'd163,8'd185} : s = 220;
	{8'd163,8'd186} : s = 377;
	{8'd163,8'd187} : s = 374;
	{8'd163,8'd188} : s = 487;
	{8'd163,8'd189} : s = 25;
	{8'd163,8'd190} : s = 99;
	{8'd163,8'd191} : s = 92;
	{8'd163,8'd192} : s = 218;
	{8'd163,8'd193} : s = 90;
	{8'd163,8'd194} : s = 217;
	{8'd163,8'd195} : s = 214;
	{8'd163,8'd196} : s = 373;
	{8'd163,8'd197} : s = 89;
	{8'd163,8'd198} : s = 213;
	{8'd163,8'd199} : s = 211;
	{8'd163,8'd200} : s = 371;
	{8'd163,8'd201} : s = 206;
	{8'd163,8'd202} : s = 366;
	{8'd163,8'd203} : s = 365;
	{8'd163,8'd204} : s = 478;
	{8'd163,8'd205} : s = 86;
	{8'd163,8'd206} : s = 205;
	{8'd163,8'd207} : s = 203;
	{8'd163,8'd208} : s = 363;
	{8'd163,8'd209} : s = 199;
	{8'd163,8'd210} : s = 359;
	{8'd163,8'd211} : s = 350;
	{8'd163,8'd212} : s = 477;
	{8'd163,8'd213} : s = 188;
	{8'd163,8'd214} : s = 349;
	{8'd163,8'd215} : s = 347;
	{8'd163,8'd216} : s = 475;
	{8'd163,8'd217} : s = 343;
	{8'd163,8'd218} : s = 471;
	{8'd163,8'd219} : s = 463;
	{8'd163,8'd220} : s = 509;
	{8'd163,8'd221} : s = 3;
	{8'd163,8'd222} : s = 22;
	{8'd163,8'd223} : s = 21;
	{8'd163,8'd224} : s = 85;
	{8'd163,8'd225} : s = 19;
	{8'd163,8'd226} : s = 83;
	{8'd163,8'd227} : s = 78;
	{8'd163,8'd228} : s = 186;
	{8'd163,8'd229} : s = 14;
	{8'd163,8'd230} : s = 77;
	{8'd163,8'd231} : s = 75;
	{8'd163,8'd232} : s = 185;
	{8'd163,8'd233} : s = 71;
	{8'd163,8'd234} : s = 182;
	{8'd163,8'd235} : s = 181;
	{8'd163,8'd236} : s = 335;
	{8'd163,8'd237} : s = 13;
	{8'd163,8'd238} : s = 60;
	{8'd163,8'd239} : s = 58;
	{8'd163,8'd240} : s = 179;
	{8'd163,8'd241} : s = 57;
	{8'd163,8'd242} : s = 174;
	{8'd163,8'd243} : s = 173;
	{8'd163,8'd244} : s = 318;
	{8'd163,8'd245} : s = 54;
	{8'd163,8'd246} : s = 171;
	{8'd163,8'd247} : s = 167;
	{8'd163,8'd248} : s = 317;
	{8'd163,8'd249} : s = 158;
	{8'd163,8'd250} : s = 315;
	{8'd163,8'd251} : s = 311;
	{8'd163,8'd252} : s = 446;
	{8'd163,8'd253} : s = 11;
	{8'd163,8'd254} : s = 53;
	{8'd163,8'd255} : s = 51;
	{8'd164,8'd0} : s = 133;
	{8'd164,8'd1} : s = 284;
	{8'd164,8'd2} : s = 282;
	{8'd164,8'd3} : s = 410;
	{8'd164,8'd4} : s = 131;
	{8'd164,8'd5} : s = 281;
	{8'd164,8'd6} : s = 278;
	{8'd164,8'd7} : s = 409;
	{8'd164,8'd8} : s = 277;
	{8'd164,8'd9} : s = 406;
	{8'd164,8'd10} : s = 405;
	{8'd164,8'd11} : s = 485;
	{8'd164,8'd12} : s = 112;
	{8'd164,8'd13} : s = 275;
	{8'd164,8'd14} : s = 270;
	{8'd164,8'd15} : s = 403;
	{8'd164,8'd16} : s = 269;
	{8'd164,8'd17} : s = 398;
	{8'd164,8'd18} : s = 397;
	{8'd164,8'd19} : s = 483;
	{8'd164,8'd20} : s = 267;
	{8'd164,8'd21} : s = 395;
	{8'd164,8'd22} : s = 391;
	{8'd164,8'd23} : s = 476;
	{8'd164,8'd24} : s = 376;
	{8'd164,8'd25} : s = 474;
	{8'd164,8'd26} : s = 473;
	{8'd164,8'd27} : s = 506;
	{8'd164,8'd28} : s = 20;
	{8'd164,8'd29} : s = 104;
	{8'd164,8'd30} : s = 100;
	{8'd164,8'd31} : s = 263;
	{8'd164,8'd32} : s = 98;
	{8'd164,8'd33} : s = 240;
	{8'd164,8'd34} : s = 232;
	{8'd164,8'd35} : s = 372;
	{8'd164,8'd36} : s = 97;
	{8'd164,8'd37} : s = 228;
	{8'd164,8'd38} : s = 226;
	{8'd164,8'd39} : s = 370;
	{8'd164,8'd40} : s = 225;
	{8'd164,8'd41} : s = 369;
	{8'd164,8'd42} : s = 364;
	{8'd164,8'd43} : s = 470;
	{8'd164,8'd44} : s = 88;
	{8'd164,8'd45} : s = 216;
	{8'd164,8'd46} : s = 212;
	{8'd164,8'd47} : s = 362;
	{8'd164,8'd48} : s = 210;
	{8'd164,8'd49} : s = 361;
	{8'd164,8'd50} : s = 358;
	{8'd164,8'd51} : s = 469;
	{8'd164,8'd52} : s = 209;
	{8'd164,8'd53} : s = 357;
	{8'd164,8'd54} : s = 355;
	{8'd164,8'd55} : s = 467;
	{8'd164,8'd56} : s = 348;
	{8'd164,8'd57} : s = 462;
	{8'd164,8'd58} : s = 461;
	{8'd164,8'd59} : s = 505;
	{8'd164,8'd60} : s = 84;
	{8'd164,8'd61} : s = 204;
	{8'd164,8'd62} : s = 202;
	{8'd164,8'd63} : s = 346;
	{8'd164,8'd64} : s = 201;
	{8'd164,8'd65} : s = 345;
	{8'd164,8'd66} : s = 342;
	{8'd164,8'd67} : s = 459;
	{8'd164,8'd68} : s = 198;
	{8'd164,8'd69} : s = 341;
	{8'd164,8'd70} : s = 339;
	{8'd164,8'd71} : s = 455;
	{8'd164,8'd72} : s = 334;
	{8'd164,8'd73} : s = 444;
	{8'd164,8'd74} : s = 442;
	{8'd164,8'd75} : s = 502;
	{8'd164,8'd76} : s = 197;
	{8'd164,8'd77} : s = 333;
	{8'd164,8'd78} : s = 331;
	{8'd164,8'd79} : s = 441;
	{8'd164,8'd80} : s = 327;
	{8'd164,8'd81} : s = 438;
	{8'd164,8'd82} : s = 437;
	{8'd164,8'd83} : s = 501;
	{8'd164,8'd84} : s = 316;
	{8'd164,8'd85} : s = 435;
	{8'd164,8'd86} : s = 430;
	{8'd164,8'd87} : s = 499;
	{8'd164,8'd88} : s = 429;
	{8'd164,8'd89} : s = 494;
	{8'd164,8'd90} : s = 493;
	{8'd164,8'd91} : s = 510;
	{8'd164,8'd92} : s = 1;
	{8'd164,8'd93} : s = 18;
	{8'd164,8'd94} : s = 17;
	{8'd164,8'd95} : s = 82;
	{8'd164,8'd96} : s = 12;
	{8'd164,8'd97} : s = 81;
	{8'd164,8'd98} : s = 76;
	{8'd164,8'd99} : s = 195;
	{8'd164,8'd100} : s = 10;
	{8'd164,8'd101} : s = 74;
	{8'd164,8'd102} : s = 73;
	{8'd164,8'd103} : s = 184;
	{8'd164,8'd104} : s = 70;
	{8'd164,8'd105} : s = 180;
	{8'd164,8'd106} : s = 178;
	{8'd164,8'd107} : s = 314;
	{8'd164,8'd108} : s = 9;
	{8'd164,8'd109} : s = 69;
	{8'd164,8'd110} : s = 67;
	{8'd164,8'd111} : s = 177;
	{8'd164,8'd112} : s = 56;
	{8'd164,8'd113} : s = 172;
	{8'd164,8'd114} : s = 170;
	{8'd164,8'd115} : s = 313;
	{8'd164,8'd116} : s = 52;
	{8'd164,8'd117} : s = 169;
	{8'd164,8'd118} : s = 166;
	{8'd164,8'd119} : s = 310;
	{8'd164,8'd120} : s = 165;
	{8'd164,8'd121} : s = 309;
	{8'd164,8'd122} : s = 307;
	{8'd164,8'd123} : s = 427;
	{8'd164,8'd124} : s = 6;
	{8'd164,8'd125} : s = 50;
	{8'd164,8'd126} : s = 49;
	{8'd164,8'd127} : s = 163;
	{8'd164,8'd128} : s = 44;
	{8'd164,8'd129} : s = 156;
	{8'd164,8'd130} : s = 154;
	{8'd164,8'd131} : s = 302;
	{8'd164,8'd132} : s = 42;
	{8'd164,8'd133} : s = 153;
	{8'd164,8'd134} : s = 150;
	{8'd164,8'd135} : s = 301;
	{8'd164,8'd136} : s = 149;
	{8'd164,8'd137} : s = 299;
	{8'd164,8'd138} : s = 295;
	{8'd164,8'd139} : s = 423;
	{8'd164,8'd140} : s = 41;
	{8'd164,8'd141} : s = 147;
	{8'd164,8'd142} : s = 142;
	{8'd164,8'd143} : s = 286;
	{8'd164,8'd144} : s = 141;
	{8'd164,8'd145} : s = 285;
	{8'd164,8'd146} : s = 283;
	{8'd164,8'd147} : s = 414;
	{8'd164,8'd148} : s = 139;
	{8'd164,8'd149} : s = 279;
	{8'd164,8'd150} : s = 271;
	{8'd164,8'd151} : s = 413;
	{8'd164,8'd152} : s = 248;
	{8'd164,8'd153} : s = 411;
	{8'd164,8'd154} : s = 407;
	{8'd164,8'd155} : s = 491;
	{8'd164,8'd156} : s = 5;
	{8'd164,8'd157} : s = 38;
	{8'd164,8'd158} : s = 37;
	{8'd164,8'd159} : s = 135;
	{8'd164,8'd160} : s = 35;
	{8'd164,8'd161} : s = 120;
	{8'd164,8'd162} : s = 116;
	{8'd164,8'd163} : s = 244;
	{8'd164,8'd164} : s = 28;
	{8'd164,8'd165} : s = 114;
	{8'd164,8'd166} : s = 113;
	{8'd164,8'd167} : s = 242;
	{8'd164,8'd168} : s = 108;
	{8'd164,8'd169} : s = 241;
	{8'd164,8'd170} : s = 236;
	{8'd164,8'd171} : s = 399;
	{8'd164,8'd172} : s = 26;
	{8'd164,8'd173} : s = 106;
	{8'd164,8'd174} : s = 105;
	{8'd164,8'd175} : s = 234;
	{8'd164,8'd176} : s = 102;
	{8'd164,8'd177} : s = 233;
	{8'd164,8'd178} : s = 230;
	{8'd164,8'd179} : s = 380;
	{8'd164,8'd180} : s = 101;
	{8'd164,8'd181} : s = 229;
	{8'd164,8'd182} : s = 227;
	{8'd164,8'd183} : s = 378;
	{8'd164,8'd184} : s = 220;
	{8'd164,8'd185} : s = 377;
	{8'd164,8'd186} : s = 374;
	{8'd164,8'd187} : s = 487;
	{8'd164,8'd188} : s = 25;
	{8'd164,8'd189} : s = 99;
	{8'd164,8'd190} : s = 92;
	{8'd164,8'd191} : s = 218;
	{8'd164,8'd192} : s = 90;
	{8'd164,8'd193} : s = 217;
	{8'd164,8'd194} : s = 214;
	{8'd164,8'd195} : s = 373;
	{8'd164,8'd196} : s = 89;
	{8'd164,8'd197} : s = 213;
	{8'd164,8'd198} : s = 211;
	{8'd164,8'd199} : s = 371;
	{8'd164,8'd200} : s = 206;
	{8'd164,8'd201} : s = 366;
	{8'd164,8'd202} : s = 365;
	{8'd164,8'd203} : s = 478;
	{8'd164,8'd204} : s = 86;
	{8'd164,8'd205} : s = 205;
	{8'd164,8'd206} : s = 203;
	{8'd164,8'd207} : s = 363;
	{8'd164,8'd208} : s = 199;
	{8'd164,8'd209} : s = 359;
	{8'd164,8'd210} : s = 350;
	{8'd164,8'd211} : s = 477;
	{8'd164,8'd212} : s = 188;
	{8'd164,8'd213} : s = 349;
	{8'd164,8'd214} : s = 347;
	{8'd164,8'd215} : s = 475;
	{8'd164,8'd216} : s = 343;
	{8'd164,8'd217} : s = 471;
	{8'd164,8'd218} : s = 463;
	{8'd164,8'd219} : s = 509;
	{8'd164,8'd220} : s = 3;
	{8'd164,8'd221} : s = 22;
	{8'd164,8'd222} : s = 21;
	{8'd164,8'd223} : s = 85;
	{8'd164,8'd224} : s = 19;
	{8'd164,8'd225} : s = 83;
	{8'd164,8'd226} : s = 78;
	{8'd164,8'd227} : s = 186;
	{8'd164,8'd228} : s = 14;
	{8'd164,8'd229} : s = 77;
	{8'd164,8'd230} : s = 75;
	{8'd164,8'd231} : s = 185;
	{8'd164,8'd232} : s = 71;
	{8'd164,8'd233} : s = 182;
	{8'd164,8'd234} : s = 181;
	{8'd164,8'd235} : s = 335;
	{8'd164,8'd236} : s = 13;
	{8'd164,8'd237} : s = 60;
	{8'd164,8'd238} : s = 58;
	{8'd164,8'd239} : s = 179;
	{8'd164,8'd240} : s = 57;
	{8'd164,8'd241} : s = 174;
	{8'd164,8'd242} : s = 173;
	{8'd164,8'd243} : s = 318;
	{8'd164,8'd244} : s = 54;
	{8'd164,8'd245} : s = 171;
	{8'd164,8'd246} : s = 167;
	{8'd164,8'd247} : s = 317;
	{8'd164,8'd248} : s = 158;
	{8'd164,8'd249} : s = 315;
	{8'd164,8'd250} : s = 311;
	{8'd164,8'd251} : s = 446;
	{8'd164,8'd252} : s = 11;
	{8'd164,8'd253} : s = 53;
	{8'd164,8'd254} : s = 51;
	{8'd164,8'd255} : s = 157;
	{8'd165,8'd0} : s = 284;
	{8'd165,8'd1} : s = 282;
	{8'd165,8'd2} : s = 410;
	{8'd165,8'd3} : s = 131;
	{8'd165,8'd4} : s = 281;
	{8'd165,8'd5} : s = 278;
	{8'd165,8'd6} : s = 409;
	{8'd165,8'd7} : s = 277;
	{8'd165,8'd8} : s = 406;
	{8'd165,8'd9} : s = 405;
	{8'd165,8'd10} : s = 485;
	{8'd165,8'd11} : s = 112;
	{8'd165,8'd12} : s = 275;
	{8'd165,8'd13} : s = 270;
	{8'd165,8'd14} : s = 403;
	{8'd165,8'd15} : s = 269;
	{8'd165,8'd16} : s = 398;
	{8'd165,8'd17} : s = 397;
	{8'd165,8'd18} : s = 483;
	{8'd165,8'd19} : s = 267;
	{8'd165,8'd20} : s = 395;
	{8'd165,8'd21} : s = 391;
	{8'd165,8'd22} : s = 476;
	{8'd165,8'd23} : s = 376;
	{8'd165,8'd24} : s = 474;
	{8'd165,8'd25} : s = 473;
	{8'd165,8'd26} : s = 506;
	{8'd165,8'd27} : s = 20;
	{8'd165,8'd28} : s = 104;
	{8'd165,8'd29} : s = 100;
	{8'd165,8'd30} : s = 263;
	{8'd165,8'd31} : s = 98;
	{8'd165,8'd32} : s = 240;
	{8'd165,8'd33} : s = 232;
	{8'd165,8'd34} : s = 372;
	{8'd165,8'd35} : s = 97;
	{8'd165,8'd36} : s = 228;
	{8'd165,8'd37} : s = 226;
	{8'd165,8'd38} : s = 370;
	{8'd165,8'd39} : s = 225;
	{8'd165,8'd40} : s = 369;
	{8'd165,8'd41} : s = 364;
	{8'd165,8'd42} : s = 470;
	{8'd165,8'd43} : s = 88;
	{8'd165,8'd44} : s = 216;
	{8'd165,8'd45} : s = 212;
	{8'd165,8'd46} : s = 362;
	{8'd165,8'd47} : s = 210;
	{8'd165,8'd48} : s = 361;
	{8'd165,8'd49} : s = 358;
	{8'd165,8'd50} : s = 469;
	{8'd165,8'd51} : s = 209;
	{8'd165,8'd52} : s = 357;
	{8'd165,8'd53} : s = 355;
	{8'd165,8'd54} : s = 467;
	{8'd165,8'd55} : s = 348;
	{8'd165,8'd56} : s = 462;
	{8'd165,8'd57} : s = 461;
	{8'd165,8'd58} : s = 505;
	{8'd165,8'd59} : s = 84;
	{8'd165,8'd60} : s = 204;
	{8'd165,8'd61} : s = 202;
	{8'd165,8'd62} : s = 346;
	{8'd165,8'd63} : s = 201;
	{8'd165,8'd64} : s = 345;
	{8'd165,8'd65} : s = 342;
	{8'd165,8'd66} : s = 459;
	{8'd165,8'd67} : s = 198;
	{8'd165,8'd68} : s = 341;
	{8'd165,8'd69} : s = 339;
	{8'd165,8'd70} : s = 455;
	{8'd165,8'd71} : s = 334;
	{8'd165,8'd72} : s = 444;
	{8'd165,8'd73} : s = 442;
	{8'd165,8'd74} : s = 502;
	{8'd165,8'd75} : s = 197;
	{8'd165,8'd76} : s = 333;
	{8'd165,8'd77} : s = 331;
	{8'd165,8'd78} : s = 441;
	{8'd165,8'd79} : s = 327;
	{8'd165,8'd80} : s = 438;
	{8'd165,8'd81} : s = 437;
	{8'd165,8'd82} : s = 501;
	{8'd165,8'd83} : s = 316;
	{8'd165,8'd84} : s = 435;
	{8'd165,8'd85} : s = 430;
	{8'd165,8'd86} : s = 499;
	{8'd165,8'd87} : s = 429;
	{8'd165,8'd88} : s = 494;
	{8'd165,8'd89} : s = 493;
	{8'd165,8'd90} : s = 510;
	{8'd165,8'd91} : s = 1;
	{8'd165,8'd92} : s = 18;
	{8'd165,8'd93} : s = 17;
	{8'd165,8'd94} : s = 82;
	{8'd165,8'd95} : s = 12;
	{8'd165,8'd96} : s = 81;
	{8'd165,8'd97} : s = 76;
	{8'd165,8'd98} : s = 195;
	{8'd165,8'd99} : s = 10;
	{8'd165,8'd100} : s = 74;
	{8'd165,8'd101} : s = 73;
	{8'd165,8'd102} : s = 184;
	{8'd165,8'd103} : s = 70;
	{8'd165,8'd104} : s = 180;
	{8'd165,8'd105} : s = 178;
	{8'd165,8'd106} : s = 314;
	{8'd165,8'd107} : s = 9;
	{8'd165,8'd108} : s = 69;
	{8'd165,8'd109} : s = 67;
	{8'd165,8'd110} : s = 177;
	{8'd165,8'd111} : s = 56;
	{8'd165,8'd112} : s = 172;
	{8'd165,8'd113} : s = 170;
	{8'd165,8'd114} : s = 313;
	{8'd165,8'd115} : s = 52;
	{8'd165,8'd116} : s = 169;
	{8'd165,8'd117} : s = 166;
	{8'd165,8'd118} : s = 310;
	{8'd165,8'd119} : s = 165;
	{8'd165,8'd120} : s = 309;
	{8'd165,8'd121} : s = 307;
	{8'd165,8'd122} : s = 427;
	{8'd165,8'd123} : s = 6;
	{8'd165,8'd124} : s = 50;
	{8'd165,8'd125} : s = 49;
	{8'd165,8'd126} : s = 163;
	{8'd165,8'd127} : s = 44;
	{8'd165,8'd128} : s = 156;
	{8'd165,8'd129} : s = 154;
	{8'd165,8'd130} : s = 302;
	{8'd165,8'd131} : s = 42;
	{8'd165,8'd132} : s = 153;
	{8'd165,8'd133} : s = 150;
	{8'd165,8'd134} : s = 301;
	{8'd165,8'd135} : s = 149;
	{8'd165,8'd136} : s = 299;
	{8'd165,8'd137} : s = 295;
	{8'd165,8'd138} : s = 423;
	{8'd165,8'd139} : s = 41;
	{8'd165,8'd140} : s = 147;
	{8'd165,8'd141} : s = 142;
	{8'd165,8'd142} : s = 286;
	{8'd165,8'd143} : s = 141;
	{8'd165,8'd144} : s = 285;
	{8'd165,8'd145} : s = 283;
	{8'd165,8'd146} : s = 414;
	{8'd165,8'd147} : s = 139;
	{8'd165,8'd148} : s = 279;
	{8'd165,8'd149} : s = 271;
	{8'd165,8'd150} : s = 413;
	{8'd165,8'd151} : s = 248;
	{8'd165,8'd152} : s = 411;
	{8'd165,8'd153} : s = 407;
	{8'd165,8'd154} : s = 491;
	{8'd165,8'd155} : s = 5;
	{8'd165,8'd156} : s = 38;
	{8'd165,8'd157} : s = 37;
	{8'd165,8'd158} : s = 135;
	{8'd165,8'd159} : s = 35;
	{8'd165,8'd160} : s = 120;
	{8'd165,8'd161} : s = 116;
	{8'd165,8'd162} : s = 244;
	{8'd165,8'd163} : s = 28;
	{8'd165,8'd164} : s = 114;
	{8'd165,8'd165} : s = 113;
	{8'd165,8'd166} : s = 242;
	{8'd165,8'd167} : s = 108;
	{8'd165,8'd168} : s = 241;
	{8'd165,8'd169} : s = 236;
	{8'd165,8'd170} : s = 399;
	{8'd165,8'd171} : s = 26;
	{8'd165,8'd172} : s = 106;
	{8'd165,8'd173} : s = 105;
	{8'd165,8'd174} : s = 234;
	{8'd165,8'd175} : s = 102;
	{8'd165,8'd176} : s = 233;
	{8'd165,8'd177} : s = 230;
	{8'd165,8'd178} : s = 380;
	{8'd165,8'd179} : s = 101;
	{8'd165,8'd180} : s = 229;
	{8'd165,8'd181} : s = 227;
	{8'd165,8'd182} : s = 378;
	{8'd165,8'd183} : s = 220;
	{8'd165,8'd184} : s = 377;
	{8'd165,8'd185} : s = 374;
	{8'd165,8'd186} : s = 487;
	{8'd165,8'd187} : s = 25;
	{8'd165,8'd188} : s = 99;
	{8'd165,8'd189} : s = 92;
	{8'd165,8'd190} : s = 218;
	{8'd165,8'd191} : s = 90;
	{8'd165,8'd192} : s = 217;
	{8'd165,8'd193} : s = 214;
	{8'd165,8'd194} : s = 373;
	{8'd165,8'd195} : s = 89;
	{8'd165,8'd196} : s = 213;
	{8'd165,8'd197} : s = 211;
	{8'd165,8'd198} : s = 371;
	{8'd165,8'd199} : s = 206;
	{8'd165,8'd200} : s = 366;
	{8'd165,8'd201} : s = 365;
	{8'd165,8'd202} : s = 478;
	{8'd165,8'd203} : s = 86;
	{8'd165,8'd204} : s = 205;
	{8'd165,8'd205} : s = 203;
	{8'd165,8'd206} : s = 363;
	{8'd165,8'd207} : s = 199;
	{8'd165,8'd208} : s = 359;
	{8'd165,8'd209} : s = 350;
	{8'd165,8'd210} : s = 477;
	{8'd165,8'd211} : s = 188;
	{8'd165,8'd212} : s = 349;
	{8'd165,8'd213} : s = 347;
	{8'd165,8'd214} : s = 475;
	{8'd165,8'd215} : s = 343;
	{8'd165,8'd216} : s = 471;
	{8'd165,8'd217} : s = 463;
	{8'd165,8'd218} : s = 509;
	{8'd165,8'd219} : s = 3;
	{8'd165,8'd220} : s = 22;
	{8'd165,8'd221} : s = 21;
	{8'd165,8'd222} : s = 85;
	{8'd165,8'd223} : s = 19;
	{8'd165,8'd224} : s = 83;
	{8'd165,8'd225} : s = 78;
	{8'd165,8'd226} : s = 186;
	{8'd165,8'd227} : s = 14;
	{8'd165,8'd228} : s = 77;
	{8'd165,8'd229} : s = 75;
	{8'd165,8'd230} : s = 185;
	{8'd165,8'd231} : s = 71;
	{8'd165,8'd232} : s = 182;
	{8'd165,8'd233} : s = 181;
	{8'd165,8'd234} : s = 335;
	{8'd165,8'd235} : s = 13;
	{8'd165,8'd236} : s = 60;
	{8'd165,8'd237} : s = 58;
	{8'd165,8'd238} : s = 179;
	{8'd165,8'd239} : s = 57;
	{8'd165,8'd240} : s = 174;
	{8'd165,8'd241} : s = 173;
	{8'd165,8'd242} : s = 318;
	{8'd165,8'd243} : s = 54;
	{8'd165,8'd244} : s = 171;
	{8'd165,8'd245} : s = 167;
	{8'd165,8'd246} : s = 317;
	{8'd165,8'd247} : s = 158;
	{8'd165,8'd248} : s = 315;
	{8'd165,8'd249} : s = 311;
	{8'd165,8'd250} : s = 446;
	{8'd165,8'd251} : s = 11;
	{8'd165,8'd252} : s = 53;
	{8'd165,8'd253} : s = 51;
	{8'd165,8'd254} : s = 157;
	{8'd165,8'd255} : s = 46;
	{8'd166,8'd0} : s = 282;
	{8'd166,8'd1} : s = 410;
	{8'd166,8'd2} : s = 131;
	{8'd166,8'd3} : s = 281;
	{8'd166,8'd4} : s = 278;
	{8'd166,8'd5} : s = 409;
	{8'd166,8'd6} : s = 277;
	{8'd166,8'd7} : s = 406;
	{8'd166,8'd8} : s = 405;
	{8'd166,8'd9} : s = 485;
	{8'd166,8'd10} : s = 112;
	{8'd166,8'd11} : s = 275;
	{8'd166,8'd12} : s = 270;
	{8'd166,8'd13} : s = 403;
	{8'd166,8'd14} : s = 269;
	{8'd166,8'd15} : s = 398;
	{8'd166,8'd16} : s = 397;
	{8'd166,8'd17} : s = 483;
	{8'd166,8'd18} : s = 267;
	{8'd166,8'd19} : s = 395;
	{8'd166,8'd20} : s = 391;
	{8'd166,8'd21} : s = 476;
	{8'd166,8'd22} : s = 376;
	{8'd166,8'd23} : s = 474;
	{8'd166,8'd24} : s = 473;
	{8'd166,8'd25} : s = 506;
	{8'd166,8'd26} : s = 20;
	{8'd166,8'd27} : s = 104;
	{8'd166,8'd28} : s = 100;
	{8'd166,8'd29} : s = 263;
	{8'd166,8'd30} : s = 98;
	{8'd166,8'd31} : s = 240;
	{8'd166,8'd32} : s = 232;
	{8'd166,8'd33} : s = 372;
	{8'd166,8'd34} : s = 97;
	{8'd166,8'd35} : s = 228;
	{8'd166,8'd36} : s = 226;
	{8'd166,8'd37} : s = 370;
	{8'd166,8'd38} : s = 225;
	{8'd166,8'd39} : s = 369;
	{8'd166,8'd40} : s = 364;
	{8'd166,8'd41} : s = 470;
	{8'd166,8'd42} : s = 88;
	{8'd166,8'd43} : s = 216;
	{8'd166,8'd44} : s = 212;
	{8'd166,8'd45} : s = 362;
	{8'd166,8'd46} : s = 210;
	{8'd166,8'd47} : s = 361;
	{8'd166,8'd48} : s = 358;
	{8'd166,8'd49} : s = 469;
	{8'd166,8'd50} : s = 209;
	{8'd166,8'd51} : s = 357;
	{8'd166,8'd52} : s = 355;
	{8'd166,8'd53} : s = 467;
	{8'd166,8'd54} : s = 348;
	{8'd166,8'd55} : s = 462;
	{8'd166,8'd56} : s = 461;
	{8'd166,8'd57} : s = 505;
	{8'd166,8'd58} : s = 84;
	{8'd166,8'd59} : s = 204;
	{8'd166,8'd60} : s = 202;
	{8'd166,8'd61} : s = 346;
	{8'd166,8'd62} : s = 201;
	{8'd166,8'd63} : s = 345;
	{8'd166,8'd64} : s = 342;
	{8'd166,8'd65} : s = 459;
	{8'd166,8'd66} : s = 198;
	{8'd166,8'd67} : s = 341;
	{8'd166,8'd68} : s = 339;
	{8'd166,8'd69} : s = 455;
	{8'd166,8'd70} : s = 334;
	{8'd166,8'd71} : s = 444;
	{8'd166,8'd72} : s = 442;
	{8'd166,8'd73} : s = 502;
	{8'd166,8'd74} : s = 197;
	{8'd166,8'd75} : s = 333;
	{8'd166,8'd76} : s = 331;
	{8'd166,8'd77} : s = 441;
	{8'd166,8'd78} : s = 327;
	{8'd166,8'd79} : s = 438;
	{8'd166,8'd80} : s = 437;
	{8'd166,8'd81} : s = 501;
	{8'd166,8'd82} : s = 316;
	{8'd166,8'd83} : s = 435;
	{8'd166,8'd84} : s = 430;
	{8'd166,8'd85} : s = 499;
	{8'd166,8'd86} : s = 429;
	{8'd166,8'd87} : s = 494;
	{8'd166,8'd88} : s = 493;
	{8'd166,8'd89} : s = 510;
	{8'd166,8'd90} : s = 1;
	{8'd166,8'd91} : s = 18;
	{8'd166,8'd92} : s = 17;
	{8'd166,8'd93} : s = 82;
	{8'd166,8'd94} : s = 12;
	{8'd166,8'd95} : s = 81;
	{8'd166,8'd96} : s = 76;
	{8'd166,8'd97} : s = 195;
	{8'd166,8'd98} : s = 10;
	{8'd166,8'd99} : s = 74;
	{8'd166,8'd100} : s = 73;
	{8'd166,8'd101} : s = 184;
	{8'd166,8'd102} : s = 70;
	{8'd166,8'd103} : s = 180;
	{8'd166,8'd104} : s = 178;
	{8'd166,8'd105} : s = 314;
	{8'd166,8'd106} : s = 9;
	{8'd166,8'd107} : s = 69;
	{8'd166,8'd108} : s = 67;
	{8'd166,8'd109} : s = 177;
	{8'd166,8'd110} : s = 56;
	{8'd166,8'd111} : s = 172;
	{8'd166,8'd112} : s = 170;
	{8'd166,8'd113} : s = 313;
	{8'd166,8'd114} : s = 52;
	{8'd166,8'd115} : s = 169;
	{8'd166,8'd116} : s = 166;
	{8'd166,8'd117} : s = 310;
	{8'd166,8'd118} : s = 165;
	{8'd166,8'd119} : s = 309;
	{8'd166,8'd120} : s = 307;
	{8'd166,8'd121} : s = 427;
	{8'd166,8'd122} : s = 6;
	{8'd166,8'd123} : s = 50;
	{8'd166,8'd124} : s = 49;
	{8'd166,8'd125} : s = 163;
	{8'd166,8'd126} : s = 44;
	{8'd166,8'd127} : s = 156;
	{8'd166,8'd128} : s = 154;
	{8'd166,8'd129} : s = 302;
	{8'd166,8'd130} : s = 42;
	{8'd166,8'd131} : s = 153;
	{8'd166,8'd132} : s = 150;
	{8'd166,8'd133} : s = 301;
	{8'd166,8'd134} : s = 149;
	{8'd166,8'd135} : s = 299;
	{8'd166,8'd136} : s = 295;
	{8'd166,8'd137} : s = 423;
	{8'd166,8'd138} : s = 41;
	{8'd166,8'd139} : s = 147;
	{8'd166,8'd140} : s = 142;
	{8'd166,8'd141} : s = 286;
	{8'd166,8'd142} : s = 141;
	{8'd166,8'd143} : s = 285;
	{8'd166,8'd144} : s = 283;
	{8'd166,8'd145} : s = 414;
	{8'd166,8'd146} : s = 139;
	{8'd166,8'd147} : s = 279;
	{8'd166,8'd148} : s = 271;
	{8'd166,8'd149} : s = 413;
	{8'd166,8'd150} : s = 248;
	{8'd166,8'd151} : s = 411;
	{8'd166,8'd152} : s = 407;
	{8'd166,8'd153} : s = 491;
	{8'd166,8'd154} : s = 5;
	{8'd166,8'd155} : s = 38;
	{8'd166,8'd156} : s = 37;
	{8'd166,8'd157} : s = 135;
	{8'd166,8'd158} : s = 35;
	{8'd166,8'd159} : s = 120;
	{8'd166,8'd160} : s = 116;
	{8'd166,8'd161} : s = 244;
	{8'd166,8'd162} : s = 28;
	{8'd166,8'd163} : s = 114;
	{8'd166,8'd164} : s = 113;
	{8'd166,8'd165} : s = 242;
	{8'd166,8'd166} : s = 108;
	{8'd166,8'd167} : s = 241;
	{8'd166,8'd168} : s = 236;
	{8'd166,8'd169} : s = 399;
	{8'd166,8'd170} : s = 26;
	{8'd166,8'd171} : s = 106;
	{8'd166,8'd172} : s = 105;
	{8'd166,8'd173} : s = 234;
	{8'd166,8'd174} : s = 102;
	{8'd166,8'd175} : s = 233;
	{8'd166,8'd176} : s = 230;
	{8'd166,8'd177} : s = 380;
	{8'd166,8'd178} : s = 101;
	{8'd166,8'd179} : s = 229;
	{8'd166,8'd180} : s = 227;
	{8'd166,8'd181} : s = 378;
	{8'd166,8'd182} : s = 220;
	{8'd166,8'd183} : s = 377;
	{8'd166,8'd184} : s = 374;
	{8'd166,8'd185} : s = 487;
	{8'd166,8'd186} : s = 25;
	{8'd166,8'd187} : s = 99;
	{8'd166,8'd188} : s = 92;
	{8'd166,8'd189} : s = 218;
	{8'd166,8'd190} : s = 90;
	{8'd166,8'd191} : s = 217;
	{8'd166,8'd192} : s = 214;
	{8'd166,8'd193} : s = 373;
	{8'd166,8'd194} : s = 89;
	{8'd166,8'd195} : s = 213;
	{8'd166,8'd196} : s = 211;
	{8'd166,8'd197} : s = 371;
	{8'd166,8'd198} : s = 206;
	{8'd166,8'd199} : s = 366;
	{8'd166,8'd200} : s = 365;
	{8'd166,8'd201} : s = 478;
	{8'd166,8'd202} : s = 86;
	{8'd166,8'd203} : s = 205;
	{8'd166,8'd204} : s = 203;
	{8'd166,8'd205} : s = 363;
	{8'd166,8'd206} : s = 199;
	{8'd166,8'd207} : s = 359;
	{8'd166,8'd208} : s = 350;
	{8'd166,8'd209} : s = 477;
	{8'd166,8'd210} : s = 188;
	{8'd166,8'd211} : s = 349;
	{8'd166,8'd212} : s = 347;
	{8'd166,8'd213} : s = 475;
	{8'd166,8'd214} : s = 343;
	{8'd166,8'd215} : s = 471;
	{8'd166,8'd216} : s = 463;
	{8'd166,8'd217} : s = 509;
	{8'd166,8'd218} : s = 3;
	{8'd166,8'd219} : s = 22;
	{8'd166,8'd220} : s = 21;
	{8'd166,8'd221} : s = 85;
	{8'd166,8'd222} : s = 19;
	{8'd166,8'd223} : s = 83;
	{8'd166,8'd224} : s = 78;
	{8'd166,8'd225} : s = 186;
	{8'd166,8'd226} : s = 14;
	{8'd166,8'd227} : s = 77;
	{8'd166,8'd228} : s = 75;
	{8'd166,8'd229} : s = 185;
	{8'd166,8'd230} : s = 71;
	{8'd166,8'd231} : s = 182;
	{8'd166,8'd232} : s = 181;
	{8'd166,8'd233} : s = 335;
	{8'd166,8'd234} : s = 13;
	{8'd166,8'd235} : s = 60;
	{8'd166,8'd236} : s = 58;
	{8'd166,8'd237} : s = 179;
	{8'd166,8'd238} : s = 57;
	{8'd166,8'd239} : s = 174;
	{8'd166,8'd240} : s = 173;
	{8'd166,8'd241} : s = 318;
	{8'd166,8'd242} : s = 54;
	{8'd166,8'd243} : s = 171;
	{8'd166,8'd244} : s = 167;
	{8'd166,8'd245} : s = 317;
	{8'd166,8'd246} : s = 158;
	{8'd166,8'd247} : s = 315;
	{8'd166,8'd248} : s = 311;
	{8'd166,8'd249} : s = 446;
	{8'd166,8'd250} : s = 11;
	{8'd166,8'd251} : s = 53;
	{8'd166,8'd252} : s = 51;
	{8'd166,8'd253} : s = 157;
	{8'd166,8'd254} : s = 46;
	{8'd166,8'd255} : s = 155;
	{8'd167,8'd0} : s = 410;
	{8'd167,8'd1} : s = 131;
	{8'd167,8'd2} : s = 281;
	{8'd167,8'd3} : s = 278;
	{8'd167,8'd4} : s = 409;
	{8'd167,8'd5} : s = 277;
	{8'd167,8'd6} : s = 406;
	{8'd167,8'd7} : s = 405;
	{8'd167,8'd8} : s = 485;
	{8'd167,8'd9} : s = 112;
	{8'd167,8'd10} : s = 275;
	{8'd167,8'd11} : s = 270;
	{8'd167,8'd12} : s = 403;
	{8'd167,8'd13} : s = 269;
	{8'd167,8'd14} : s = 398;
	{8'd167,8'd15} : s = 397;
	{8'd167,8'd16} : s = 483;
	{8'd167,8'd17} : s = 267;
	{8'd167,8'd18} : s = 395;
	{8'd167,8'd19} : s = 391;
	{8'd167,8'd20} : s = 476;
	{8'd167,8'd21} : s = 376;
	{8'd167,8'd22} : s = 474;
	{8'd167,8'd23} : s = 473;
	{8'd167,8'd24} : s = 506;
	{8'd167,8'd25} : s = 20;
	{8'd167,8'd26} : s = 104;
	{8'd167,8'd27} : s = 100;
	{8'd167,8'd28} : s = 263;
	{8'd167,8'd29} : s = 98;
	{8'd167,8'd30} : s = 240;
	{8'd167,8'd31} : s = 232;
	{8'd167,8'd32} : s = 372;
	{8'd167,8'd33} : s = 97;
	{8'd167,8'd34} : s = 228;
	{8'd167,8'd35} : s = 226;
	{8'd167,8'd36} : s = 370;
	{8'd167,8'd37} : s = 225;
	{8'd167,8'd38} : s = 369;
	{8'd167,8'd39} : s = 364;
	{8'd167,8'd40} : s = 470;
	{8'd167,8'd41} : s = 88;
	{8'd167,8'd42} : s = 216;
	{8'd167,8'd43} : s = 212;
	{8'd167,8'd44} : s = 362;
	{8'd167,8'd45} : s = 210;
	{8'd167,8'd46} : s = 361;
	{8'd167,8'd47} : s = 358;
	{8'd167,8'd48} : s = 469;
	{8'd167,8'd49} : s = 209;
	{8'd167,8'd50} : s = 357;
	{8'd167,8'd51} : s = 355;
	{8'd167,8'd52} : s = 467;
	{8'd167,8'd53} : s = 348;
	{8'd167,8'd54} : s = 462;
	{8'd167,8'd55} : s = 461;
	{8'd167,8'd56} : s = 505;
	{8'd167,8'd57} : s = 84;
	{8'd167,8'd58} : s = 204;
	{8'd167,8'd59} : s = 202;
	{8'd167,8'd60} : s = 346;
	{8'd167,8'd61} : s = 201;
	{8'd167,8'd62} : s = 345;
	{8'd167,8'd63} : s = 342;
	{8'd167,8'd64} : s = 459;
	{8'd167,8'd65} : s = 198;
	{8'd167,8'd66} : s = 341;
	{8'd167,8'd67} : s = 339;
	{8'd167,8'd68} : s = 455;
	{8'd167,8'd69} : s = 334;
	{8'd167,8'd70} : s = 444;
	{8'd167,8'd71} : s = 442;
	{8'd167,8'd72} : s = 502;
	{8'd167,8'd73} : s = 197;
	{8'd167,8'd74} : s = 333;
	{8'd167,8'd75} : s = 331;
	{8'd167,8'd76} : s = 441;
	{8'd167,8'd77} : s = 327;
	{8'd167,8'd78} : s = 438;
	{8'd167,8'd79} : s = 437;
	{8'd167,8'd80} : s = 501;
	{8'd167,8'd81} : s = 316;
	{8'd167,8'd82} : s = 435;
	{8'd167,8'd83} : s = 430;
	{8'd167,8'd84} : s = 499;
	{8'd167,8'd85} : s = 429;
	{8'd167,8'd86} : s = 494;
	{8'd167,8'd87} : s = 493;
	{8'd167,8'd88} : s = 510;
	{8'd167,8'd89} : s = 1;
	{8'd167,8'd90} : s = 18;
	{8'd167,8'd91} : s = 17;
	{8'd167,8'd92} : s = 82;
	{8'd167,8'd93} : s = 12;
	{8'd167,8'd94} : s = 81;
	{8'd167,8'd95} : s = 76;
	{8'd167,8'd96} : s = 195;
	{8'd167,8'd97} : s = 10;
	{8'd167,8'd98} : s = 74;
	{8'd167,8'd99} : s = 73;
	{8'd167,8'd100} : s = 184;
	{8'd167,8'd101} : s = 70;
	{8'd167,8'd102} : s = 180;
	{8'd167,8'd103} : s = 178;
	{8'd167,8'd104} : s = 314;
	{8'd167,8'd105} : s = 9;
	{8'd167,8'd106} : s = 69;
	{8'd167,8'd107} : s = 67;
	{8'd167,8'd108} : s = 177;
	{8'd167,8'd109} : s = 56;
	{8'd167,8'd110} : s = 172;
	{8'd167,8'd111} : s = 170;
	{8'd167,8'd112} : s = 313;
	{8'd167,8'd113} : s = 52;
	{8'd167,8'd114} : s = 169;
	{8'd167,8'd115} : s = 166;
	{8'd167,8'd116} : s = 310;
	{8'd167,8'd117} : s = 165;
	{8'd167,8'd118} : s = 309;
	{8'd167,8'd119} : s = 307;
	{8'd167,8'd120} : s = 427;
	{8'd167,8'd121} : s = 6;
	{8'd167,8'd122} : s = 50;
	{8'd167,8'd123} : s = 49;
	{8'd167,8'd124} : s = 163;
	{8'd167,8'd125} : s = 44;
	{8'd167,8'd126} : s = 156;
	{8'd167,8'd127} : s = 154;
	{8'd167,8'd128} : s = 302;
	{8'd167,8'd129} : s = 42;
	{8'd167,8'd130} : s = 153;
	{8'd167,8'd131} : s = 150;
	{8'd167,8'd132} : s = 301;
	{8'd167,8'd133} : s = 149;
	{8'd167,8'd134} : s = 299;
	{8'd167,8'd135} : s = 295;
	{8'd167,8'd136} : s = 423;
	{8'd167,8'd137} : s = 41;
	{8'd167,8'd138} : s = 147;
	{8'd167,8'd139} : s = 142;
	{8'd167,8'd140} : s = 286;
	{8'd167,8'd141} : s = 141;
	{8'd167,8'd142} : s = 285;
	{8'd167,8'd143} : s = 283;
	{8'd167,8'd144} : s = 414;
	{8'd167,8'd145} : s = 139;
	{8'd167,8'd146} : s = 279;
	{8'd167,8'd147} : s = 271;
	{8'd167,8'd148} : s = 413;
	{8'd167,8'd149} : s = 248;
	{8'd167,8'd150} : s = 411;
	{8'd167,8'd151} : s = 407;
	{8'd167,8'd152} : s = 491;
	{8'd167,8'd153} : s = 5;
	{8'd167,8'd154} : s = 38;
	{8'd167,8'd155} : s = 37;
	{8'd167,8'd156} : s = 135;
	{8'd167,8'd157} : s = 35;
	{8'd167,8'd158} : s = 120;
	{8'd167,8'd159} : s = 116;
	{8'd167,8'd160} : s = 244;
	{8'd167,8'd161} : s = 28;
	{8'd167,8'd162} : s = 114;
	{8'd167,8'd163} : s = 113;
	{8'd167,8'd164} : s = 242;
	{8'd167,8'd165} : s = 108;
	{8'd167,8'd166} : s = 241;
	{8'd167,8'd167} : s = 236;
	{8'd167,8'd168} : s = 399;
	{8'd167,8'd169} : s = 26;
	{8'd167,8'd170} : s = 106;
	{8'd167,8'd171} : s = 105;
	{8'd167,8'd172} : s = 234;
	{8'd167,8'd173} : s = 102;
	{8'd167,8'd174} : s = 233;
	{8'd167,8'd175} : s = 230;
	{8'd167,8'd176} : s = 380;
	{8'd167,8'd177} : s = 101;
	{8'd167,8'd178} : s = 229;
	{8'd167,8'd179} : s = 227;
	{8'd167,8'd180} : s = 378;
	{8'd167,8'd181} : s = 220;
	{8'd167,8'd182} : s = 377;
	{8'd167,8'd183} : s = 374;
	{8'd167,8'd184} : s = 487;
	{8'd167,8'd185} : s = 25;
	{8'd167,8'd186} : s = 99;
	{8'd167,8'd187} : s = 92;
	{8'd167,8'd188} : s = 218;
	{8'd167,8'd189} : s = 90;
	{8'd167,8'd190} : s = 217;
	{8'd167,8'd191} : s = 214;
	{8'd167,8'd192} : s = 373;
	{8'd167,8'd193} : s = 89;
	{8'd167,8'd194} : s = 213;
	{8'd167,8'd195} : s = 211;
	{8'd167,8'd196} : s = 371;
	{8'd167,8'd197} : s = 206;
	{8'd167,8'd198} : s = 366;
	{8'd167,8'd199} : s = 365;
	{8'd167,8'd200} : s = 478;
	{8'd167,8'd201} : s = 86;
	{8'd167,8'd202} : s = 205;
	{8'd167,8'd203} : s = 203;
	{8'd167,8'd204} : s = 363;
	{8'd167,8'd205} : s = 199;
	{8'd167,8'd206} : s = 359;
	{8'd167,8'd207} : s = 350;
	{8'd167,8'd208} : s = 477;
	{8'd167,8'd209} : s = 188;
	{8'd167,8'd210} : s = 349;
	{8'd167,8'd211} : s = 347;
	{8'd167,8'd212} : s = 475;
	{8'd167,8'd213} : s = 343;
	{8'd167,8'd214} : s = 471;
	{8'd167,8'd215} : s = 463;
	{8'd167,8'd216} : s = 509;
	{8'd167,8'd217} : s = 3;
	{8'd167,8'd218} : s = 22;
	{8'd167,8'd219} : s = 21;
	{8'd167,8'd220} : s = 85;
	{8'd167,8'd221} : s = 19;
	{8'd167,8'd222} : s = 83;
	{8'd167,8'd223} : s = 78;
	{8'd167,8'd224} : s = 186;
	{8'd167,8'd225} : s = 14;
	{8'd167,8'd226} : s = 77;
	{8'd167,8'd227} : s = 75;
	{8'd167,8'd228} : s = 185;
	{8'd167,8'd229} : s = 71;
	{8'd167,8'd230} : s = 182;
	{8'd167,8'd231} : s = 181;
	{8'd167,8'd232} : s = 335;
	{8'd167,8'd233} : s = 13;
	{8'd167,8'd234} : s = 60;
	{8'd167,8'd235} : s = 58;
	{8'd167,8'd236} : s = 179;
	{8'd167,8'd237} : s = 57;
	{8'd167,8'd238} : s = 174;
	{8'd167,8'd239} : s = 173;
	{8'd167,8'd240} : s = 318;
	{8'd167,8'd241} : s = 54;
	{8'd167,8'd242} : s = 171;
	{8'd167,8'd243} : s = 167;
	{8'd167,8'd244} : s = 317;
	{8'd167,8'd245} : s = 158;
	{8'd167,8'd246} : s = 315;
	{8'd167,8'd247} : s = 311;
	{8'd167,8'd248} : s = 446;
	{8'd167,8'd249} : s = 11;
	{8'd167,8'd250} : s = 53;
	{8'd167,8'd251} : s = 51;
	{8'd167,8'd252} : s = 157;
	{8'd167,8'd253} : s = 46;
	{8'd167,8'd254} : s = 155;
	{8'd167,8'd255} : s = 151;
	{8'd168,8'd0} : s = 131;
	{8'd168,8'd1} : s = 281;
	{8'd168,8'd2} : s = 278;
	{8'd168,8'd3} : s = 409;
	{8'd168,8'd4} : s = 277;
	{8'd168,8'd5} : s = 406;
	{8'd168,8'd6} : s = 405;
	{8'd168,8'd7} : s = 485;
	{8'd168,8'd8} : s = 112;
	{8'd168,8'd9} : s = 275;
	{8'd168,8'd10} : s = 270;
	{8'd168,8'd11} : s = 403;
	{8'd168,8'd12} : s = 269;
	{8'd168,8'd13} : s = 398;
	{8'd168,8'd14} : s = 397;
	{8'd168,8'd15} : s = 483;
	{8'd168,8'd16} : s = 267;
	{8'd168,8'd17} : s = 395;
	{8'd168,8'd18} : s = 391;
	{8'd168,8'd19} : s = 476;
	{8'd168,8'd20} : s = 376;
	{8'd168,8'd21} : s = 474;
	{8'd168,8'd22} : s = 473;
	{8'd168,8'd23} : s = 506;
	{8'd168,8'd24} : s = 20;
	{8'd168,8'd25} : s = 104;
	{8'd168,8'd26} : s = 100;
	{8'd168,8'd27} : s = 263;
	{8'd168,8'd28} : s = 98;
	{8'd168,8'd29} : s = 240;
	{8'd168,8'd30} : s = 232;
	{8'd168,8'd31} : s = 372;
	{8'd168,8'd32} : s = 97;
	{8'd168,8'd33} : s = 228;
	{8'd168,8'd34} : s = 226;
	{8'd168,8'd35} : s = 370;
	{8'd168,8'd36} : s = 225;
	{8'd168,8'd37} : s = 369;
	{8'd168,8'd38} : s = 364;
	{8'd168,8'd39} : s = 470;
	{8'd168,8'd40} : s = 88;
	{8'd168,8'd41} : s = 216;
	{8'd168,8'd42} : s = 212;
	{8'd168,8'd43} : s = 362;
	{8'd168,8'd44} : s = 210;
	{8'd168,8'd45} : s = 361;
	{8'd168,8'd46} : s = 358;
	{8'd168,8'd47} : s = 469;
	{8'd168,8'd48} : s = 209;
	{8'd168,8'd49} : s = 357;
	{8'd168,8'd50} : s = 355;
	{8'd168,8'd51} : s = 467;
	{8'd168,8'd52} : s = 348;
	{8'd168,8'd53} : s = 462;
	{8'd168,8'd54} : s = 461;
	{8'd168,8'd55} : s = 505;
	{8'd168,8'd56} : s = 84;
	{8'd168,8'd57} : s = 204;
	{8'd168,8'd58} : s = 202;
	{8'd168,8'd59} : s = 346;
	{8'd168,8'd60} : s = 201;
	{8'd168,8'd61} : s = 345;
	{8'd168,8'd62} : s = 342;
	{8'd168,8'd63} : s = 459;
	{8'd168,8'd64} : s = 198;
	{8'd168,8'd65} : s = 341;
	{8'd168,8'd66} : s = 339;
	{8'd168,8'd67} : s = 455;
	{8'd168,8'd68} : s = 334;
	{8'd168,8'd69} : s = 444;
	{8'd168,8'd70} : s = 442;
	{8'd168,8'd71} : s = 502;
	{8'd168,8'd72} : s = 197;
	{8'd168,8'd73} : s = 333;
	{8'd168,8'd74} : s = 331;
	{8'd168,8'd75} : s = 441;
	{8'd168,8'd76} : s = 327;
	{8'd168,8'd77} : s = 438;
	{8'd168,8'd78} : s = 437;
	{8'd168,8'd79} : s = 501;
	{8'd168,8'd80} : s = 316;
	{8'd168,8'd81} : s = 435;
	{8'd168,8'd82} : s = 430;
	{8'd168,8'd83} : s = 499;
	{8'd168,8'd84} : s = 429;
	{8'd168,8'd85} : s = 494;
	{8'd168,8'd86} : s = 493;
	{8'd168,8'd87} : s = 510;
	{8'd168,8'd88} : s = 1;
	{8'd168,8'd89} : s = 18;
	{8'd168,8'd90} : s = 17;
	{8'd168,8'd91} : s = 82;
	{8'd168,8'd92} : s = 12;
	{8'd168,8'd93} : s = 81;
	{8'd168,8'd94} : s = 76;
	{8'd168,8'd95} : s = 195;
	{8'd168,8'd96} : s = 10;
	{8'd168,8'd97} : s = 74;
	{8'd168,8'd98} : s = 73;
	{8'd168,8'd99} : s = 184;
	{8'd168,8'd100} : s = 70;
	{8'd168,8'd101} : s = 180;
	{8'd168,8'd102} : s = 178;
	{8'd168,8'd103} : s = 314;
	{8'd168,8'd104} : s = 9;
	{8'd168,8'd105} : s = 69;
	{8'd168,8'd106} : s = 67;
	{8'd168,8'd107} : s = 177;
	{8'd168,8'd108} : s = 56;
	{8'd168,8'd109} : s = 172;
	{8'd168,8'd110} : s = 170;
	{8'd168,8'd111} : s = 313;
	{8'd168,8'd112} : s = 52;
	{8'd168,8'd113} : s = 169;
	{8'd168,8'd114} : s = 166;
	{8'd168,8'd115} : s = 310;
	{8'd168,8'd116} : s = 165;
	{8'd168,8'd117} : s = 309;
	{8'd168,8'd118} : s = 307;
	{8'd168,8'd119} : s = 427;
	{8'd168,8'd120} : s = 6;
	{8'd168,8'd121} : s = 50;
	{8'd168,8'd122} : s = 49;
	{8'd168,8'd123} : s = 163;
	{8'd168,8'd124} : s = 44;
	{8'd168,8'd125} : s = 156;
	{8'd168,8'd126} : s = 154;
	{8'd168,8'd127} : s = 302;
	{8'd168,8'd128} : s = 42;
	{8'd168,8'd129} : s = 153;
	{8'd168,8'd130} : s = 150;
	{8'd168,8'd131} : s = 301;
	{8'd168,8'd132} : s = 149;
	{8'd168,8'd133} : s = 299;
	{8'd168,8'd134} : s = 295;
	{8'd168,8'd135} : s = 423;
	{8'd168,8'd136} : s = 41;
	{8'd168,8'd137} : s = 147;
	{8'd168,8'd138} : s = 142;
	{8'd168,8'd139} : s = 286;
	{8'd168,8'd140} : s = 141;
	{8'd168,8'd141} : s = 285;
	{8'd168,8'd142} : s = 283;
	{8'd168,8'd143} : s = 414;
	{8'd168,8'd144} : s = 139;
	{8'd168,8'd145} : s = 279;
	{8'd168,8'd146} : s = 271;
	{8'd168,8'd147} : s = 413;
	{8'd168,8'd148} : s = 248;
	{8'd168,8'd149} : s = 411;
	{8'd168,8'd150} : s = 407;
	{8'd168,8'd151} : s = 491;
	{8'd168,8'd152} : s = 5;
	{8'd168,8'd153} : s = 38;
	{8'd168,8'd154} : s = 37;
	{8'd168,8'd155} : s = 135;
	{8'd168,8'd156} : s = 35;
	{8'd168,8'd157} : s = 120;
	{8'd168,8'd158} : s = 116;
	{8'd168,8'd159} : s = 244;
	{8'd168,8'd160} : s = 28;
	{8'd168,8'd161} : s = 114;
	{8'd168,8'd162} : s = 113;
	{8'd168,8'd163} : s = 242;
	{8'd168,8'd164} : s = 108;
	{8'd168,8'd165} : s = 241;
	{8'd168,8'd166} : s = 236;
	{8'd168,8'd167} : s = 399;
	{8'd168,8'd168} : s = 26;
	{8'd168,8'd169} : s = 106;
	{8'd168,8'd170} : s = 105;
	{8'd168,8'd171} : s = 234;
	{8'd168,8'd172} : s = 102;
	{8'd168,8'd173} : s = 233;
	{8'd168,8'd174} : s = 230;
	{8'd168,8'd175} : s = 380;
	{8'd168,8'd176} : s = 101;
	{8'd168,8'd177} : s = 229;
	{8'd168,8'd178} : s = 227;
	{8'd168,8'd179} : s = 378;
	{8'd168,8'd180} : s = 220;
	{8'd168,8'd181} : s = 377;
	{8'd168,8'd182} : s = 374;
	{8'd168,8'd183} : s = 487;
	{8'd168,8'd184} : s = 25;
	{8'd168,8'd185} : s = 99;
	{8'd168,8'd186} : s = 92;
	{8'd168,8'd187} : s = 218;
	{8'd168,8'd188} : s = 90;
	{8'd168,8'd189} : s = 217;
	{8'd168,8'd190} : s = 214;
	{8'd168,8'd191} : s = 373;
	{8'd168,8'd192} : s = 89;
	{8'd168,8'd193} : s = 213;
	{8'd168,8'd194} : s = 211;
	{8'd168,8'd195} : s = 371;
	{8'd168,8'd196} : s = 206;
	{8'd168,8'd197} : s = 366;
	{8'd168,8'd198} : s = 365;
	{8'd168,8'd199} : s = 478;
	{8'd168,8'd200} : s = 86;
	{8'd168,8'd201} : s = 205;
	{8'd168,8'd202} : s = 203;
	{8'd168,8'd203} : s = 363;
	{8'd168,8'd204} : s = 199;
	{8'd168,8'd205} : s = 359;
	{8'd168,8'd206} : s = 350;
	{8'd168,8'd207} : s = 477;
	{8'd168,8'd208} : s = 188;
	{8'd168,8'd209} : s = 349;
	{8'd168,8'd210} : s = 347;
	{8'd168,8'd211} : s = 475;
	{8'd168,8'd212} : s = 343;
	{8'd168,8'd213} : s = 471;
	{8'd168,8'd214} : s = 463;
	{8'd168,8'd215} : s = 509;
	{8'd168,8'd216} : s = 3;
	{8'd168,8'd217} : s = 22;
	{8'd168,8'd218} : s = 21;
	{8'd168,8'd219} : s = 85;
	{8'd168,8'd220} : s = 19;
	{8'd168,8'd221} : s = 83;
	{8'd168,8'd222} : s = 78;
	{8'd168,8'd223} : s = 186;
	{8'd168,8'd224} : s = 14;
	{8'd168,8'd225} : s = 77;
	{8'd168,8'd226} : s = 75;
	{8'd168,8'd227} : s = 185;
	{8'd168,8'd228} : s = 71;
	{8'd168,8'd229} : s = 182;
	{8'd168,8'd230} : s = 181;
	{8'd168,8'd231} : s = 335;
	{8'd168,8'd232} : s = 13;
	{8'd168,8'd233} : s = 60;
	{8'd168,8'd234} : s = 58;
	{8'd168,8'd235} : s = 179;
	{8'd168,8'd236} : s = 57;
	{8'd168,8'd237} : s = 174;
	{8'd168,8'd238} : s = 173;
	{8'd168,8'd239} : s = 318;
	{8'd168,8'd240} : s = 54;
	{8'd168,8'd241} : s = 171;
	{8'd168,8'd242} : s = 167;
	{8'd168,8'd243} : s = 317;
	{8'd168,8'd244} : s = 158;
	{8'd168,8'd245} : s = 315;
	{8'd168,8'd246} : s = 311;
	{8'd168,8'd247} : s = 446;
	{8'd168,8'd248} : s = 11;
	{8'd168,8'd249} : s = 53;
	{8'd168,8'd250} : s = 51;
	{8'd168,8'd251} : s = 157;
	{8'd168,8'd252} : s = 46;
	{8'd168,8'd253} : s = 155;
	{8'd168,8'd254} : s = 151;
	{8'd168,8'd255} : s = 303;
	{8'd169,8'd0} : s = 281;
	{8'd169,8'd1} : s = 278;
	{8'd169,8'd2} : s = 409;
	{8'd169,8'd3} : s = 277;
	{8'd169,8'd4} : s = 406;
	{8'd169,8'd5} : s = 405;
	{8'd169,8'd6} : s = 485;
	{8'd169,8'd7} : s = 112;
	{8'd169,8'd8} : s = 275;
	{8'd169,8'd9} : s = 270;
	{8'd169,8'd10} : s = 403;
	{8'd169,8'd11} : s = 269;
	{8'd169,8'd12} : s = 398;
	{8'd169,8'd13} : s = 397;
	{8'd169,8'd14} : s = 483;
	{8'd169,8'd15} : s = 267;
	{8'd169,8'd16} : s = 395;
	{8'd169,8'd17} : s = 391;
	{8'd169,8'd18} : s = 476;
	{8'd169,8'd19} : s = 376;
	{8'd169,8'd20} : s = 474;
	{8'd169,8'd21} : s = 473;
	{8'd169,8'd22} : s = 506;
	{8'd169,8'd23} : s = 20;
	{8'd169,8'd24} : s = 104;
	{8'd169,8'd25} : s = 100;
	{8'd169,8'd26} : s = 263;
	{8'd169,8'd27} : s = 98;
	{8'd169,8'd28} : s = 240;
	{8'd169,8'd29} : s = 232;
	{8'd169,8'd30} : s = 372;
	{8'd169,8'd31} : s = 97;
	{8'd169,8'd32} : s = 228;
	{8'd169,8'd33} : s = 226;
	{8'd169,8'd34} : s = 370;
	{8'd169,8'd35} : s = 225;
	{8'd169,8'd36} : s = 369;
	{8'd169,8'd37} : s = 364;
	{8'd169,8'd38} : s = 470;
	{8'd169,8'd39} : s = 88;
	{8'd169,8'd40} : s = 216;
	{8'd169,8'd41} : s = 212;
	{8'd169,8'd42} : s = 362;
	{8'd169,8'd43} : s = 210;
	{8'd169,8'd44} : s = 361;
	{8'd169,8'd45} : s = 358;
	{8'd169,8'd46} : s = 469;
	{8'd169,8'd47} : s = 209;
	{8'd169,8'd48} : s = 357;
	{8'd169,8'd49} : s = 355;
	{8'd169,8'd50} : s = 467;
	{8'd169,8'd51} : s = 348;
	{8'd169,8'd52} : s = 462;
	{8'd169,8'd53} : s = 461;
	{8'd169,8'd54} : s = 505;
	{8'd169,8'd55} : s = 84;
	{8'd169,8'd56} : s = 204;
	{8'd169,8'd57} : s = 202;
	{8'd169,8'd58} : s = 346;
	{8'd169,8'd59} : s = 201;
	{8'd169,8'd60} : s = 345;
	{8'd169,8'd61} : s = 342;
	{8'd169,8'd62} : s = 459;
	{8'd169,8'd63} : s = 198;
	{8'd169,8'd64} : s = 341;
	{8'd169,8'd65} : s = 339;
	{8'd169,8'd66} : s = 455;
	{8'd169,8'd67} : s = 334;
	{8'd169,8'd68} : s = 444;
	{8'd169,8'd69} : s = 442;
	{8'd169,8'd70} : s = 502;
	{8'd169,8'd71} : s = 197;
	{8'd169,8'd72} : s = 333;
	{8'd169,8'd73} : s = 331;
	{8'd169,8'd74} : s = 441;
	{8'd169,8'd75} : s = 327;
	{8'd169,8'd76} : s = 438;
	{8'd169,8'd77} : s = 437;
	{8'd169,8'd78} : s = 501;
	{8'd169,8'd79} : s = 316;
	{8'd169,8'd80} : s = 435;
	{8'd169,8'd81} : s = 430;
	{8'd169,8'd82} : s = 499;
	{8'd169,8'd83} : s = 429;
	{8'd169,8'd84} : s = 494;
	{8'd169,8'd85} : s = 493;
	{8'd169,8'd86} : s = 510;
	{8'd169,8'd87} : s = 1;
	{8'd169,8'd88} : s = 18;
	{8'd169,8'd89} : s = 17;
	{8'd169,8'd90} : s = 82;
	{8'd169,8'd91} : s = 12;
	{8'd169,8'd92} : s = 81;
	{8'd169,8'd93} : s = 76;
	{8'd169,8'd94} : s = 195;
	{8'd169,8'd95} : s = 10;
	{8'd169,8'd96} : s = 74;
	{8'd169,8'd97} : s = 73;
	{8'd169,8'd98} : s = 184;
	{8'd169,8'd99} : s = 70;
	{8'd169,8'd100} : s = 180;
	{8'd169,8'd101} : s = 178;
	{8'd169,8'd102} : s = 314;
	{8'd169,8'd103} : s = 9;
	{8'd169,8'd104} : s = 69;
	{8'd169,8'd105} : s = 67;
	{8'd169,8'd106} : s = 177;
	{8'd169,8'd107} : s = 56;
	{8'd169,8'd108} : s = 172;
	{8'd169,8'd109} : s = 170;
	{8'd169,8'd110} : s = 313;
	{8'd169,8'd111} : s = 52;
	{8'd169,8'd112} : s = 169;
	{8'd169,8'd113} : s = 166;
	{8'd169,8'd114} : s = 310;
	{8'd169,8'd115} : s = 165;
	{8'd169,8'd116} : s = 309;
	{8'd169,8'd117} : s = 307;
	{8'd169,8'd118} : s = 427;
	{8'd169,8'd119} : s = 6;
	{8'd169,8'd120} : s = 50;
	{8'd169,8'd121} : s = 49;
	{8'd169,8'd122} : s = 163;
	{8'd169,8'd123} : s = 44;
	{8'd169,8'd124} : s = 156;
	{8'd169,8'd125} : s = 154;
	{8'd169,8'd126} : s = 302;
	{8'd169,8'd127} : s = 42;
	{8'd169,8'd128} : s = 153;
	{8'd169,8'd129} : s = 150;
	{8'd169,8'd130} : s = 301;
	{8'd169,8'd131} : s = 149;
	{8'd169,8'd132} : s = 299;
	{8'd169,8'd133} : s = 295;
	{8'd169,8'd134} : s = 423;
	{8'd169,8'd135} : s = 41;
	{8'd169,8'd136} : s = 147;
	{8'd169,8'd137} : s = 142;
	{8'd169,8'd138} : s = 286;
	{8'd169,8'd139} : s = 141;
	{8'd169,8'd140} : s = 285;
	{8'd169,8'd141} : s = 283;
	{8'd169,8'd142} : s = 414;
	{8'd169,8'd143} : s = 139;
	{8'd169,8'd144} : s = 279;
	{8'd169,8'd145} : s = 271;
	{8'd169,8'd146} : s = 413;
	{8'd169,8'd147} : s = 248;
	{8'd169,8'd148} : s = 411;
	{8'd169,8'd149} : s = 407;
	{8'd169,8'd150} : s = 491;
	{8'd169,8'd151} : s = 5;
	{8'd169,8'd152} : s = 38;
	{8'd169,8'd153} : s = 37;
	{8'd169,8'd154} : s = 135;
	{8'd169,8'd155} : s = 35;
	{8'd169,8'd156} : s = 120;
	{8'd169,8'd157} : s = 116;
	{8'd169,8'd158} : s = 244;
	{8'd169,8'd159} : s = 28;
	{8'd169,8'd160} : s = 114;
	{8'd169,8'd161} : s = 113;
	{8'd169,8'd162} : s = 242;
	{8'd169,8'd163} : s = 108;
	{8'd169,8'd164} : s = 241;
	{8'd169,8'd165} : s = 236;
	{8'd169,8'd166} : s = 399;
	{8'd169,8'd167} : s = 26;
	{8'd169,8'd168} : s = 106;
	{8'd169,8'd169} : s = 105;
	{8'd169,8'd170} : s = 234;
	{8'd169,8'd171} : s = 102;
	{8'd169,8'd172} : s = 233;
	{8'd169,8'd173} : s = 230;
	{8'd169,8'd174} : s = 380;
	{8'd169,8'd175} : s = 101;
	{8'd169,8'd176} : s = 229;
	{8'd169,8'd177} : s = 227;
	{8'd169,8'd178} : s = 378;
	{8'd169,8'd179} : s = 220;
	{8'd169,8'd180} : s = 377;
	{8'd169,8'd181} : s = 374;
	{8'd169,8'd182} : s = 487;
	{8'd169,8'd183} : s = 25;
	{8'd169,8'd184} : s = 99;
	{8'd169,8'd185} : s = 92;
	{8'd169,8'd186} : s = 218;
	{8'd169,8'd187} : s = 90;
	{8'd169,8'd188} : s = 217;
	{8'd169,8'd189} : s = 214;
	{8'd169,8'd190} : s = 373;
	{8'd169,8'd191} : s = 89;
	{8'd169,8'd192} : s = 213;
	{8'd169,8'd193} : s = 211;
	{8'd169,8'd194} : s = 371;
	{8'd169,8'd195} : s = 206;
	{8'd169,8'd196} : s = 366;
	{8'd169,8'd197} : s = 365;
	{8'd169,8'd198} : s = 478;
	{8'd169,8'd199} : s = 86;
	{8'd169,8'd200} : s = 205;
	{8'd169,8'd201} : s = 203;
	{8'd169,8'd202} : s = 363;
	{8'd169,8'd203} : s = 199;
	{8'd169,8'd204} : s = 359;
	{8'd169,8'd205} : s = 350;
	{8'd169,8'd206} : s = 477;
	{8'd169,8'd207} : s = 188;
	{8'd169,8'd208} : s = 349;
	{8'd169,8'd209} : s = 347;
	{8'd169,8'd210} : s = 475;
	{8'd169,8'd211} : s = 343;
	{8'd169,8'd212} : s = 471;
	{8'd169,8'd213} : s = 463;
	{8'd169,8'd214} : s = 509;
	{8'd169,8'd215} : s = 3;
	{8'd169,8'd216} : s = 22;
	{8'd169,8'd217} : s = 21;
	{8'd169,8'd218} : s = 85;
	{8'd169,8'd219} : s = 19;
	{8'd169,8'd220} : s = 83;
	{8'd169,8'd221} : s = 78;
	{8'd169,8'd222} : s = 186;
	{8'd169,8'd223} : s = 14;
	{8'd169,8'd224} : s = 77;
	{8'd169,8'd225} : s = 75;
	{8'd169,8'd226} : s = 185;
	{8'd169,8'd227} : s = 71;
	{8'd169,8'd228} : s = 182;
	{8'd169,8'd229} : s = 181;
	{8'd169,8'd230} : s = 335;
	{8'd169,8'd231} : s = 13;
	{8'd169,8'd232} : s = 60;
	{8'd169,8'd233} : s = 58;
	{8'd169,8'd234} : s = 179;
	{8'd169,8'd235} : s = 57;
	{8'd169,8'd236} : s = 174;
	{8'd169,8'd237} : s = 173;
	{8'd169,8'd238} : s = 318;
	{8'd169,8'd239} : s = 54;
	{8'd169,8'd240} : s = 171;
	{8'd169,8'd241} : s = 167;
	{8'd169,8'd242} : s = 317;
	{8'd169,8'd243} : s = 158;
	{8'd169,8'd244} : s = 315;
	{8'd169,8'd245} : s = 311;
	{8'd169,8'd246} : s = 446;
	{8'd169,8'd247} : s = 11;
	{8'd169,8'd248} : s = 53;
	{8'd169,8'd249} : s = 51;
	{8'd169,8'd250} : s = 157;
	{8'd169,8'd251} : s = 46;
	{8'd169,8'd252} : s = 155;
	{8'd169,8'd253} : s = 151;
	{8'd169,8'd254} : s = 303;
	{8'd169,8'd255} : s = 45;
	{8'd170,8'd0} : s = 278;
	{8'd170,8'd1} : s = 409;
	{8'd170,8'd2} : s = 277;
	{8'd170,8'd3} : s = 406;
	{8'd170,8'd4} : s = 405;
	{8'd170,8'd5} : s = 485;
	{8'd170,8'd6} : s = 112;
	{8'd170,8'd7} : s = 275;
	{8'd170,8'd8} : s = 270;
	{8'd170,8'd9} : s = 403;
	{8'd170,8'd10} : s = 269;
	{8'd170,8'd11} : s = 398;
	{8'd170,8'd12} : s = 397;
	{8'd170,8'd13} : s = 483;
	{8'd170,8'd14} : s = 267;
	{8'd170,8'd15} : s = 395;
	{8'd170,8'd16} : s = 391;
	{8'd170,8'd17} : s = 476;
	{8'd170,8'd18} : s = 376;
	{8'd170,8'd19} : s = 474;
	{8'd170,8'd20} : s = 473;
	{8'd170,8'd21} : s = 506;
	{8'd170,8'd22} : s = 20;
	{8'd170,8'd23} : s = 104;
	{8'd170,8'd24} : s = 100;
	{8'd170,8'd25} : s = 263;
	{8'd170,8'd26} : s = 98;
	{8'd170,8'd27} : s = 240;
	{8'd170,8'd28} : s = 232;
	{8'd170,8'd29} : s = 372;
	{8'd170,8'd30} : s = 97;
	{8'd170,8'd31} : s = 228;
	{8'd170,8'd32} : s = 226;
	{8'd170,8'd33} : s = 370;
	{8'd170,8'd34} : s = 225;
	{8'd170,8'd35} : s = 369;
	{8'd170,8'd36} : s = 364;
	{8'd170,8'd37} : s = 470;
	{8'd170,8'd38} : s = 88;
	{8'd170,8'd39} : s = 216;
	{8'd170,8'd40} : s = 212;
	{8'd170,8'd41} : s = 362;
	{8'd170,8'd42} : s = 210;
	{8'd170,8'd43} : s = 361;
	{8'd170,8'd44} : s = 358;
	{8'd170,8'd45} : s = 469;
	{8'd170,8'd46} : s = 209;
	{8'd170,8'd47} : s = 357;
	{8'd170,8'd48} : s = 355;
	{8'd170,8'd49} : s = 467;
	{8'd170,8'd50} : s = 348;
	{8'd170,8'd51} : s = 462;
	{8'd170,8'd52} : s = 461;
	{8'd170,8'd53} : s = 505;
	{8'd170,8'd54} : s = 84;
	{8'd170,8'd55} : s = 204;
	{8'd170,8'd56} : s = 202;
	{8'd170,8'd57} : s = 346;
	{8'd170,8'd58} : s = 201;
	{8'd170,8'd59} : s = 345;
	{8'd170,8'd60} : s = 342;
	{8'd170,8'd61} : s = 459;
	{8'd170,8'd62} : s = 198;
	{8'd170,8'd63} : s = 341;
	{8'd170,8'd64} : s = 339;
	{8'd170,8'd65} : s = 455;
	{8'd170,8'd66} : s = 334;
	{8'd170,8'd67} : s = 444;
	{8'd170,8'd68} : s = 442;
	{8'd170,8'd69} : s = 502;
	{8'd170,8'd70} : s = 197;
	{8'd170,8'd71} : s = 333;
	{8'd170,8'd72} : s = 331;
	{8'd170,8'd73} : s = 441;
	{8'd170,8'd74} : s = 327;
	{8'd170,8'd75} : s = 438;
	{8'd170,8'd76} : s = 437;
	{8'd170,8'd77} : s = 501;
	{8'd170,8'd78} : s = 316;
	{8'd170,8'd79} : s = 435;
	{8'd170,8'd80} : s = 430;
	{8'd170,8'd81} : s = 499;
	{8'd170,8'd82} : s = 429;
	{8'd170,8'd83} : s = 494;
	{8'd170,8'd84} : s = 493;
	{8'd170,8'd85} : s = 510;
	{8'd170,8'd86} : s = 1;
	{8'd170,8'd87} : s = 18;
	{8'd170,8'd88} : s = 17;
	{8'd170,8'd89} : s = 82;
	{8'd170,8'd90} : s = 12;
	{8'd170,8'd91} : s = 81;
	{8'd170,8'd92} : s = 76;
	{8'd170,8'd93} : s = 195;
	{8'd170,8'd94} : s = 10;
	{8'd170,8'd95} : s = 74;
	{8'd170,8'd96} : s = 73;
	{8'd170,8'd97} : s = 184;
	{8'd170,8'd98} : s = 70;
	{8'd170,8'd99} : s = 180;
	{8'd170,8'd100} : s = 178;
	{8'd170,8'd101} : s = 314;
	{8'd170,8'd102} : s = 9;
	{8'd170,8'd103} : s = 69;
	{8'd170,8'd104} : s = 67;
	{8'd170,8'd105} : s = 177;
	{8'd170,8'd106} : s = 56;
	{8'd170,8'd107} : s = 172;
	{8'd170,8'd108} : s = 170;
	{8'd170,8'd109} : s = 313;
	{8'd170,8'd110} : s = 52;
	{8'd170,8'd111} : s = 169;
	{8'd170,8'd112} : s = 166;
	{8'd170,8'd113} : s = 310;
	{8'd170,8'd114} : s = 165;
	{8'd170,8'd115} : s = 309;
	{8'd170,8'd116} : s = 307;
	{8'd170,8'd117} : s = 427;
	{8'd170,8'd118} : s = 6;
	{8'd170,8'd119} : s = 50;
	{8'd170,8'd120} : s = 49;
	{8'd170,8'd121} : s = 163;
	{8'd170,8'd122} : s = 44;
	{8'd170,8'd123} : s = 156;
	{8'd170,8'd124} : s = 154;
	{8'd170,8'd125} : s = 302;
	{8'd170,8'd126} : s = 42;
	{8'd170,8'd127} : s = 153;
	{8'd170,8'd128} : s = 150;
	{8'd170,8'd129} : s = 301;
	{8'd170,8'd130} : s = 149;
	{8'd170,8'd131} : s = 299;
	{8'd170,8'd132} : s = 295;
	{8'd170,8'd133} : s = 423;
	{8'd170,8'd134} : s = 41;
	{8'd170,8'd135} : s = 147;
	{8'd170,8'd136} : s = 142;
	{8'd170,8'd137} : s = 286;
	{8'd170,8'd138} : s = 141;
	{8'd170,8'd139} : s = 285;
	{8'd170,8'd140} : s = 283;
	{8'd170,8'd141} : s = 414;
	{8'd170,8'd142} : s = 139;
	{8'd170,8'd143} : s = 279;
	{8'd170,8'd144} : s = 271;
	{8'd170,8'd145} : s = 413;
	{8'd170,8'd146} : s = 248;
	{8'd170,8'd147} : s = 411;
	{8'd170,8'd148} : s = 407;
	{8'd170,8'd149} : s = 491;
	{8'd170,8'd150} : s = 5;
	{8'd170,8'd151} : s = 38;
	{8'd170,8'd152} : s = 37;
	{8'd170,8'd153} : s = 135;
	{8'd170,8'd154} : s = 35;
	{8'd170,8'd155} : s = 120;
	{8'd170,8'd156} : s = 116;
	{8'd170,8'd157} : s = 244;
	{8'd170,8'd158} : s = 28;
	{8'd170,8'd159} : s = 114;
	{8'd170,8'd160} : s = 113;
	{8'd170,8'd161} : s = 242;
	{8'd170,8'd162} : s = 108;
	{8'd170,8'd163} : s = 241;
	{8'd170,8'd164} : s = 236;
	{8'd170,8'd165} : s = 399;
	{8'd170,8'd166} : s = 26;
	{8'd170,8'd167} : s = 106;
	{8'd170,8'd168} : s = 105;
	{8'd170,8'd169} : s = 234;
	{8'd170,8'd170} : s = 102;
	{8'd170,8'd171} : s = 233;
	{8'd170,8'd172} : s = 230;
	{8'd170,8'd173} : s = 380;
	{8'd170,8'd174} : s = 101;
	{8'd170,8'd175} : s = 229;
	{8'd170,8'd176} : s = 227;
	{8'd170,8'd177} : s = 378;
	{8'd170,8'd178} : s = 220;
	{8'd170,8'd179} : s = 377;
	{8'd170,8'd180} : s = 374;
	{8'd170,8'd181} : s = 487;
	{8'd170,8'd182} : s = 25;
	{8'd170,8'd183} : s = 99;
	{8'd170,8'd184} : s = 92;
	{8'd170,8'd185} : s = 218;
	{8'd170,8'd186} : s = 90;
	{8'd170,8'd187} : s = 217;
	{8'd170,8'd188} : s = 214;
	{8'd170,8'd189} : s = 373;
	{8'd170,8'd190} : s = 89;
	{8'd170,8'd191} : s = 213;
	{8'd170,8'd192} : s = 211;
	{8'd170,8'd193} : s = 371;
	{8'd170,8'd194} : s = 206;
	{8'd170,8'd195} : s = 366;
	{8'd170,8'd196} : s = 365;
	{8'd170,8'd197} : s = 478;
	{8'd170,8'd198} : s = 86;
	{8'd170,8'd199} : s = 205;
	{8'd170,8'd200} : s = 203;
	{8'd170,8'd201} : s = 363;
	{8'd170,8'd202} : s = 199;
	{8'd170,8'd203} : s = 359;
	{8'd170,8'd204} : s = 350;
	{8'd170,8'd205} : s = 477;
	{8'd170,8'd206} : s = 188;
	{8'd170,8'd207} : s = 349;
	{8'd170,8'd208} : s = 347;
	{8'd170,8'd209} : s = 475;
	{8'd170,8'd210} : s = 343;
	{8'd170,8'd211} : s = 471;
	{8'd170,8'd212} : s = 463;
	{8'd170,8'd213} : s = 509;
	{8'd170,8'd214} : s = 3;
	{8'd170,8'd215} : s = 22;
	{8'd170,8'd216} : s = 21;
	{8'd170,8'd217} : s = 85;
	{8'd170,8'd218} : s = 19;
	{8'd170,8'd219} : s = 83;
	{8'd170,8'd220} : s = 78;
	{8'd170,8'd221} : s = 186;
	{8'd170,8'd222} : s = 14;
	{8'd170,8'd223} : s = 77;
	{8'd170,8'd224} : s = 75;
	{8'd170,8'd225} : s = 185;
	{8'd170,8'd226} : s = 71;
	{8'd170,8'd227} : s = 182;
	{8'd170,8'd228} : s = 181;
	{8'd170,8'd229} : s = 335;
	{8'd170,8'd230} : s = 13;
	{8'd170,8'd231} : s = 60;
	{8'd170,8'd232} : s = 58;
	{8'd170,8'd233} : s = 179;
	{8'd170,8'd234} : s = 57;
	{8'd170,8'd235} : s = 174;
	{8'd170,8'd236} : s = 173;
	{8'd170,8'd237} : s = 318;
	{8'd170,8'd238} : s = 54;
	{8'd170,8'd239} : s = 171;
	{8'd170,8'd240} : s = 167;
	{8'd170,8'd241} : s = 317;
	{8'd170,8'd242} : s = 158;
	{8'd170,8'd243} : s = 315;
	{8'd170,8'd244} : s = 311;
	{8'd170,8'd245} : s = 446;
	{8'd170,8'd246} : s = 11;
	{8'd170,8'd247} : s = 53;
	{8'd170,8'd248} : s = 51;
	{8'd170,8'd249} : s = 157;
	{8'd170,8'd250} : s = 46;
	{8'd170,8'd251} : s = 155;
	{8'd170,8'd252} : s = 151;
	{8'd170,8'd253} : s = 303;
	{8'd170,8'd254} : s = 45;
	{8'd170,8'd255} : s = 143;
	{8'd171,8'd0} : s = 409;
	{8'd171,8'd1} : s = 277;
	{8'd171,8'd2} : s = 406;
	{8'd171,8'd3} : s = 405;
	{8'd171,8'd4} : s = 485;
	{8'd171,8'd5} : s = 112;
	{8'd171,8'd6} : s = 275;
	{8'd171,8'd7} : s = 270;
	{8'd171,8'd8} : s = 403;
	{8'd171,8'd9} : s = 269;
	{8'd171,8'd10} : s = 398;
	{8'd171,8'd11} : s = 397;
	{8'd171,8'd12} : s = 483;
	{8'd171,8'd13} : s = 267;
	{8'd171,8'd14} : s = 395;
	{8'd171,8'd15} : s = 391;
	{8'd171,8'd16} : s = 476;
	{8'd171,8'd17} : s = 376;
	{8'd171,8'd18} : s = 474;
	{8'd171,8'd19} : s = 473;
	{8'd171,8'd20} : s = 506;
	{8'd171,8'd21} : s = 20;
	{8'd171,8'd22} : s = 104;
	{8'd171,8'd23} : s = 100;
	{8'd171,8'd24} : s = 263;
	{8'd171,8'd25} : s = 98;
	{8'd171,8'd26} : s = 240;
	{8'd171,8'd27} : s = 232;
	{8'd171,8'd28} : s = 372;
	{8'd171,8'd29} : s = 97;
	{8'd171,8'd30} : s = 228;
	{8'd171,8'd31} : s = 226;
	{8'd171,8'd32} : s = 370;
	{8'd171,8'd33} : s = 225;
	{8'd171,8'd34} : s = 369;
	{8'd171,8'd35} : s = 364;
	{8'd171,8'd36} : s = 470;
	{8'd171,8'd37} : s = 88;
	{8'd171,8'd38} : s = 216;
	{8'd171,8'd39} : s = 212;
	{8'd171,8'd40} : s = 362;
	{8'd171,8'd41} : s = 210;
	{8'd171,8'd42} : s = 361;
	{8'd171,8'd43} : s = 358;
	{8'd171,8'd44} : s = 469;
	{8'd171,8'd45} : s = 209;
	{8'd171,8'd46} : s = 357;
	{8'd171,8'd47} : s = 355;
	{8'd171,8'd48} : s = 467;
	{8'd171,8'd49} : s = 348;
	{8'd171,8'd50} : s = 462;
	{8'd171,8'd51} : s = 461;
	{8'd171,8'd52} : s = 505;
	{8'd171,8'd53} : s = 84;
	{8'd171,8'd54} : s = 204;
	{8'd171,8'd55} : s = 202;
	{8'd171,8'd56} : s = 346;
	{8'd171,8'd57} : s = 201;
	{8'd171,8'd58} : s = 345;
	{8'd171,8'd59} : s = 342;
	{8'd171,8'd60} : s = 459;
	{8'd171,8'd61} : s = 198;
	{8'd171,8'd62} : s = 341;
	{8'd171,8'd63} : s = 339;
	{8'd171,8'd64} : s = 455;
	{8'd171,8'd65} : s = 334;
	{8'd171,8'd66} : s = 444;
	{8'd171,8'd67} : s = 442;
	{8'd171,8'd68} : s = 502;
	{8'd171,8'd69} : s = 197;
	{8'd171,8'd70} : s = 333;
	{8'd171,8'd71} : s = 331;
	{8'd171,8'd72} : s = 441;
	{8'd171,8'd73} : s = 327;
	{8'd171,8'd74} : s = 438;
	{8'd171,8'd75} : s = 437;
	{8'd171,8'd76} : s = 501;
	{8'd171,8'd77} : s = 316;
	{8'd171,8'd78} : s = 435;
	{8'd171,8'd79} : s = 430;
	{8'd171,8'd80} : s = 499;
	{8'd171,8'd81} : s = 429;
	{8'd171,8'd82} : s = 494;
	{8'd171,8'd83} : s = 493;
	{8'd171,8'd84} : s = 510;
	{8'd171,8'd85} : s = 1;
	{8'd171,8'd86} : s = 18;
	{8'd171,8'd87} : s = 17;
	{8'd171,8'd88} : s = 82;
	{8'd171,8'd89} : s = 12;
	{8'd171,8'd90} : s = 81;
	{8'd171,8'd91} : s = 76;
	{8'd171,8'd92} : s = 195;
	{8'd171,8'd93} : s = 10;
	{8'd171,8'd94} : s = 74;
	{8'd171,8'd95} : s = 73;
	{8'd171,8'd96} : s = 184;
	{8'd171,8'd97} : s = 70;
	{8'd171,8'd98} : s = 180;
	{8'd171,8'd99} : s = 178;
	{8'd171,8'd100} : s = 314;
	{8'd171,8'd101} : s = 9;
	{8'd171,8'd102} : s = 69;
	{8'd171,8'd103} : s = 67;
	{8'd171,8'd104} : s = 177;
	{8'd171,8'd105} : s = 56;
	{8'd171,8'd106} : s = 172;
	{8'd171,8'd107} : s = 170;
	{8'd171,8'd108} : s = 313;
	{8'd171,8'd109} : s = 52;
	{8'd171,8'd110} : s = 169;
	{8'd171,8'd111} : s = 166;
	{8'd171,8'd112} : s = 310;
	{8'd171,8'd113} : s = 165;
	{8'd171,8'd114} : s = 309;
	{8'd171,8'd115} : s = 307;
	{8'd171,8'd116} : s = 427;
	{8'd171,8'd117} : s = 6;
	{8'd171,8'd118} : s = 50;
	{8'd171,8'd119} : s = 49;
	{8'd171,8'd120} : s = 163;
	{8'd171,8'd121} : s = 44;
	{8'd171,8'd122} : s = 156;
	{8'd171,8'd123} : s = 154;
	{8'd171,8'd124} : s = 302;
	{8'd171,8'd125} : s = 42;
	{8'd171,8'd126} : s = 153;
	{8'd171,8'd127} : s = 150;
	{8'd171,8'd128} : s = 301;
	{8'd171,8'd129} : s = 149;
	{8'd171,8'd130} : s = 299;
	{8'd171,8'd131} : s = 295;
	{8'd171,8'd132} : s = 423;
	{8'd171,8'd133} : s = 41;
	{8'd171,8'd134} : s = 147;
	{8'd171,8'd135} : s = 142;
	{8'd171,8'd136} : s = 286;
	{8'd171,8'd137} : s = 141;
	{8'd171,8'd138} : s = 285;
	{8'd171,8'd139} : s = 283;
	{8'd171,8'd140} : s = 414;
	{8'd171,8'd141} : s = 139;
	{8'd171,8'd142} : s = 279;
	{8'd171,8'd143} : s = 271;
	{8'd171,8'd144} : s = 413;
	{8'd171,8'd145} : s = 248;
	{8'd171,8'd146} : s = 411;
	{8'd171,8'd147} : s = 407;
	{8'd171,8'd148} : s = 491;
	{8'd171,8'd149} : s = 5;
	{8'd171,8'd150} : s = 38;
	{8'd171,8'd151} : s = 37;
	{8'd171,8'd152} : s = 135;
	{8'd171,8'd153} : s = 35;
	{8'd171,8'd154} : s = 120;
	{8'd171,8'd155} : s = 116;
	{8'd171,8'd156} : s = 244;
	{8'd171,8'd157} : s = 28;
	{8'd171,8'd158} : s = 114;
	{8'd171,8'd159} : s = 113;
	{8'd171,8'd160} : s = 242;
	{8'd171,8'd161} : s = 108;
	{8'd171,8'd162} : s = 241;
	{8'd171,8'd163} : s = 236;
	{8'd171,8'd164} : s = 399;
	{8'd171,8'd165} : s = 26;
	{8'd171,8'd166} : s = 106;
	{8'd171,8'd167} : s = 105;
	{8'd171,8'd168} : s = 234;
	{8'd171,8'd169} : s = 102;
	{8'd171,8'd170} : s = 233;
	{8'd171,8'd171} : s = 230;
	{8'd171,8'd172} : s = 380;
	{8'd171,8'd173} : s = 101;
	{8'd171,8'd174} : s = 229;
	{8'd171,8'd175} : s = 227;
	{8'd171,8'd176} : s = 378;
	{8'd171,8'd177} : s = 220;
	{8'd171,8'd178} : s = 377;
	{8'd171,8'd179} : s = 374;
	{8'd171,8'd180} : s = 487;
	{8'd171,8'd181} : s = 25;
	{8'd171,8'd182} : s = 99;
	{8'd171,8'd183} : s = 92;
	{8'd171,8'd184} : s = 218;
	{8'd171,8'd185} : s = 90;
	{8'd171,8'd186} : s = 217;
	{8'd171,8'd187} : s = 214;
	{8'd171,8'd188} : s = 373;
	{8'd171,8'd189} : s = 89;
	{8'd171,8'd190} : s = 213;
	{8'd171,8'd191} : s = 211;
	{8'd171,8'd192} : s = 371;
	{8'd171,8'd193} : s = 206;
	{8'd171,8'd194} : s = 366;
	{8'd171,8'd195} : s = 365;
	{8'd171,8'd196} : s = 478;
	{8'd171,8'd197} : s = 86;
	{8'd171,8'd198} : s = 205;
	{8'd171,8'd199} : s = 203;
	{8'd171,8'd200} : s = 363;
	{8'd171,8'd201} : s = 199;
	{8'd171,8'd202} : s = 359;
	{8'd171,8'd203} : s = 350;
	{8'd171,8'd204} : s = 477;
	{8'd171,8'd205} : s = 188;
	{8'd171,8'd206} : s = 349;
	{8'd171,8'd207} : s = 347;
	{8'd171,8'd208} : s = 475;
	{8'd171,8'd209} : s = 343;
	{8'd171,8'd210} : s = 471;
	{8'd171,8'd211} : s = 463;
	{8'd171,8'd212} : s = 509;
	{8'd171,8'd213} : s = 3;
	{8'd171,8'd214} : s = 22;
	{8'd171,8'd215} : s = 21;
	{8'd171,8'd216} : s = 85;
	{8'd171,8'd217} : s = 19;
	{8'd171,8'd218} : s = 83;
	{8'd171,8'd219} : s = 78;
	{8'd171,8'd220} : s = 186;
	{8'd171,8'd221} : s = 14;
	{8'd171,8'd222} : s = 77;
	{8'd171,8'd223} : s = 75;
	{8'd171,8'd224} : s = 185;
	{8'd171,8'd225} : s = 71;
	{8'd171,8'd226} : s = 182;
	{8'd171,8'd227} : s = 181;
	{8'd171,8'd228} : s = 335;
	{8'd171,8'd229} : s = 13;
	{8'd171,8'd230} : s = 60;
	{8'd171,8'd231} : s = 58;
	{8'd171,8'd232} : s = 179;
	{8'd171,8'd233} : s = 57;
	{8'd171,8'd234} : s = 174;
	{8'd171,8'd235} : s = 173;
	{8'd171,8'd236} : s = 318;
	{8'd171,8'd237} : s = 54;
	{8'd171,8'd238} : s = 171;
	{8'd171,8'd239} : s = 167;
	{8'd171,8'd240} : s = 317;
	{8'd171,8'd241} : s = 158;
	{8'd171,8'd242} : s = 315;
	{8'd171,8'd243} : s = 311;
	{8'd171,8'd244} : s = 446;
	{8'd171,8'd245} : s = 11;
	{8'd171,8'd246} : s = 53;
	{8'd171,8'd247} : s = 51;
	{8'd171,8'd248} : s = 157;
	{8'd171,8'd249} : s = 46;
	{8'd171,8'd250} : s = 155;
	{8'd171,8'd251} : s = 151;
	{8'd171,8'd252} : s = 303;
	{8'd171,8'd253} : s = 45;
	{8'd171,8'd254} : s = 143;
	{8'd171,8'd255} : s = 124;
	{8'd172,8'd0} : s = 277;
	{8'd172,8'd1} : s = 406;
	{8'd172,8'd2} : s = 405;
	{8'd172,8'd3} : s = 485;
	{8'd172,8'd4} : s = 112;
	{8'd172,8'd5} : s = 275;
	{8'd172,8'd6} : s = 270;
	{8'd172,8'd7} : s = 403;
	{8'd172,8'd8} : s = 269;
	{8'd172,8'd9} : s = 398;
	{8'd172,8'd10} : s = 397;
	{8'd172,8'd11} : s = 483;
	{8'd172,8'd12} : s = 267;
	{8'd172,8'd13} : s = 395;
	{8'd172,8'd14} : s = 391;
	{8'd172,8'd15} : s = 476;
	{8'd172,8'd16} : s = 376;
	{8'd172,8'd17} : s = 474;
	{8'd172,8'd18} : s = 473;
	{8'd172,8'd19} : s = 506;
	{8'd172,8'd20} : s = 20;
	{8'd172,8'd21} : s = 104;
	{8'd172,8'd22} : s = 100;
	{8'd172,8'd23} : s = 263;
	{8'd172,8'd24} : s = 98;
	{8'd172,8'd25} : s = 240;
	{8'd172,8'd26} : s = 232;
	{8'd172,8'd27} : s = 372;
	{8'd172,8'd28} : s = 97;
	{8'd172,8'd29} : s = 228;
	{8'd172,8'd30} : s = 226;
	{8'd172,8'd31} : s = 370;
	{8'd172,8'd32} : s = 225;
	{8'd172,8'd33} : s = 369;
	{8'd172,8'd34} : s = 364;
	{8'd172,8'd35} : s = 470;
	{8'd172,8'd36} : s = 88;
	{8'd172,8'd37} : s = 216;
	{8'd172,8'd38} : s = 212;
	{8'd172,8'd39} : s = 362;
	{8'd172,8'd40} : s = 210;
	{8'd172,8'd41} : s = 361;
	{8'd172,8'd42} : s = 358;
	{8'd172,8'd43} : s = 469;
	{8'd172,8'd44} : s = 209;
	{8'd172,8'd45} : s = 357;
	{8'd172,8'd46} : s = 355;
	{8'd172,8'd47} : s = 467;
	{8'd172,8'd48} : s = 348;
	{8'd172,8'd49} : s = 462;
	{8'd172,8'd50} : s = 461;
	{8'd172,8'd51} : s = 505;
	{8'd172,8'd52} : s = 84;
	{8'd172,8'd53} : s = 204;
	{8'd172,8'd54} : s = 202;
	{8'd172,8'd55} : s = 346;
	{8'd172,8'd56} : s = 201;
	{8'd172,8'd57} : s = 345;
	{8'd172,8'd58} : s = 342;
	{8'd172,8'd59} : s = 459;
	{8'd172,8'd60} : s = 198;
	{8'd172,8'd61} : s = 341;
	{8'd172,8'd62} : s = 339;
	{8'd172,8'd63} : s = 455;
	{8'd172,8'd64} : s = 334;
	{8'd172,8'd65} : s = 444;
	{8'd172,8'd66} : s = 442;
	{8'd172,8'd67} : s = 502;
	{8'd172,8'd68} : s = 197;
	{8'd172,8'd69} : s = 333;
	{8'd172,8'd70} : s = 331;
	{8'd172,8'd71} : s = 441;
	{8'd172,8'd72} : s = 327;
	{8'd172,8'd73} : s = 438;
	{8'd172,8'd74} : s = 437;
	{8'd172,8'd75} : s = 501;
	{8'd172,8'd76} : s = 316;
	{8'd172,8'd77} : s = 435;
	{8'd172,8'd78} : s = 430;
	{8'd172,8'd79} : s = 499;
	{8'd172,8'd80} : s = 429;
	{8'd172,8'd81} : s = 494;
	{8'd172,8'd82} : s = 493;
	{8'd172,8'd83} : s = 510;
	{8'd172,8'd84} : s = 1;
	{8'd172,8'd85} : s = 18;
	{8'd172,8'd86} : s = 17;
	{8'd172,8'd87} : s = 82;
	{8'd172,8'd88} : s = 12;
	{8'd172,8'd89} : s = 81;
	{8'd172,8'd90} : s = 76;
	{8'd172,8'd91} : s = 195;
	{8'd172,8'd92} : s = 10;
	{8'd172,8'd93} : s = 74;
	{8'd172,8'd94} : s = 73;
	{8'd172,8'd95} : s = 184;
	{8'd172,8'd96} : s = 70;
	{8'd172,8'd97} : s = 180;
	{8'd172,8'd98} : s = 178;
	{8'd172,8'd99} : s = 314;
	{8'd172,8'd100} : s = 9;
	{8'd172,8'd101} : s = 69;
	{8'd172,8'd102} : s = 67;
	{8'd172,8'd103} : s = 177;
	{8'd172,8'd104} : s = 56;
	{8'd172,8'd105} : s = 172;
	{8'd172,8'd106} : s = 170;
	{8'd172,8'd107} : s = 313;
	{8'd172,8'd108} : s = 52;
	{8'd172,8'd109} : s = 169;
	{8'd172,8'd110} : s = 166;
	{8'd172,8'd111} : s = 310;
	{8'd172,8'd112} : s = 165;
	{8'd172,8'd113} : s = 309;
	{8'd172,8'd114} : s = 307;
	{8'd172,8'd115} : s = 427;
	{8'd172,8'd116} : s = 6;
	{8'd172,8'd117} : s = 50;
	{8'd172,8'd118} : s = 49;
	{8'd172,8'd119} : s = 163;
	{8'd172,8'd120} : s = 44;
	{8'd172,8'd121} : s = 156;
	{8'd172,8'd122} : s = 154;
	{8'd172,8'd123} : s = 302;
	{8'd172,8'd124} : s = 42;
	{8'd172,8'd125} : s = 153;
	{8'd172,8'd126} : s = 150;
	{8'd172,8'd127} : s = 301;
	{8'd172,8'd128} : s = 149;
	{8'd172,8'd129} : s = 299;
	{8'd172,8'd130} : s = 295;
	{8'd172,8'd131} : s = 423;
	{8'd172,8'd132} : s = 41;
	{8'd172,8'd133} : s = 147;
	{8'd172,8'd134} : s = 142;
	{8'd172,8'd135} : s = 286;
	{8'd172,8'd136} : s = 141;
	{8'd172,8'd137} : s = 285;
	{8'd172,8'd138} : s = 283;
	{8'd172,8'd139} : s = 414;
	{8'd172,8'd140} : s = 139;
	{8'd172,8'd141} : s = 279;
	{8'd172,8'd142} : s = 271;
	{8'd172,8'd143} : s = 413;
	{8'd172,8'd144} : s = 248;
	{8'd172,8'd145} : s = 411;
	{8'd172,8'd146} : s = 407;
	{8'd172,8'd147} : s = 491;
	{8'd172,8'd148} : s = 5;
	{8'd172,8'd149} : s = 38;
	{8'd172,8'd150} : s = 37;
	{8'd172,8'd151} : s = 135;
	{8'd172,8'd152} : s = 35;
	{8'd172,8'd153} : s = 120;
	{8'd172,8'd154} : s = 116;
	{8'd172,8'd155} : s = 244;
	{8'd172,8'd156} : s = 28;
	{8'd172,8'd157} : s = 114;
	{8'd172,8'd158} : s = 113;
	{8'd172,8'd159} : s = 242;
	{8'd172,8'd160} : s = 108;
	{8'd172,8'd161} : s = 241;
	{8'd172,8'd162} : s = 236;
	{8'd172,8'd163} : s = 399;
	{8'd172,8'd164} : s = 26;
	{8'd172,8'd165} : s = 106;
	{8'd172,8'd166} : s = 105;
	{8'd172,8'd167} : s = 234;
	{8'd172,8'd168} : s = 102;
	{8'd172,8'd169} : s = 233;
	{8'd172,8'd170} : s = 230;
	{8'd172,8'd171} : s = 380;
	{8'd172,8'd172} : s = 101;
	{8'd172,8'd173} : s = 229;
	{8'd172,8'd174} : s = 227;
	{8'd172,8'd175} : s = 378;
	{8'd172,8'd176} : s = 220;
	{8'd172,8'd177} : s = 377;
	{8'd172,8'd178} : s = 374;
	{8'd172,8'd179} : s = 487;
	{8'd172,8'd180} : s = 25;
	{8'd172,8'd181} : s = 99;
	{8'd172,8'd182} : s = 92;
	{8'd172,8'd183} : s = 218;
	{8'd172,8'd184} : s = 90;
	{8'd172,8'd185} : s = 217;
	{8'd172,8'd186} : s = 214;
	{8'd172,8'd187} : s = 373;
	{8'd172,8'd188} : s = 89;
	{8'd172,8'd189} : s = 213;
	{8'd172,8'd190} : s = 211;
	{8'd172,8'd191} : s = 371;
	{8'd172,8'd192} : s = 206;
	{8'd172,8'd193} : s = 366;
	{8'd172,8'd194} : s = 365;
	{8'd172,8'd195} : s = 478;
	{8'd172,8'd196} : s = 86;
	{8'd172,8'd197} : s = 205;
	{8'd172,8'd198} : s = 203;
	{8'd172,8'd199} : s = 363;
	{8'd172,8'd200} : s = 199;
	{8'd172,8'd201} : s = 359;
	{8'd172,8'd202} : s = 350;
	{8'd172,8'd203} : s = 477;
	{8'd172,8'd204} : s = 188;
	{8'd172,8'd205} : s = 349;
	{8'd172,8'd206} : s = 347;
	{8'd172,8'd207} : s = 475;
	{8'd172,8'd208} : s = 343;
	{8'd172,8'd209} : s = 471;
	{8'd172,8'd210} : s = 463;
	{8'd172,8'd211} : s = 509;
	{8'd172,8'd212} : s = 3;
	{8'd172,8'd213} : s = 22;
	{8'd172,8'd214} : s = 21;
	{8'd172,8'd215} : s = 85;
	{8'd172,8'd216} : s = 19;
	{8'd172,8'd217} : s = 83;
	{8'd172,8'd218} : s = 78;
	{8'd172,8'd219} : s = 186;
	{8'd172,8'd220} : s = 14;
	{8'd172,8'd221} : s = 77;
	{8'd172,8'd222} : s = 75;
	{8'd172,8'd223} : s = 185;
	{8'd172,8'd224} : s = 71;
	{8'd172,8'd225} : s = 182;
	{8'd172,8'd226} : s = 181;
	{8'd172,8'd227} : s = 335;
	{8'd172,8'd228} : s = 13;
	{8'd172,8'd229} : s = 60;
	{8'd172,8'd230} : s = 58;
	{8'd172,8'd231} : s = 179;
	{8'd172,8'd232} : s = 57;
	{8'd172,8'd233} : s = 174;
	{8'd172,8'd234} : s = 173;
	{8'd172,8'd235} : s = 318;
	{8'd172,8'd236} : s = 54;
	{8'd172,8'd237} : s = 171;
	{8'd172,8'd238} : s = 167;
	{8'd172,8'd239} : s = 317;
	{8'd172,8'd240} : s = 158;
	{8'd172,8'd241} : s = 315;
	{8'd172,8'd242} : s = 311;
	{8'd172,8'd243} : s = 446;
	{8'd172,8'd244} : s = 11;
	{8'd172,8'd245} : s = 53;
	{8'd172,8'd246} : s = 51;
	{8'd172,8'd247} : s = 157;
	{8'd172,8'd248} : s = 46;
	{8'd172,8'd249} : s = 155;
	{8'd172,8'd250} : s = 151;
	{8'd172,8'd251} : s = 303;
	{8'd172,8'd252} : s = 45;
	{8'd172,8'd253} : s = 143;
	{8'd172,8'd254} : s = 124;
	{8'd172,8'd255} : s = 287;
	{8'd173,8'd0} : s = 406;
	{8'd173,8'd1} : s = 405;
	{8'd173,8'd2} : s = 485;
	{8'd173,8'd3} : s = 112;
	{8'd173,8'd4} : s = 275;
	{8'd173,8'd5} : s = 270;
	{8'd173,8'd6} : s = 403;
	{8'd173,8'd7} : s = 269;
	{8'd173,8'd8} : s = 398;
	{8'd173,8'd9} : s = 397;
	{8'd173,8'd10} : s = 483;
	{8'd173,8'd11} : s = 267;
	{8'd173,8'd12} : s = 395;
	{8'd173,8'd13} : s = 391;
	{8'd173,8'd14} : s = 476;
	{8'd173,8'd15} : s = 376;
	{8'd173,8'd16} : s = 474;
	{8'd173,8'd17} : s = 473;
	{8'd173,8'd18} : s = 506;
	{8'd173,8'd19} : s = 20;
	{8'd173,8'd20} : s = 104;
	{8'd173,8'd21} : s = 100;
	{8'd173,8'd22} : s = 263;
	{8'd173,8'd23} : s = 98;
	{8'd173,8'd24} : s = 240;
	{8'd173,8'd25} : s = 232;
	{8'd173,8'd26} : s = 372;
	{8'd173,8'd27} : s = 97;
	{8'd173,8'd28} : s = 228;
	{8'd173,8'd29} : s = 226;
	{8'd173,8'd30} : s = 370;
	{8'd173,8'd31} : s = 225;
	{8'd173,8'd32} : s = 369;
	{8'd173,8'd33} : s = 364;
	{8'd173,8'd34} : s = 470;
	{8'd173,8'd35} : s = 88;
	{8'd173,8'd36} : s = 216;
	{8'd173,8'd37} : s = 212;
	{8'd173,8'd38} : s = 362;
	{8'd173,8'd39} : s = 210;
	{8'd173,8'd40} : s = 361;
	{8'd173,8'd41} : s = 358;
	{8'd173,8'd42} : s = 469;
	{8'd173,8'd43} : s = 209;
	{8'd173,8'd44} : s = 357;
	{8'd173,8'd45} : s = 355;
	{8'd173,8'd46} : s = 467;
	{8'd173,8'd47} : s = 348;
	{8'd173,8'd48} : s = 462;
	{8'd173,8'd49} : s = 461;
	{8'd173,8'd50} : s = 505;
	{8'd173,8'd51} : s = 84;
	{8'd173,8'd52} : s = 204;
	{8'd173,8'd53} : s = 202;
	{8'd173,8'd54} : s = 346;
	{8'd173,8'd55} : s = 201;
	{8'd173,8'd56} : s = 345;
	{8'd173,8'd57} : s = 342;
	{8'd173,8'd58} : s = 459;
	{8'd173,8'd59} : s = 198;
	{8'd173,8'd60} : s = 341;
	{8'd173,8'd61} : s = 339;
	{8'd173,8'd62} : s = 455;
	{8'd173,8'd63} : s = 334;
	{8'd173,8'd64} : s = 444;
	{8'd173,8'd65} : s = 442;
	{8'd173,8'd66} : s = 502;
	{8'd173,8'd67} : s = 197;
	{8'd173,8'd68} : s = 333;
	{8'd173,8'd69} : s = 331;
	{8'd173,8'd70} : s = 441;
	{8'd173,8'd71} : s = 327;
	{8'd173,8'd72} : s = 438;
	{8'd173,8'd73} : s = 437;
	{8'd173,8'd74} : s = 501;
	{8'd173,8'd75} : s = 316;
	{8'd173,8'd76} : s = 435;
	{8'd173,8'd77} : s = 430;
	{8'd173,8'd78} : s = 499;
	{8'd173,8'd79} : s = 429;
	{8'd173,8'd80} : s = 494;
	{8'd173,8'd81} : s = 493;
	{8'd173,8'd82} : s = 510;
	{8'd173,8'd83} : s = 1;
	{8'd173,8'd84} : s = 18;
	{8'd173,8'd85} : s = 17;
	{8'd173,8'd86} : s = 82;
	{8'd173,8'd87} : s = 12;
	{8'd173,8'd88} : s = 81;
	{8'd173,8'd89} : s = 76;
	{8'd173,8'd90} : s = 195;
	{8'd173,8'd91} : s = 10;
	{8'd173,8'd92} : s = 74;
	{8'd173,8'd93} : s = 73;
	{8'd173,8'd94} : s = 184;
	{8'd173,8'd95} : s = 70;
	{8'd173,8'd96} : s = 180;
	{8'd173,8'd97} : s = 178;
	{8'd173,8'd98} : s = 314;
	{8'd173,8'd99} : s = 9;
	{8'd173,8'd100} : s = 69;
	{8'd173,8'd101} : s = 67;
	{8'd173,8'd102} : s = 177;
	{8'd173,8'd103} : s = 56;
	{8'd173,8'd104} : s = 172;
	{8'd173,8'd105} : s = 170;
	{8'd173,8'd106} : s = 313;
	{8'd173,8'd107} : s = 52;
	{8'd173,8'd108} : s = 169;
	{8'd173,8'd109} : s = 166;
	{8'd173,8'd110} : s = 310;
	{8'd173,8'd111} : s = 165;
	{8'd173,8'd112} : s = 309;
	{8'd173,8'd113} : s = 307;
	{8'd173,8'd114} : s = 427;
	{8'd173,8'd115} : s = 6;
	{8'd173,8'd116} : s = 50;
	{8'd173,8'd117} : s = 49;
	{8'd173,8'd118} : s = 163;
	{8'd173,8'd119} : s = 44;
	{8'd173,8'd120} : s = 156;
	{8'd173,8'd121} : s = 154;
	{8'd173,8'd122} : s = 302;
	{8'd173,8'd123} : s = 42;
	{8'd173,8'd124} : s = 153;
	{8'd173,8'd125} : s = 150;
	{8'd173,8'd126} : s = 301;
	{8'd173,8'd127} : s = 149;
	{8'd173,8'd128} : s = 299;
	{8'd173,8'd129} : s = 295;
	{8'd173,8'd130} : s = 423;
	{8'd173,8'd131} : s = 41;
	{8'd173,8'd132} : s = 147;
	{8'd173,8'd133} : s = 142;
	{8'd173,8'd134} : s = 286;
	{8'd173,8'd135} : s = 141;
	{8'd173,8'd136} : s = 285;
	{8'd173,8'd137} : s = 283;
	{8'd173,8'd138} : s = 414;
	{8'd173,8'd139} : s = 139;
	{8'd173,8'd140} : s = 279;
	{8'd173,8'd141} : s = 271;
	{8'd173,8'd142} : s = 413;
	{8'd173,8'd143} : s = 248;
	{8'd173,8'd144} : s = 411;
	{8'd173,8'd145} : s = 407;
	{8'd173,8'd146} : s = 491;
	{8'd173,8'd147} : s = 5;
	{8'd173,8'd148} : s = 38;
	{8'd173,8'd149} : s = 37;
	{8'd173,8'd150} : s = 135;
	{8'd173,8'd151} : s = 35;
	{8'd173,8'd152} : s = 120;
	{8'd173,8'd153} : s = 116;
	{8'd173,8'd154} : s = 244;
	{8'd173,8'd155} : s = 28;
	{8'd173,8'd156} : s = 114;
	{8'd173,8'd157} : s = 113;
	{8'd173,8'd158} : s = 242;
	{8'd173,8'd159} : s = 108;
	{8'd173,8'd160} : s = 241;
	{8'd173,8'd161} : s = 236;
	{8'd173,8'd162} : s = 399;
	{8'd173,8'd163} : s = 26;
	{8'd173,8'd164} : s = 106;
	{8'd173,8'd165} : s = 105;
	{8'd173,8'd166} : s = 234;
	{8'd173,8'd167} : s = 102;
	{8'd173,8'd168} : s = 233;
	{8'd173,8'd169} : s = 230;
	{8'd173,8'd170} : s = 380;
	{8'd173,8'd171} : s = 101;
	{8'd173,8'd172} : s = 229;
	{8'd173,8'd173} : s = 227;
	{8'd173,8'd174} : s = 378;
	{8'd173,8'd175} : s = 220;
	{8'd173,8'd176} : s = 377;
	{8'd173,8'd177} : s = 374;
	{8'd173,8'd178} : s = 487;
	{8'd173,8'd179} : s = 25;
	{8'd173,8'd180} : s = 99;
	{8'd173,8'd181} : s = 92;
	{8'd173,8'd182} : s = 218;
	{8'd173,8'd183} : s = 90;
	{8'd173,8'd184} : s = 217;
	{8'd173,8'd185} : s = 214;
	{8'd173,8'd186} : s = 373;
	{8'd173,8'd187} : s = 89;
	{8'd173,8'd188} : s = 213;
	{8'd173,8'd189} : s = 211;
	{8'd173,8'd190} : s = 371;
	{8'd173,8'd191} : s = 206;
	{8'd173,8'd192} : s = 366;
	{8'd173,8'd193} : s = 365;
	{8'd173,8'd194} : s = 478;
	{8'd173,8'd195} : s = 86;
	{8'd173,8'd196} : s = 205;
	{8'd173,8'd197} : s = 203;
	{8'd173,8'd198} : s = 363;
	{8'd173,8'd199} : s = 199;
	{8'd173,8'd200} : s = 359;
	{8'd173,8'd201} : s = 350;
	{8'd173,8'd202} : s = 477;
	{8'd173,8'd203} : s = 188;
	{8'd173,8'd204} : s = 349;
	{8'd173,8'd205} : s = 347;
	{8'd173,8'd206} : s = 475;
	{8'd173,8'd207} : s = 343;
	{8'd173,8'd208} : s = 471;
	{8'd173,8'd209} : s = 463;
	{8'd173,8'd210} : s = 509;
	{8'd173,8'd211} : s = 3;
	{8'd173,8'd212} : s = 22;
	{8'd173,8'd213} : s = 21;
	{8'd173,8'd214} : s = 85;
	{8'd173,8'd215} : s = 19;
	{8'd173,8'd216} : s = 83;
	{8'd173,8'd217} : s = 78;
	{8'd173,8'd218} : s = 186;
	{8'd173,8'd219} : s = 14;
	{8'd173,8'd220} : s = 77;
	{8'd173,8'd221} : s = 75;
	{8'd173,8'd222} : s = 185;
	{8'd173,8'd223} : s = 71;
	{8'd173,8'd224} : s = 182;
	{8'd173,8'd225} : s = 181;
	{8'd173,8'd226} : s = 335;
	{8'd173,8'd227} : s = 13;
	{8'd173,8'd228} : s = 60;
	{8'd173,8'd229} : s = 58;
	{8'd173,8'd230} : s = 179;
	{8'd173,8'd231} : s = 57;
	{8'd173,8'd232} : s = 174;
	{8'd173,8'd233} : s = 173;
	{8'd173,8'd234} : s = 318;
	{8'd173,8'd235} : s = 54;
	{8'd173,8'd236} : s = 171;
	{8'd173,8'd237} : s = 167;
	{8'd173,8'd238} : s = 317;
	{8'd173,8'd239} : s = 158;
	{8'd173,8'd240} : s = 315;
	{8'd173,8'd241} : s = 311;
	{8'd173,8'd242} : s = 446;
	{8'd173,8'd243} : s = 11;
	{8'd173,8'd244} : s = 53;
	{8'd173,8'd245} : s = 51;
	{8'd173,8'd246} : s = 157;
	{8'd173,8'd247} : s = 46;
	{8'd173,8'd248} : s = 155;
	{8'd173,8'd249} : s = 151;
	{8'd173,8'd250} : s = 303;
	{8'd173,8'd251} : s = 45;
	{8'd173,8'd252} : s = 143;
	{8'd173,8'd253} : s = 124;
	{8'd173,8'd254} : s = 287;
	{8'd173,8'd255} : s = 122;
	{8'd174,8'd0} : s = 405;
	{8'd174,8'd1} : s = 485;
	{8'd174,8'd2} : s = 112;
	{8'd174,8'd3} : s = 275;
	{8'd174,8'd4} : s = 270;
	{8'd174,8'd5} : s = 403;
	{8'd174,8'd6} : s = 269;
	{8'd174,8'd7} : s = 398;
	{8'd174,8'd8} : s = 397;
	{8'd174,8'd9} : s = 483;
	{8'd174,8'd10} : s = 267;
	{8'd174,8'd11} : s = 395;
	{8'd174,8'd12} : s = 391;
	{8'd174,8'd13} : s = 476;
	{8'd174,8'd14} : s = 376;
	{8'd174,8'd15} : s = 474;
	{8'd174,8'd16} : s = 473;
	{8'd174,8'd17} : s = 506;
	{8'd174,8'd18} : s = 20;
	{8'd174,8'd19} : s = 104;
	{8'd174,8'd20} : s = 100;
	{8'd174,8'd21} : s = 263;
	{8'd174,8'd22} : s = 98;
	{8'd174,8'd23} : s = 240;
	{8'd174,8'd24} : s = 232;
	{8'd174,8'd25} : s = 372;
	{8'd174,8'd26} : s = 97;
	{8'd174,8'd27} : s = 228;
	{8'd174,8'd28} : s = 226;
	{8'd174,8'd29} : s = 370;
	{8'd174,8'd30} : s = 225;
	{8'd174,8'd31} : s = 369;
	{8'd174,8'd32} : s = 364;
	{8'd174,8'd33} : s = 470;
	{8'd174,8'd34} : s = 88;
	{8'd174,8'd35} : s = 216;
	{8'd174,8'd36} : s = 212;
	{8'd174,8'd37} : s = 362;
	{8'd174,8'd38} : s = 210;
	{8'd174,8'd39} : s = 361;
	{8'd174,8'd40} : s = 358;
	{8'd174,8'd41} : s = 469;
	{8'd174,8'd42} : s = 209;
	{8'd174,8'd43} : s = 357;
	{8'd174,8'd44} : s = 355;
	{8'd174,8'd45} : s = 467;
	{8'd174,8'd46} : s = 348;
	{8'd174,8'd47} : s = 462;
	{8'd174,8'd48} : s = 461;
	{8'd174,8'd49} : s = 505;
	{8'd174,8'd50} : s = 84;
	{8'd174,8'd51} : s = 204;
	{8'd174,8'd52} : s = 202;
	{8'd174,8'd53} : s = 346;
	{8'd174,8'd54} : s = 201;
	{8'd174,8'd55} : s = 345;
	{8'd174,8'd56} : s = 342;
	{8'd174,8'd57} : s = 459;
	{8'd174,8'd58} : s = 198;
	{8'd174,8'd59} : s = 341;
	{8'd174,8'd60} : s = 339;
	{8'd174,8'd61} : s = 455;
	{8'd174,8'd62} : s = 334;
	{8'd174,8'd63} : s = 444;
	{8'd174,8'd64} : s = 442;
	{8'd174,8'd65} : s = 502;
	{8'd174,8'd66} : s = 197;
	{8'd174,8'd67} : s = 333;
	{8'd174,8'd68} : s = 331;
	{8'd174,8'd69} : s = 441;
	{8'd174,8'd70} : s = 327;
	{8'd174,8'd71} : s = 438;
	{8'd174,8'd72} : s = 437;
	{8'd174,8'd73} : s = 501;
	{8'd174,8'd74} : s = 316;
	{8'd174,8'd75} : s = 435;
	{8'd174,8'd76} : s = 430;
	{8'd174,8'd77} : s = 499;
	{8'd174,8'd78} : s = 429;
	{8'd174,8'd79} : s = 494;
	{8'd174,8'd80} : s = 493;
	{8'd174,8'd81} : s = 510;
	{8'd174,8'd82} : s = 1;
	{8'd174,8'd83} : s = 18;
	{8'd174,8'd84} : s = 17;
	{8'd174,8'd85} : s = 82;
	{8'd174,8'd86} : s = 12;
	{8'd174,8'd87} : s = 81;
	{8'd174,8'd88} : s = 76;
	{8'd174,8'd89} : s = 195;
	{8'd174,8'd90} : s = 10;
	{8'd174,8'd91} : s = 74;
	{8'd174,8'd92} : s = 73;
	{8'd174,8'd93} : s = 184;
	{8'd174,8'd94} : s = 70;
	{8'd174,8'd95} : s = 180;
	{8'd174,8'd96} : s = 178;
	{8'd174,8'd97} : s = 314;
	{8'd174,8'd98} : s = 9;
	{8'd174,8'd99} : s = 69;
	{8'd174,8'd100} : s = 67;
	{8'd174,8'd101} : s = 177;
	{8'd174,8'd102} : s = 56;
	{8'd174,8'd103} : s = 172;
	{8'd174,8'd104} : s = 170;
	{8'd174,8'd105} : s = 313;
	{8'd174,8'd106} : s = 52;
	{8'd174,8'd107} : s = 169;
	{8'd174,8'd108} : s = 166;
	{8'd174,8'd109} : s = 310;
	{8'd174,8'd110} : s = 165;
	{8'd174,8'd111} : s = 309;
	{8'd174,8'd112} : s = 307;
	{8'd174,8'd113} : s = 427;
	{8'd174,8'd114} : s = 6;
	{8'd174,8'd115} : s = 50;
	{8'd174,8'd116} : s = 49;
	{8'd174,8'd117} : s = 163;
	{8'd174,8'd118} : s = 44;
	{8'd174,8'd119} : s = 156;
	{8'd174,8'd120} : s = 154;
	{8'd174,8'd121} : s = 302;
	{8'd174,8'd122} : s = 42;
	{8'd174,8'd123} : s = 153;
	{8'd174,8'd124} : s = 150;
	{8'd174,8'd125} : s = 301;
	{8'd174,8'd126} : s = 149;
	{8'd174,8'd127} : s = 299;
	{8'd174,8'd128} : s = 295;
	{8'd174,8'd129} : s = 423;
	{8'd174,8'd130} : s = 41;
	{8'd174,8'd131} : s = 147;
	{8'd174,8'd132} : s = 142;
	{8'd174,8'd133} : s = 286;
	{8'd174,8'd134} : s = 141;
	{8'd174,8'd135} : s = 285;
	{8'd174,8'd136} : s = 283;
	{8'd174,8'd137} : s = 414;
	{8'd174,8'd138} : s = 139;
	{8'd174,8'd139} : s = 279;
	{8'd174,8'd140} : s = 271;
	{8'd174,8'd141} : s = 413;
	{8'd174,8'd142} : s = 248;
	{8'd174,8'd143} : s = 411;
	{8'd174,8'd144} : s = 407;
	{8'd174,8'd145} : s = 491;
	{8'd174,8'd146} : s = 5;
	{8'd174,8'd147} : s = 38;
	{8'd174,8'd148} : s = 37;
	{8'd174,8'd149} : s = 135;
	{8'd174,8'd150} : s = 35;
	{8'd174,8'd151} : s = 120;
	{8'd174,8'd152} : s = 116;
	{8'd174,8'd153} : s = 244;
	{8'd174,8'd154} : s = 28;
	{8'd174,8'd155} : s = 114;
	{8'd174,8'd156} : s = 113;
	{8'd174,8'd157} : s = 242;
	{8'd174,8'd158} : s = 108;
	{8'd174,8'd159} : s = 241;
	{8'd174,8'd160} : s = 236;
	{8'd174,8'd161} : s = 399;
	{8'd174,8'd162} : s = 26;
	{8'd174,8'd163} : s = 106;
	{8'd174,8'd164} : s = 105;
	{8'd174,8'd165} : s = 234;
	{8'd174,8'd166} : s = 102;
	{8'd174,8'd167} : s = 233;
	{8'd174,8'd168} : s = 230;
	{8'd174,8'd169} : s = 380;
	{8'd174,8'd170} : s = 101;
	{8'd174,8'd171} : s = 229;
	{8'd174,8'd172} : s = 227;
	{8'd174,8'd173} : s = 378;
	{8'd174,8'd174} : s = 220;
	{8'd174,8'd175} : s = 377;
	{8'd174,8'd176} : s = 374;
	{8'd174,8'd177} : s = 487;
	{8'd174,8'd178} : s = 25;
	{8'd174,8'd179} : s = 99;
	{8'd174,8'd180} : s = 92;
	{8'd174,8'd181} : s = 218;
	{8'd174,8'd182} : s = 90;
	{8'd174,8'd183} : s = 217;
	{8'd174,8'd184} : s = 214;
	{8'd174,8'd185} : s = 373;
	{8'd174,8'd186} : s = 89;
	{8'd174,8'd187} : s = 213;
	{8'd174,8'd188} : s = 211;
	{8'd174,8'd189} : s = 371;
	{8'd174,8'd190} : s = 206;
	{8'd174,8'd191} : s = 366;
	{8'd174,8'd192} : s = 365;
	{8'd174,8'd193} : s = 478;
	{8'd174,8'd194} : s = 86;
	{8'd174,8'd195} : s = 205;
	{8'd174,8'd196} : s = 203;
	{8'd174,8'd197} : s = 363;
	{8'd174,8'd198} : s = 199;
	{8'd174,8'd199} : s = 359;
	{8'd174,8'd200} : s = 350;
	{8'd174,8'd201} : s = 477;
	{8'd174,8'd202} : s = 188;
	{8'd174,8'd203} : s = 349;
	{8'd174,8'd204} : s = 347;
	{8'd174,8'd205} : s = 475;
	{8'd174,8'd206} : s = 343;
	{8'd174,8'd207} : s = 471;
	{8'd174,8'd208} : s = 463;
	{8'd174,8'd209} : s = 509;
	{8'd174,8'd210} : s = 3;
	{8'd174,8'd211} : s = 22;
	{8'd174,8'd212} : s = 21;
	{8'd174,8'd213} : s = 85;
	{8'd174,8'd214} : s = 19;
	{8'd174,8'd215} : s = 83;
	{8'd174,8'd216} : s = 78;
	{8'd174,8'd217} : s = 186;
	{8'd174,8'd218} : s = 14;
	{8'd174,8'd219} : s = 77;
	{8'd174,8'd220} : s = 75;
	{8'd174,8'd221} : s = 185;
	{8'd174,8'd222} : s = 71;
	{8'd174,8'd223} : s = 182;
	{8'd174,8'd224} : s = 181;
	{8'd174,8'd225} : s = 335;
	{8'd174,8'd226} : s = 13;
	{8'd174,8'd227} : s = 60;
	{8'd174,8'd228} : s = 58;
	{8'd174,8'd229} : s = 179;
	{8'd174,8'd230} : s = 57;
	{8'd174,8'd231} : s = 174;
	{8'd174,8'd232} : s = 173;
	{8'd174,8'd233} : s = 318;
	{8'd174,8'd234} : s = 54;
	{8'd174,8'd235} : s = 171;
	{8'd174,8'd236} : s = 167;
	{8'd174,8'd237} : s = 317;
	{8'd174,8'd238} : s = 158;
	{8'd174,8'd239} : s = 315;
	{8'd174,8'd240} : s = 311;
	{8'd174,8'd241} : s = 446;
	{8'd174,8'd242} : s = 11;
	{8'd174,8'd243} : s = 53;
	{8'd174,8'd244} : s = 51;
	{8'd174,8'd245} : s = 157;
	{8'd174,8'd246} : s = 46;
	{8'd174,8'd247} : s = 155;
	{8'd174,8'd248} : s = 151;
	{8'd174,8'd249} : s = 303;
	{8'd174,8'd250} : s = 45;
	{8'd174,8'd251} : s = 143;
	{8'd174,8'd252} : s = 124;
	{8'd174,8'd253} : s = 287;
	{8'd174,8'd254} : s = 122;
	{8'd174,8'd255} : s = 252;
	{8'd175,8'd0} : s = 485;
	{8'd175,8'd1} : s = 112;
	{8'd175,8'd2} : s = 275;
	{8'd175,8'd3} : s = 270;
	{8'd175,8'd4} : s = 403;
	{8'd175,8'd5} : s = 269;
	{8'd175,8'd6} : s = 398;
	{8'd175,8'd7} : s = 397;
	{8'd175,8'd8} : s = 483;
	{8'd175,8'd9} : s = 267;
	{8'd175,8'd10} : s = 395;
	{8'd175,8'd11} : s = 391;
	{8'd175,8'd12} : s = 476;
	{8'd175,8'd13} : s = 376;
	{8'd175,8'd14} : s = 474;
	{8'd175,8'd15} : s = 473;
	{8'd175,8'd16} : s = 506;
	{8'd175,8'd17} : s = 20;
	{8'd175,8'd18} : s = 104;
	{8'd175,8'd19} : s = 100;
	{8'd175,8'd20} : s = 263;
	{8'd175,8'd21} : s = 98;
	{8'd175,8'd22} : s = 240;
	{8'd175,8'd23} : s = 232;
	{8'd175,8'd24} : s = 372;
	{8'd175,8'd25} : s = 97;
	{8'd175,8'd26} : s = 228;
	{8'd175,8'd27} : s = 226;
	{8'd175,8'd28} : s = 370;
	{8'd175,8'd29} : s = 225;
	{8'd175,8'd30} : s = 369;
	{8'd175,8'd31} : s = 364;
	{8'd175,8'd32} : s = 470;
	{8'd175,8'd33} : s = 88;
	{8'd175,8'd34} : s = 216;
	{8'd175,8'd35} : s = 212;
	{8'd175,8'd36} : s = 362;
	{8'd175,8'd37} : s = 210;
	{8'd175,8'd38} : s = 361;
	{8'd175,8'd39} : s = 358;
	{8'd175,8'd40} : s = 469;
	{8'd175,8'd41} : s = 209;
	{8'd175,8'd42} : s = 357;
	{8'd175,8'd43} : s = 355;
	{8'd175,8'd44} : s = 467;
	{8'd175,8'd45} : s = 348;
	{8'd175,8'd46} : s = 462;
	{8'd175,8'd47} : s = 461;
	{8'd175,8'd48} : s = 505;
	{8'd175,8'd49} : s = 84;
	{8'd175,8'd50} : s = 204;
	{8'd175,8'd51} : s = 202;
	{8'd175,8'd52} : s = 346;
	{8'd175,8'd53} : s = 201;
	{8'd175,8'd54} : s = 345;
	{8'd175,8'd55} : s = 342;
	{8'd175,8'd56} : s = 459;
	{8'd175,8'd57} : s = 198;
	{8'd175,8'd58} : s = 341;
	{8'd175,8'd59} : s = 339;
	{8'd175,8'd60} : s = 455;
	{8'd175,8'd61} : s = 334;
	{8'd175,8'd62} : s = 444;
	{8'd175,8'd63} : s = 442;
	{8'd175,8'd64} : s = 502;
	{8'd175,8'd65} : s = 197;
	{8'd175,8'd66} : s = 333;
	{8'd175,8'd67} : s = 331;
	{8'd175,8'd68} : s = 441;
	{8'd175,8'd69} : s = 327;
	{8'd175,8'd70} : s = 438;
	{8'd175,8'd71} : s = 437;
	{8'd175,8'd72} : s = 501;
	{8'd175,8'd73} : s = 316;
	{8'd175,8'd74} : s = 435;
	{8'd175,8'd75} : s = 430;
	{8'd175,8'd76} : s = 499;
	{8'd175,8'd77} : s = 429;
	{8'd175,8'd78} : s = 494;
	{8'd175,8'd79} : s = 493;
	{8'd175,8'd80} : s = 510;
	{8'd175,8'd81} : s = 1;
	{8'd175,8'd82} : s = 18;
	{8'd175,8'd83} : s = 17;
	{8'd175,8'd84} : s = 82;
	{8'd175,8'd85} : s = 12;
	{8'd175,8'd86} : s = 81;
	{8'd175,8'd87} : s = 76;
	{8'd175,8'd88} : s = 195;
	{8'd175,8'd89} : s = 10;
	{8'd175,8'd90} : s = 74;
	{8'd175,8'd91} : s = 73;
	{8'd175,8'd92} : s = 184;
	{8'd175,8'd93} : s = 70;
	{8'd175,8'd94} : s = 180;
	{8'd175,8'd95} : s = 178;
	{8'd175,8'd96} : s = 314;
	{8'd175,8'd97} : s = 9;
	{8'd175,8'd98} : s = 69;
	{8'd175,8'd99} : s = 67;
	{8'd175,8'd100} : s = 177;
	{8'd175,8'd101} : s = 56;
	{8'd175,8'd102} : s = 172;
	{8'd175,8'd103} : s = 170;
	{8'd175,8'd104} : s = 313;
	{8'd175,8'd105} : s = 52;
	{8'd175,8'd106} : s = 169;
	{8'd175,8'd107} : s = 166;
	{8'd175,8'd108} : s = 310;
	{8'd175,8'd109} : s = 165;
	{8'd175,8'd110} : s = 309;
	{8'd175,8'd111} : s = 307;
	{8'd175,8'd112} : s = 427;
	{8'd175,8'd113} : s = 6;
	{8'd175,8'd114} : s = 50;
	{8'd175,8'd115} : s = 49;
	{8'd175,8'd116} : s = 163;
	{8'd175,8'd117} : s = 44;
	{8'd175,8'd118} : s = 156;
	{8'd175,8'd119} : s = 154;
	{8'd175,8'd120} : s = 302;
	{8'd175,8'd121} : s = 42;
	{8'd175,8'd122} : s = 153;
	{8'd175,8'd123} : s = 150;
	{8'd175,8'd124} : s = 301;
	{8'd175,8'd125} : s = 149;
	{8'd175,8'd126} : s = 299;
	{8'd175,8'd127} : s = 295;
	{8'd175,8'd128} : s = 423;
	{8'd175,8'd129} : s = 41;
	{8'd175,8'd130} : s = 147;
	{8'd175,8'd131} : s = 142;
	{8'd175,8'd132} : s = 286;
	{8'd175,8'd133} : s = 141;
	{8'd175,8'd134} : s = 285;
	{8'd175,8'd135} : s = 283;
	{8'd175,8'd136} : s = 414;
	{8'd175,8'd137} : s = 139;
	{8'd175,8'd138} : s = 279;
	{8'd175,8'd139} : s = 271;
	{8'd175,8'd140} : s = 413;
	{8'd175,8'd141} : s = 248;
	{8'd175,8'd142} : s = 411;
	{8'd175,8'd143} : s = 407;
	{8'd175,8'd144} : s = 491;
	{8'd175,8'd145} : s = 5;
	{8'd175,8'd146} : s = 38;
	{8'd175,8'd147} : s = 37;
	{8'd175,8'd148} : s = 135;
	{8'd175,8'd149} : s = 35;
	{8'd175,8'd150} : s = 120;
	{8'd175,8'd151} : s = 116;
	{8'd175,8'd152} : s = 244;
	{8'd175,8'd153} : s = 28;
	{8'd175,8'd154} : s = 114;
	{8'd175,8'd155} : s = 113;
	{8'd175,8'd156} : s = 242;
	{8'd175,8'd157} : s = 108;
	{8'd175,8'd158} : s = 241;
	{8'd175,8'd159} : s = 236;
	{8'd175,8'd160} : s = 399;
	{8'd175,8'd161} : s = 26;
	{8'd175,8'd162} : s = 106;
	{8'd175,8'd163} : s = 105;
	{8'd175,8'd164} : s = 234;
	{8'd175,8'd165} : s = 102;
	{8'd175,8'd166} : s = 233;
	{8'd175,8'd167} : s = 230;
	{8'd175,8'd168} : s = 380;
	{8'd175,8'd169} : s = 101;
	{8'd175,8'd170} : s = 229;
	{8'd175,8'd171} : s = 227;
	{8'd175,8'd172} : s = 378;
	{8'd175,8'd173} : s = 220;
	{8'd175,8'd174} : s = 377;
	{8'd175,8'd175} : s = 374;
	{8'd175,8'd176} : s = 487;
	{8'd175,8'd177} : s = 25;
	{8'd175,8'd178} : s = 99;
	{8'd175,8'd179} : s = 92;
	{8'd175,8'd180} : s = 218;
	{8'd175,8'd181} : s = 90;
	{8'd175,8'd182} : s = 217;
	{8'd175,8'd183} : s = 214;
	{8'd175,8'd184} : s = 373;
	{8'd175,8'd185} : s = 89;
	{8'd175,8'd186} : s = 213;
	{8'd175,8'd187} : s = 211;
	{8'd175,8'd188} : s = 371;
	{8'd175,8'd189} : s = 206;
	{8'd175,8'd190} : s = 366;
	{8'd175,8'd191} : s = 365;
	{8'd175,8'd192} : s = 478;
	{8'd175,8'd193} : s = 86;
	{8'd175,8'd194} : s = 205;
	{8'd175,8'd195} : s = 203;
	{8'd175,8'd196} : s = 363;
	{8'd175,8'd197} : s = 199;
	{8'd175,8'd198} : s = 359;
	{8'd175,8'd199} : s = 350;
	{8'd175,8'd200} : s = 477;
	{8'd175,8'd201} : s = 188;
	{8'd175,8'd202} : s = 349;
	{8'd175,8'd203} : s = 347;
	{8'd175,8'd204} : s = 475;
	{8'd175,8'd205} : s = 343;
	{8'd175,8'd206} : s = 471;
	{8'd175,8'd207} : s = 463;
	{8'd175,8'd208} : s = 509;
	{8'd175,8'd209} : s = 3;
	{8'd175,8'd210} : s = 22;
	{8'd175,8'd211} : s = 21;
	{8'd175,8'd212} : s = 85;
	{8'd175,8'd213} : s = 19;
	{8'd175,8'd214} : s = 83;
	{8'd175,8'd215} : s = 78;
	{8'd175,8'd216} : s = 186;
	{8'd175,8'd217} : s = 14;
	{8'd175,8'd218} : s = 77;
	{8'd175,8'd219} : s = 75;
	{8'd175,8'd220} : s = 185;
	{8'd175,8'd221} : s = 71;
	{8'd175,8'd222} : s = 182;
	{8'd175,8'd223} : s = 181;
	{8'd175,8'd224} : s = 335;
	{8'd175,8'd225} : s = 13;
	{8'd175,8'd226} : s = 60;
	{8'd175,8'd227} : s = 58;
	{8'd175,8'd228} : s = 179;
	{8'd175,8'd229} : s = 57;
	{8'd175,8'd230} : s = 174;
	{8'd175,8'd231} : s = 173;
	{8'd175,8'd232} : s = 318;
	{8'd175,8'd233} : s = 54;
	{8'd175,8'd234} : s = 171;
	{8'd175,8'd235} : s = 167;
	{8'd175,8'd236} : s = 317;
	{8'd175,8'd237} : s = 158;
	{8'd175,8'd238} : s = 315;
	{8'd175,8'd239} : s = 311;
	{8'd175,8'd240} : s = 446;
	{8'd175,8'd241} : s = 11;
	{8'd175,8'd242} : s = 53;
	{8'd175,8'd243} : s = 51;
	{8'd175,8'd244} : s = 157;
	{8'd175,8'd245} : s = 46;
	{8'd175,8'd246} : s = 155;
	{8'd175,8'd247} : s = 151;
	{8'd175,8'd248} : s = 303;
	{8'd175,8'd249} : s = 45;
	{8'd175,8'd250} : s = 143;
	{8'd175,8'd251} : s = 124;
	{8'd175,8'd252} : s = 287;
	{8'd175,8'd253} : s = 122;
	{8'd175,8'd254} : s = 252;
	{8'd175,8'd255} : s = 250;
	{8'd176,8'd0} : s = 112;
	{8'd176,8'd1} : s = 275;
	{8'd176,8'd2} : s = 270;
	{8'd176,8'd3} : s = 403;
	{8'd176,8'd4} : s = 269;
	{8'd176,8'd5} : s = 398;
	{8'd176,8'd6} : s = 397;
	{8'd176,8'd7} : s = 483;
	{8'd176,8'd8} : s = 267;
	{8'd176,8'd9} : s = 395;
	{8'd176,8'd10} : s = 391;
	{8'd176,8'd11} : s = 476;
	{8'd176,8'd12} : s = 376;
	{8'd176,8'd13} : s = 474;
	{8'd176,8'd14} : s = 473;
	{8'd176,8'd15} : s = 506;
	{8'd176,8'd16} : s = 20;
	{8'd176,8'd17} : s = 104;
	{8'd176,8'd18} : s = 100;
	{8'd176,8'd19} : s = 263;
	{8'd176,8'd20} : s = 98;
	{8'd176,8'd21} : s = 240;
	{8'd176,8'd22} : s = 232;
	{8'd176,8'd23} : s = 372;
	{8'd176,8'd24} : s = 97;
	{8'd176,8'd25} : s = 228;
	{8'd176,8'd26} : s = 226;
	{8'd176,8'd27} : s = 370;
	{8'd176,8'd28} : s = 225;
	{8'd176,8'd29} : s = 369;
	{8'd176,8'd30} : s = 364;
	{8'd176,8'd31} : s = 470;
	{8'd176,8'd32} : s = 88;
	{8'd176,8'd33} : s = 216;
	{8'd176,8'd34} : s = 212;
	{8'd176,8'd35} : s = 362;
	{8'd176,8'd36} : s = 210;
	{8'd176,8'd37} : s = 361;
	{8'd176,8'd38} : s = 358;
	{8'd176,8'd39} : s = 469;
	{8'd176,8'd40} : s = 209;
	{8'd176,8'd41} : s = 357;
	{8'd176,8'd42} : s = 355;
	{8'd176,8'd43} : s = 467;
	{8'd176,8'd44} : s = 348;
	{8'd176,8'd45} : s = 462;
	{8'd176,8'd46} : s = 461;
	{8'd176,8'd47} : s = 505;
	{8'd176,8'd48} : s = 84;
	{8'd176,8'd49} : s = 204;
	{8'd176,8'd50} : s = 202;
	{8'd176,8'd51} : s = 346;
	{8'd176,8'd52} : s = 201;
	{8'd176,8'd53} : s = 345;
	{8'd176,8'd54} : s = 342;
	{8'd176,8'd55} : s = 459;
	{8'd176,8'd56} : s = 198;
	{8'd176,8'd57} : s = 341;
	{8'd176,8'd58} : s = 339;
	{8'd176,8'd59} : s = 455;
	{8'd176,8'd60} : s = 334;
	{8'd176,8'd61} : s = 444;
	{8'd176,8'd62} : s = 442;
	{8'd176,8'd63} : s = 502;
	{8'd176,8'd64} : s = 197;
	{8'd176,8'd65} : s = 333;
	{8'd176,8'd66} : s = 331;
	{8'd176,8'd67} : s = 441;
	{8'd176,8'd68} : s = 327;
	{8'd176,8'd69} : s = 438;
	{8'd176,8'd70} : s = 437;
	{8'd176,8'd71} : s = 501;
	{8'd176,8'd72} : s = 316;
	{8'd176,8'd73} : s = 435;
	{8'd176,8'd74} : s = 430;
	{8'd176,8'd75} : s = 499;
	{8'd176,8'd76} : s = 429;
	{8'd176,8'd77} : s = 494;
	{8'd176,8'd78} : s = 493;
	{8'd176,8'd79} : s = 510;
	{8'd176,8'd80} : s = 1;
	{8'd176,8'd81} : s = 18;
	{8'd176,8'd82} : s = 17;
	{8'd176,8'd83} : s = 82;
	{8'd176,8'd84} : s = 12;
	{8'd176,8'd85} : s = 81;
	{8'd176,8'd86} : s = 76;
	{8'd176,8'd87} : s = 195;
	{8'd176,8'd88} : s = 10;
	{8'd176,8'd89} : s = 74;
	{8'd176,8'd90} : s = 73;
	{8'd176,8'd91} : s = 184;
	{8'd176,8'd92} : s = 70;
	{8'd176,8'd93} : s = 180;
	{8'd176,8'd94} : s = 178;
	{8'd176,8'd95} : s = 314;
	{8'd176,8'd96} : s = 9;
	{8'd176,8'd97} : s = 69;
	{8'd176,8'd98} : s = 67;
	{8'd176,8'd99} : s = 177;
	{8'd176,8'd100} : s = 56;
	{8'd176,8'd101} : s = 172;
	{8'd176,8'd102} : s = 170;
	{8'd176,8'd103} : s = 313;
	{8'd176,8'd104} : s = 52;
	{8'd176,8'd105} : s = 169;
	{8'd176,8'd106} : s = 166;
	{8'd176,8'd107} : s = 310;
	{8'd176,8'd108} : s = 165;
	{8'd176,8'd109} : s = 309;
	{8'd176,8'd110} : s = 307;
	{8'd176,8'd111} : s = 427;
	{8'd176,8'd112} : s = 6;
	{8'd176,8'd113} : s = 50;
	{8'd176,8'd114} : s = 49;
	{8'd176,8'd115} : s = 163;
	{8'd176,8'd116} : s = 44;
	{8'd176,8'd117} : s = 156;
	{8'd176,8'd118} : s = 154;
	{8'd176,8'd119} : s = 302;
	{8'd176,8'd120} : s = 42;
	{8'd176,8'd121} : s = 153;
	{8'd176,8'd122} : s = 150;
	{8'd176,8'd123} : s = 301;
	{8'd176,8'd124} : s = 149;
	{8'd176,8'd125} : s = 299;
	{8'd176,8'd126} : s = 295;
	{8'd176,8'd127} : s = 423;
	{8'd176,8'd128} : s = 41;
	{8'd176,8'd129} : s = 147;
	{8'd176,8'd130} : s = 142;
	{8'd176,8'd131} : s = 286;
	{8'd176,8'd132} : s = 141;
	{8'd176,8'd133} : s = 285;
	{8'd176,8'd134} : s = 283;
	{8'd176,8'd135} : s = 414;
	{8'd176,8'd136} : s = 139;
	{8'd176,8'd137} : s = 279;
	{8'd176,8'd138} : s = 271;
	{8'd176,8'd139} : s = 413;
	{8'd176,8'd140} : s = 248;
	{8'd176,8'd141} : s = 411;
	{8'd176,8'd142} : s = 407;
	{8'd176,8'd143} : s = 491;
	{8'd176,8'd144} : s = 5;
	{8'd176,8'd145} : s = 38;
	{8'd176,8'd146} : s = 37;
	{8'd176,8'd147} : s = 135;
	{8'd176,8'd148} : s = 35;
	{8'd176,8'd149} : s = 120;
	{8'd176,8'd150} : s = 116;
	{8'd176,8'd151} : s = 244;
	{8'd176,8'd152} : s = 28;
	{8'd176,8'd153} : s = 114;
	{8'd176,8'd154} : s = 113;
	{8'd176,8'd155} : s = 242;
	{8'd176,8'd156} : s = 108;
	{8'd176,8'd157} : s = 241;
	{8'd176,8'd158} : s = 236;
	{8'd176,8'd159} : s = 399;
	{8'd176,8'd160} : s = 26;
	{8'd176,8'd161} : s = 106;
	{8'd176,8'd162} : s = 105;
	{8'd176,8'd163} : s = 234;
	{8'd176,8'd164} : s = 102;
	{8'd176,8'd165} : s = 233;
	{8'd176,8'd166} : s = 230;
	{8'd176,8'd167} : s = 380;
	{8'd176,8'd168} : s = 101;
	{8'd176,8'd169} : s = 229;
	{8'd176,8'd170} : s = 227;
	{8'd176,8'd171} : s = 378;
	{8'd176,8'd172} : s = 220;
	{8'd176,8'd173} : s = 377;
	{8'd176,8'd174} : s = 374;
	{8'd176,8'd175} : s = 487;
	{8'd176,8'd176} : s = 25;
	{8'd176,8'd177} : s = 99;
	{8'd176,8'd178} : s = 92;
	{8'd176,8'd179} : s = 218;
	{8'd176,8'd180} : s = 90;
	{8'd176,8'd181} : s = 217;
	{8'd176,8'd182} : s = 214;
	{8'd176,8'd183} : s = 373;
	{8'd176,8'd184} : s = 89;
	{8'd176,8'd185} : s = 213;
	{8'd176,8'd186} : s = 211;
	{8'd176,8'd187} : s = 371;
	{8'd176,8'd188} : s = 206;
	{8'd176,8'd189} : s = 366;
	{8'd176,8'd190} : s = 365;
	{8'd176,8'd191} : s = 478;
	{8'd176,8'd192} : s = 86;
	{8'd176,8'd193} : s = 205;
	{8'd176,8'd194} : s = 203;
	{8'd176,8'd195} : s = 363;
	{8'd176,8'd196} : s = 199;
	{8'd176,8'd197} : s = 359;
	{8'd176,8'd198} : s = 350;
	{8'd176,8'd199} : s = 477;
	{8'd176,8'd200} : s = 188;
	{8'd176,8'd201} : s = 349;
	{8'd176,8'd202} : s = 347;
	{8'd176,8'd203} : s = 475;
	{8'd176,8'd204} : s = 343;
	{8'd176,8'd205} : s = 471;
	{8'd176,8'd206} : s = 463;
	{8'd176,8'd207} : s = 509;
	{8'd176,8'd208} : s = 3;
	{8'd176,8'd209} : s = 22;
	{8'd176,8'd210} : s = 21;
	{8'd176,8'd211} : s = 85;
	{8'd176,8'd212} : s = 19;
	{8'd176,8'd213} : s = 83;
	{8'd176,8'd214} : s = 78;
	{8'd176,8'd215} : s = 186;
	{8'd176,8'd216} : s = 14;
	{8'd176,8'd217} : s = 77;
	{8'd176,8'd218} : s = 75;
	{8'd176,8'd219} : s = 185;
	{8'd176,8'd220} : s = 71;
	{8'd176,8'd221} : s = 182;
	{8'd176,8'd222} : s = 181;
	{8'd176,8'd223} : s = 335;
	{8'd176,8'd224} : s = 13;
	{8'd176,8'd225} : s = 60;
	{8'd176,8'd226} : s = 58;
	{8'd176,8'd227} : s = 179;
	{8'd176,8'd228} : s = 57;
	{8'd176,8'd229} : s = 174;
	{8'd176,8'd230} : s = 173;
	{8'd176,8'd231} : s = 318;
	{8'd176,8'd232} : s = 54;
	{8'd176,8'd233} : s = 171;
	{8'd176,8'd234} : s = 167;
	{8'd176,8'd235} : s = 317;
	{8'd176,8'd236} : s = 158;
	{8'd176,8'd237} : s = 315;
	{8'd176,8'd238} : s = 311;
	{8'd176,8'd239} : s = 446;
	{8'd176,8'd240} : s = 11;
	{8'd176,8'd241} : s = 53;
	{8'd176,8'd242} : s = 51;
	{8'd176,8'd243} : s = 157;
	{8'd176,8'd244} : s = 46;
	{8'd176,8'd245} : s = 155;
	{8'd176,8'd246} : s = 151;
	{8'd176,8'd247} : s = 303;
	{8'd176,8'd248} : s = 45;
	{8'd176,8'd249} : s = 143;
	{8'd176,8'd250} : s = 124;
	{8'd176,8'd251} : s = 287;
	{8'd176,8'd252} : s = 122;
	{8'd176,8'd253} : s = 252;
	{8'd176,8'd254} : s = 250;
	{8'd176,8'd255} : s = 445;
	{8'd177,8'd0} : s = 275;
	{8'd177,8'd1} : s = 270;
	{8'd177,8'd2} : s = 403;
	{8'd177,8'd3} : s = 269;
	{8'd177,8'd4} : s = 398;
	{8'd177,8'd5} : s = 397;
	{8'd177,8'd6} : s = 483;
	{8'd177,8'd7} : s = 267;
	{8'd177,8'd8} : s = 395;
	{8'd177,8'd9} : s = 391;
	{8'd177,8'd10} : s = 476;
	{8'd177,8'd11} : s = 376;
	{8'd177,8'd12} : s = 474;
	{8'd177,8'd13} : s = 473;
	{8'd177,8'd14} : s = 506;
	{8'd177,8'd15} : s = 20;
	{8'd177,8'd16} : s = 104;
	{8'd177,8'd17} : s = 100;
	{8'd177,8'd18} : s = 263;
	{8'd177,8'd19} : s = 98;
	{8'd177,8'd20} : s = 240;
	{8'd177,8'd21} : s = 232;
	{8'd177,8'd22} : s = 372;
	{8'd177,8'd23} : s = 97;
	{8'd177,8'd24} : s = 228;
	{8'd177,8'd25} : s = 226;
	{8'd177,8'd26} : s = 370;
	{8'd177,8'd27} : s = 225;
	{8'd177,8'd28} : s = 369;
	{8'd177,8'd29} : s = 364;
	{8'd177,8'd30} : s = 470;
	{8'd177,8'd31} : s = 88;
	{8'd177,8'd32} : s = 216;
	{8'd177,8'd33} : s = 212;
	{8'd177,8'd34} : s = 362;
	{8'd177,8'd35} : s = 210;
	{8'd177,8'd36} : s = 361;
	{8'd177,8'd37} : s = 358;
	{8'd177,8'd38} : s = 469;
	{8'd177,8'd39} : s = 209;
	{8'd177,8'd40} : s = 357;
	{8'd177,8'd41} : s = 355;
	{8'd177,8'd42} : s = 467;
	{8'd177,8'd43} : s = 348;
	{8'd177,8'd44} : s = 462;
	{8'd177,8'd45} : s = 461;
	{8'd177,8'd46} : s = 505;
	{8'd177,8'd47} : s = 84;
	{8'd177,8'd48} : s = 204;
	{8'd177,8'd49} : s = 202;
	{8'd177,8'd50} : s = 346;
	{8'd177,8'd51} : s = 201;
	{8'd177,8'd52} : s = 345;
	{8'd177,8'd53} : s = 342;
	{8'd177,8'd54} : s = 459;
	{8'd177,8'd55} : s = 198;
	{8'd177,8'd56} : s = 341;
	{8'd177,8'd57} : s = 339;
	{8'd177,8'd58} : s = 455;
	{8'd177,8'd59} : s = 334;
	{8'd177,8'd60} : s = 444;
	{8'd177,8'd61} : s = 442;
	{8'd177,8'd62} : s = 502;
	{8'd177,8'd63} : s = 197;
	{8'd177,8'd64} : s = 333;
	{8'd177,8'd65} : s = 331;
	{8'd177,8'd66} : s = 441;
	{8'd177,8'd67} : s = 327;
	{8'd177,8'd68} : s = 438;
	{8'd177,8'd69} : s = 437;
	{8'd177,8'd70} : s = 501;
	{8'd177,8'd71} : s = 316;
	{8'd177,8'd72} : s = 435;
	{8'd177,8'd73} : s = 430;
	{8'd177,8'd74} : s = 499;
	{8'd177,8'd75} : s = 429;
	{8'd177,8'd76} : s = 494;
	{8'd177,8'd77} : s = 493;
	{8'd177,8'd78} : s = 510;
	{8'd177,8'd79} : s = 1;
	{8'd177,8'd80} : s = 18;
	{8'd177,8'd81} : s = 17;
	{8'd177,8'd82} : s = 82;
	{8'd177,8'd83} : s = 12;
	{8'd177,8'd84} : s = 81;
	{8'd177,8'd85} : s = 76;
	{8'd177,8'd86} : s = 195;
	{8'd177,8'd87} : s = 10;
	{8'd177,8'd88} : s = 74;
	{8'd177,8'd89} : s = 73;
	{8'd177,8'd90} : s = 184;
	{8'd177,8'd91} : s = 70;
	{8'd177,8'd92} : s = 180;
	{8'd177,8'd93} : s = 178;
	{8'd177,8'd94} : s = 314;
	{8'd177,8'd95} : s = 9;
	{8'd177,8'd96} : s = 69;
	{8'd177,8'd97} : s = 67;
	{8'd177,8'd98} : s = 177;
	{8'd177,8'd99} : s = 56;
	{8'd177,8'd100} : s = 172;
	{8'd177,8'd101} : s = 170;
	{8'd177,8'd102} : s = 313;
	{8'd177,8'd103} : s = 52;
	{8'd177,8'd104} : s = 169;
	{8'd177,8'd105} : s = 166;
	{8'd177,8'd106} : s = 310;
	{8'd177,8'd107} : s = 165;
	{8'd177,8'd108} : s = 309;
	{8'd177,8'd109} : s = 307;
	{8'd177,8'd110} : s = 427;
	{8'd177,8'd111} : s = 6;
	{8'd177,8'd112} : s = 50;
	{8'd177,8'd113} : s = 49;
	{8'd177,8'd114} : s = 163;
	{8'd177,8'd115} : s = 44;
	{8'd177,8'd116} : s = 156;
	{8'd177,8'd117} : s = 154;
	{8'd177,8'd118} : s = 302;
	{8'd177,8'd119} : s = 42;
	{8'd177,8'd120} : s = 153;
	{8'd177,8'd121} : s = 150;
	{8'd177,8'd122} : s = 301;
	{8'd177,8'd123} : s = 149;
	{8'd177,8'd124} : s = 299;
	{8'd177,8'd125} : s = 295;
	{8'd177,8'd126} : s = 423;
	{8'd177,8'd127} : s = 41;
	{8'd177,8'd128} : s = 147;
	{8'd177,8'd129} : s = 142;
	{8'd177,8'd130} : s = 286;
	{8'd177,8'd131} : s = 141;
	{8'd177,8'd132} : s = 285;
	{8'd177,8'd133} : s = 283;
	{8'd177,8'd134} : s = 414;
	{8'd177,8'd135} : s = 139;
	{8'd177,8'd136} : s = 279;
	{8'd177,8'd137} : s = 271;
	{8'd177,8'd138} : s = 413;
	{8'd177,8'd139} : s = 248;
	{8'd177,8'd140} : s = 411;
	{8'd177,8'd141} : s = 407;
	{8'd177,8'd142} : s = 491;
	{8'd177,8'd143} : s = 5;
	{8'd177,8'd144} : s = 38;
	{8'd177,8'd145} : s = 37;
	{8'd177,8'd146} : s = 135;
	{8'd177,8'd147} : s = 35;
	{8'd177,8'd148} : s = 120;
	{8'd177,8'd149} : s = 116;
	{8'd177,8'd150} : s = 244;
	{8'd177,8'd151} : s = 28;
	{8'd177,8'd152} : s = 114;
	{8'd177,8'd153} : s = 113;
	{8'd177,8'd154} : s = 242;
	{8'd177,8'd155} : s = 108;
	{8'd177,8'd156} : s = 241;
	{8'd177,8'd157} : s = 236;
	{8'd177,8'd158} : s = 399;
	{8'd177,8'd159} : s = 26;
	{8'd177,8'd160} : s = 106;
	{8'd177,8'd161} : s = 105;
	{8'd177,8'd162} : s = 234;
	{8'd177,8'd163} : s = 102;
	{8'd177,8'd164} : s = 233;
	{8'd177,8'd165} : s = 230;
	{8'd177,8'd166} : s = 380;
	{8'd177,8'd167} : s = 101;
	{8'd177,8'd168} : s = 229;
	{8'd177,8'd169} : s = 227;
	{8'd177,8'd170} : s = 378;
	{8'd177,8'd171} : s = 220;
	{8'd177,8'd172} : s = 377;
	{8'd177,8'd173} : s = 374;
	{8'd177,8'd174} : s = 487;
	{8'd177,8'd175} : s = 25;
	{8'd177,8'd176} : s = 99;
	{8'd177,8'd177} : s = 92;
	{8'd177,8'd178} : s = 218;
	{8'd177,8'd179} : s = 90;
	{8'd177,8'd180} : s = 217;
	{8'd177,8'd181} : s = 214;
	{8'd177,8'd182} : s = 373;
	{8'd177,8'd183} : s = 89;
	{8'd177,8'd184} : s = 213;
	{8'd177,8'd185} : s = 211;
	{8'd177,8'd186} : s = 371;
	{8'd177,8'd187} : s = 206;
	{8'd177,8'd188} : s = 366;
	{8'd177,8'd189} : s = 365;
	{8'd177,8'd190} : s = 478;
	{8'd177,8'd191} : s = 86;
	{8'd177,8'd192} : s = 205;
	{8'd177,8'd193} : s = 203;
	{8'd177,8'd194} : s = 363;
	{8'd177,8'd195} : s = 199;
	{8'd177,8'd196} : s = 359;
	{8'd177,8'd197} : s = 350;
	{8'd177,8'd198} : s = 477;
	{8'd177,8'd199} : s = 188;
	{8'd177,8'd200} : s = 349;
	{8'd177,8'd201} : s = 347;
	{8'd177,8'd202} : s = 475;
	{8'd177,8'd203} : s = 343;
	{8'd177,8'd204} : s = 471;
	{8'd177,8'd205} : s = 463;
	{8'd177,8'd206} : s = 509;
	{8'd177,8'd207} : s = 3;
	{8'd177,8'd208} : s = 22;
	{8'd177,8'd209} : s = 21;
	{8'd177,8'd210} : s = 85;
	{8'd177,8'd211} : s = 19;
	{8'd177,8'd212} : s = 83;
	{8'd177,8'd213} : s = 78;
	{8'd177,8'd214} : s = 186;
	{8'd177,8'd215} : s = 14;
	{8'd177,8'd216} : s = 77;
	{8'd177,8'd217} : s = 75;
	{8'd177,8'd218} : s = 185;
	{8'd177,8'd219} : s = 71;
	{8'd177,8'd220} : s = 182;
	{8'd177,8'd221} : s = 181;
	{8'd177,8'd222} : s = 335;
	{8'd177,8'd223} : s = 13;
	{8'd177,8'd224} : s = 60;
	{8'd177,8'd225} : s = 58;
	{8'd177,8'd226} : s = 179;
	{8'd177,8'd227} : s = 57;
	{8'd177,8'd228} : s = 174;
	{8'd177,8'd229} : s = 173;
	{8'd177,8'd230} : s = 318;
	{8'd177,8'd231} : s = 54;
	{8'd177,8'd232} : s = 171;
	{8'd177,8'd233} : s = 167;
	{8'd177,8'd234} : s = 317;
	{8'd177,8'd235} : s = 158;
	{8'd177,8'd236} : s = 315;
	{8'd177,8'd237} : s = 311;
	{8'd177,8'd238} : s = 446;
	{8'd177,8'd239} : s = 11;
	{8'd177,8'd240} : s = 53;
	{8'd177,8'd241} : s = 51;
	{8'd177,8'd242} : s = 157;
	{8'd177,8'd243} : s = 46;
	{8'd177,8'd244} : s = 155;
	{8'd177,8'd245} : s = 151;
	{8'd177,8'd246} : s = 303;
	{8'd177,8'd247} : s = 45;
	{8'd177,8'd248} : s = 143;
	{8'd177,8'd249} : s = 124;
	{8'd177,8'd250} : s = 287;
	{8'd177,8'd251} : s = 122;
	{8'd177,8'd252} : s = 252;
	{8'd177,8'd253} : s = 250;
	{8'd177,8'd254} : s = 445;
	{8'd177,8'd255} : s = 43;
	{8'd178,8'd0} : s = 270;
	{8'd178,8'd1} : s = 403;
	{8'd178,8'd2} : s = 269;
	{8'd178,8'd3} : s = 398;
	{8'd178,8'd4} : s = 397;
	{8'd178,8'd5} : s = 483;
	{8'd178,8'd6} : s = 267;
	{8'd178,8'd7} : s = 395;
	{8'd178,8'd8} : s = 391;
	{8'd178,8'd9} : s = 476;
	{8'd178,8'd10} : s = 376;
	{8'd178,8'd11} : s = 474;
	{8'd178,8'd12} : s = 473;
	{8'd178,8'd13} : s = 506;
	{8'd178,8'd14} : s = 20;
	{8'd178,8'd15} : s = 104;
	{8'd178,8'd16} : s = 100;
	{8'd178,8'd17} : s = 263;
	{8'd178,8'd18} : s = 98;
	{8'd178,8'd19} : s = 240;
	{8'd178,8'd20} : s = 232;
	{8'd178,8'd21} : s = 372;
	{8'd178,8'd22} : s = 97;
	{8'd178,8'd23} : s = 228;
	{8'd178,8'd24} : s = 226;
	{8'd178,8'd25} : s = 370;
	{8'd178,8'd26} : s = 225;
	{8'd178,8'd27} : s = 369;
	{8'd178,8'd28} : s = 364;
	{8'd178,8'd29} : s = 470;
	{8'd178,8'd30} : s = 88;
	{8'd178,8'd31} : s = 216;
	{8'd178,8'd32} : s = 212;
	{8'd178,8'd33} : s = 362;
	{8'd178,8'd34} : s = 210;
	{8'd178,8'd35} : s = 361;
	{8'd178,8'd36} : s = 358;
	{8'd178,8'd37} : s = 469;
	{8'd178,8'd38} : s = 209;
	{8'd178,8'd39} : s = 357;
	{8'd178,8'd40} : s = 355;
	{8'd178,8'd41} : s = 467;
	{8'd178,8'd42} : s = 348;
	{8'd178,8'd43} : s = 462;
	{8'd178,8'd44} : s = 461;
	{8'd178,8'd45} : s = 505;
	{8'd178,8'd46} : s = 84;
	{8'd178,8'd47} : s = 204;
	{8'd178,8'd48} : s = 202;
	{8'd178,8'd49} : s = 346;
	{8'd178,8'd50} : s = 201;
	{8'd178,8'd51} : s = 345;
	{8'd178,8'd52} : s = 342;
	{8'd178,8'd53} : s = 459;
	{8'd178,8'd54} : s = 198;
	{8'd178,8'd55} : s = 341;
	{8'd178,8'd56} : s = 339;
	{8'd178,8'd57} : s = 455;
	{8'd178,8'd58} : s = 334;
	{8'd178,8'd59} : s = 444;
	{8'd178,8'd60} : s = 442;
	{8'd178,8'd61} : s = 502;
	{8'd178,8'd62} : s = 197;
	{8'd178,8'd63} : s = 333;
	{8'd178,8'd64} : s = 331;
	{8'd178,8'd65} : s = 441;
	{8'd178,8'd66} : s = 327;
	{8'd178,8'd67} : s = 438;
	{8'd178,8'd68} : s = 437;
	{8'd178,8'd69} : s = 501;
	{8'd178,8'd70} : s = 316;
	{8'd178,8'd71} : s = 435;
	{8'd178,8'd72} : s = 430;
	{8'd178,8'd73} : s = 499;
	{8'd178,8'd74} : s = 429;
	{8'd178,8'd75} : s = 494;
	{8'd178,8'd76} : s = 493;
	{8'd178,8'd77} : s = 510;
	{8'd178,8'd78} : s = 1;
	{8'd178,8'd79} : s = 18;
	{8'd178,8'd80} : s = 17;
	{8'd178,8'd81} : s = 82;
	{8'd178,8'd82} : s = 12;
	{8'd178,8'd83} : s = 81;
	{8'd178,8'd84} : s = 76;
	{8'd178,8'd85} : s = 195;
	{8'd178,8'd86} : s = 10;
	{8'd178,8'd87} : s = 74;
	{8'd178,8'd88} : s = 73;
	{8'd178,8'd89} : s = 184;
	{8'd178,8'd90} : s = 70;
	{8'd178,8'd91} : s = 180;
	{8'd178,8'd92} : s = 178;
	{8'd178,8'd93} : s = 314;
	{8'd178,8'd94} : s = 9;
	{8'd178,8'd95} : s = 69;
	{8'd178,8'd96} : s = 67;
	{8'd178,8'd97} : s = 177;
	{8'd178,8'd98} : s = 56;
	{8'd178,8'd99} : s = 172;
	{8'd178,8'd100} : s = 170;
	{8'd178,8'd101} : s = 313;
	{8'd178,8'd102} : s = 52;
	{8'd178,8'd103} : s = 169;
	{8'd178,8'd104} : s = 166;
	{8'd178,8'd105} : s = 310;
	{8'd178,8'd106} : s = 165;
	{8'd178,8'd107} : s = 309;
	{8'd178,8'd108} : s = 307;
	{8'd178,8'd109} : s = 427;
	{8'd178,8'd110} : s = 6;
	{8'd178,8'd111} : s = 50;
	{8'd178,8'd112} : s = 49;
	{8'd178,8'd113} : s = 163;
	{8'd178,8'd114} : s = 44;
	{8'd178,8'd115} : s = 156;
	{8'd178,8'd116} : s = 154;
	{8'd178,8'd117} : s = 302;
	{8'd178,8'd118} : s = 42;
	{8'd178,8'd119} : s = 153;
	{8'd178,8'd120} : s = 150;
	{8'd178,8'd121} : s = 301;
	{8'd178,8'd122} : s = 149;
	{8'd178,8'd123} : s = 299;
	{8'd178,8'd124} : s = 295;
	{8'd178,8'd125} : s = 423;
	{8'd178,8'd126} : s = 41;
	{8'd178,8'd127} : s = 147;
	{8'd178,8'd128} : s = 142;
	{8'd178,8'd129} : s = 286;
	{8'd178,8'd130} : s = 141;
	{8'd178,8'd131} : s = 285;
	{8'd178,8'd132} : s = 283;
	{8'd178,8'd133} : s = 414;
	{8'd178,8'd134} : s = 139;
	{8'd178,8'd135} : s = 279;
	{8'd178,8'd136} : s = 271;
	{8'd178,8'd137} : s = 413;
	{8'd178,8'd138} : s = 248;
	{8'd178,8'd139} : s = 411;
	{8'd178,8'd140} : s = 407;
	{8'd178,8'd141} : s = 491;
	{8'd178,8'd142} : s = 5;
	{8'd178,8'd143} : s = 38;
	{8'd178,8'd144} : s = 37;
	{8'd178,8'd145} : s = 135;
	{8'd178,8'd146} : s = 35;
	{8'd178,8'd147} : s = 120;
	{8'd178,8'd148} : s = 116;
	{8'd178,8'd149} : s = 244;
	{8'd178,8'd150} : s = 28;
	{8'd178,8'd151} : s = 114;
	{8'd178,8'd152} : s = 113;
	{8'd178,8'd153} : s = 242;
	{8'd178,8'd154} : s = 108;
	{8'd178,8'd155} : s = 241;
	{8'd178,8'd156} : s = 236;
	{8'd178,8'd157} : s = 399;
	{8'd178,8'd158} : s = 26;
	{8'd178,8'd159} : s = 106;
	{8'd178,8'd160} : s = 105;
	{8'd178,8'd161} : s = 234;
	{8'd178,8'd162} : s = 102;
	{8'd178,8'd163} : s = 233;
	{8'd178,8'd164} : s = 230;
	{8'd178,8'd165} : s = 380;
	{8'd178,8'd166} : s = 101;
	{8'd178,8'd167} : s = 229;
	{8'd178,8'd168} : s = 227;
	{8'd178,8'd169} : s = 378;
	{8'd178,8'd170} : s = 220;
	{8'd178,8'd171} : s = 377;
	{8'd178,8'd172} : s = 374;
	{8'd178,8'd173} : s = 487;
	{8'd178,8'd174} : s = 25;
	{8'd178,8'd175} : s = 99;
	{8'd178,8'd176} : s = 92;
	{8'd178,8'd177} : s = 218;
	{8'd178,8'd178} : s = 90;
	{8'd178,8'd179} : s = 217;
	{8'd178,8'd180} : s = 214;
	{8'd178,8'd181} : s = 373;
	{8'd178,8'd182} : s = 89;
	{8'd178,8'd183} : s = 213;
	{8'd178,8'd184} : s = 211;
	{8'd178,8'd185} : s = 371;
	{8'd178,8'd186} : s = 206;
	{8'd178,8'd187} : s = 366;
	{8'd178,8'd188} : s = 365;
	{8'd178,8'd189} : s = 478;
	{8'd178,8'd190} : s = 86;
	{8'd178,8'd191} : s = 205;
	{8'd178,8'd192} : s = 203;
	{8'd178,8'd193} : s = 363;
	{8'd178,8'd194} : s = 199;
	{8'd178,8'd195} : s = 359;
	{8'd178,8'd196} : s = 350;
	{8'd178,8'd197} : s = 477;
	{8'd178,8'd198} : s = 188;
	{8'd178,8'd199} : s = 349;
	{8'd178,8'd200} : s = 347;
	{8'd178,8'd201} : s = 475;
	{8'd178,8'd202} : s = 343;
	{8'd178,8'd203} : s = 471;
	{8'd178,8'd204} : s = 463;
	{8'd178,8'd205} : s = 509;
	{8'd178,8'd206} : s = 3;
	{8'd178,8'd207} : s = 22;
	{8'd178,8'd208} : s = 21;
	{8'd178,8'd209} : s = 85;
	{8'd178,8'd210} : s = 19;
	{8'd178,8'd211} : s = 83;
	{8'd178,8'd212} : s = 78;
	{8'd178,8'd213} : s = 186;
	{8'd178,8'd214} : s = 14;
	{8'd178,8'd215} : s = 77;
	{8'd178,8'd216} : s = 75;
	{8'd178,8'd217} : s = 185;
	{8'd178,8'd218} : s = 71;
	{8'd178,8'd219} : s = 182;
	{8'd178,8'd220} : s = 181;
	{8'd178,8'd221} : s = 335;
	{8'd178,8'd222} : s = 13;
	{8'd178,8'd223} : s = 60;
	{8'd178,8'd224} : s = 58;
	{8'd178,8'd225} : s = 179;
	{8'd178,8'd226} : s = 57;
	{8'd178,8'd227} : s = 174;
	{8'd178,8'd228} : s = 173;
	{8'd178,8'd229} : s = 318;
	{8'd178,8'd230} : s = 54;
	{8'd178,8'd231} : s = 171;
	{8'd178,8'd232} : s = 167;
	{8'd178,8'd233} : s = 317;
	{8'd178,8'd234} : s = 158;
	{8'd178,8'd235} : s = 315;
	{8'd178,8'd236} : s = 311;
	{8'd178,8'd237} : s = 446;
	{8'd178,8'd238} : s = 11;
	{8'd178,8'd239} : s = 53;
	{8'd178,8'd240} : s = 51;
	{8'd178,8'd241} : s = 157;
	{8'd178,8'd242} : s = 46;
	{8'd178,8'd243} : s = 155;
	{8'd178,8'd244} : s = 151;
	{8'd178,8'd245} : s = 303;
	{8'd178,8'd246} : s = 45;
	{8'd178,8'd247} : s = 143;
	{8'd178,8'd248} : s = 124;
	{8'd178,8'd249} : s = 287;
	{8'd178,8'd250} : s = 122;
	{8'd178,8'd251} : s = 252;
	{8'd178,8'd252} : s = 250;
	{8'd178,8'd253} : s = 445;
	{8'd178,8'd254} : s = 43;
	{8'd178,8'd255} : s = 121;
	{8'd179,8'd0} : s = 403;
	{8'd179,8'd1} : s = 269;
	{8'd179,8'd2} : s = 398;
	{8'd179,8'd3} : s = 397;
	{8'd179,8'd4} : s = 483;
	{8'd179,8'd5} : s = 267;
	{8'd179,8'd6} : s = 395;
	{8'd179,8'd7} : s = 391;
	{8'd179,8'd8} : s = 476;
	{8'd179,8'd9} : s = 376;
	{8'd179,8'd10} : s = 474;
	{8'd179,8'd11} : s = 473;
	{8'd179,8'd12} : s = 506;
	{8'd179,8'd13} : s = 20;
	{8'd179,8'd14} : s = 104;
	{8'd179,8'd15} : s = 100;
	{8'd179,8'd16} : s = 263;
	{8'd179,8'd17} : s = 98;
	{8'd179,8'd18} : s = 240;
	{8'd179,8'd19} : s = 232;
	{8'd179,8'd20} : s = 372;
	{8'd179,8'd21} : s = 97;
	{8'd179,8'd22} : s = 228;
	{8'd179,8'd23} : s = 226;
	{8'd179,8'd24} : s = 370;
	{8'd179,8'd25} : s = 225;
	{8'd179,8'd26} : s = 369;
	{8'd179,8'd27} : s = 364;
	{8'd179,8'd28} : s = 470;
	{8'd179,8'd29} : s = 88;
	{8'd179,8'd30} : s = 216;
	{8'd179,8'd31} : s = 212;
	{8'd179,8'd32} : s = 362;
	{8'd179,8'd33} : s = 210;
	{8'd179,8'd34} : s = 361;
	{8'd179,8'd35} : s = 358;
	{8'd179,8'd36} : s = 469;
	{8'd179,8'd37} : s = 209;
	{8'd179,8'd38} : s = 357;
	{8'd179,8'd39} : s = 355;
	{8'd179,8'd40} : s = 467;
	{8'd179,8'd41} : s = 348;
	{8'd179,8'd42} : s = 462;
	{8'd179,8'd43} : s = 461;
	{8'd179,8'd44} : s = 505;
	{8'd179,8'd45} : s = 84;
	{8'd179,8'd46} : s = 204;
	{8'd179,8'd47} : s = 202;
	{8'd179,8'd48} : s = 346;
	{8'd179,8'd49} : s = 201;
	{8'd179,8'd50} : s = 345;
	{8'd179,8'd51} : s = 342;
	{8'd179,8'd52} : s = 459;
	{8'd179,8'd53} : s = 198;
	{8'd179,8'd54} : s = 341;
	{8'd179,8'd55} : s = 339;
	{8'd179,8'd56} : s = 455;
	{8'd179,8'd57} : s = 334;
	{8'd179,8'd58} : s = 444;
	{8'd179,8'd59} : s = 442;
	{8'd179,8'd60} : s = 502;
	{8'd179,8'd61} : s = 197;
	{8'd179,8'd62} : s = 333;
	{8'd179,8'd63} : s = 331;
	{8'd179,8'd64} : s = 441;
	{8'd179,8'd65} : s = 327;
	{8'd179,8'd66} : s = 438;
	{8'd179,8'd67} : s = 437;
	{8'd179,8'd68} : s = 501;
	{8'd179,8'd69} : s = 316;
	{8'd179,8'd70} : s = 435;
	{8'd179,8'd71} : s = 430;
	{8'd179,8'd72} : s = 499;
	{8'd179,8'd73} : s = 429;
	{8'd179,8'd74} : s = 494;
	{8'd179,8'd75} : s = 493;
	{8'd179,8'd76} : s = 510;
	{8'd179,8'd77} : s = 1;
	{8'd179,8'd78} : s = 18;
	{8'd179,8'd79} : s = 17;
	{8'd179,8'd80} : s = 82;
	{8'd179,8'd81} : s = 12;
	{8'd179,8'd82} : s = 81;
	{8'd179,8'd83} : s = 76;
	{8'd179,8'd84} : s = 195;
	{8'd179,8'd85} : s = 10;
	{8'd179,8'd86} : s = 74;
	{8'd179,8'd87} : s = 73;
	{8'd179,8'd88} : s = 184;
	{8'd179,8'd89} : s = 70;
	{8'd179,8'd90} : s = 180;
	{8'd179,8'd91} : s = 178;
	{8'd179,8'd92} : s = 314;
	{8'd179,8'd93} : s = 9;
	{8'd179,8'd94} : s = 69;
	{8'd179,8'd95} : s = 67;
	{8'd179,8'd96} : s = 177;
	{8'd179,8'd97} : s = 56;
	{8'd179,8'd98} : s = 172;
	{8'd179,8'd99} : s = 170;
	{8'd179,8'd100} : s = 313;
	{8'd179,8'd101} : s = 52;
	{8'd179,8'd102} : s = 169;
	{8'd179,8'd103} : s = 166;
	{8'd179,8'd104} : s = 310;
	{8'd179,8'd105} : s = 165;
	{8'd179,8'd106} : s = 309;
	{8'd179,8'd107} : s = 307;
	{8'd179,8'd108} : s = 427;
	{8'd179,8'd109} : s = 6;
	{8'd179,8'd110} : s = 50;
	{8'd179,8'd111} : s = 49;
	{8'd179,8'd112} : s = 163;
	{8'd179,8'd113} : s = 44;
	{8'd179,8'd114} : s = 156;
	{8'd179,8'd115} : s = 154;
	{8'd179,8'd116} : s = 302;
	{8'd179,8'd117} : s = 42;
	{8'd179,8'd118} : s = 153;
	{8'd179,8'd119} : s = 150;
	{8'd179,8'd120} : s = 301;
	{8'd179,8'd121} : s = 149;
	{8'd179,8'd122} : s = 299;
	{8'd179,8'd123} : s = 295;
	{8'd179,8'd124} : s = 423;
	{8'd179,8'd125} : s = 41;
	{8'd179,8'd126} : s = 147;
	{8'd179,8'd127} : s = 142;
	{8'd179,8'd128} : s = 286;
	{8'd179,8'd129} : s = 141;
	{8'd179,8'd130} : s = 285;
	{8'd179,8'd131} : s = 283;
	{8'd179,8'd132} : s = 414;
	{8'd179,8'd133} : s = 139;
	{8'd179,8'd134} : s = 279;
	{8'd179,8'd135} : s = 271;
	{8'd179,8'd136} : s = 413;
	{8'd179,8'd137} : s = 248;
	{8'd179,8'd138} : s = 411;
	{8'd179,8'd139} : s = 407;
	{8'd179,8'd140} : s = 491;
	{8'd179,8'd141} : s = 5;
	{8'd179,8'd142} : s = 38;
	{8'd179,8'd143} : s = 37;
	{8'd179,8'd144} : s = 135;
	{8'd179,8'd145} : s = 35;
	{8'd179,8'd146} : s = 120;
	{8'd179,8'd147} : s = 116;
	{8'd179,8'd148} : s = 244;
	{8'd179,8'd149} : s = 28;
	{8'd179,8'd150} : s = 114;
	{8'd179,8'd151} : s = 113;
	{8'd179,8'd152} : s = 242;
	{8'd179,8'd153} : s = 108;
	{8'd179,8'd154} : s = 241;
	{8'd179,8'd155} : s = 236;
	{8'd179,8'd156} : s = 399;
	{8'd179,8'd157} : s = 26;
	{8'd179,8'd158} : s = 106;
	{8'd179,8'd159} : s = 105;
	{8'd179,8'd160} : s = 234;
	{8'd179,8'd161} : s = 102;
	{8'd179,8'd162} : s = 233;
	{8'd179,8'd163} : s = 230;
	{8'd179,8'd164} : s = 380;
	{8'd179,8'd165} : s = 101;
	{8'd179,8'd166} : s = 229;
	{8'd179,8'd167} : s = 227;
	{8'd179,8'd168} : s = 378;
	{8'd179,8'd169} : s = 220;
	{8'd179,8'd170} : s = 377;
	{8'd179,8'd171} : s = 374;
	{8'd179,8'd172} : s = 487;
	{8'd179,8'd173} : s = 25;
	{8'd179,8'd174} : s = 99;
	{8'd179,8'd175} : s = 92;
	{8'd179,8'd176} : s = 218;
	{8'd179,8'd177} : s = 90;
	{8'd179,8'd178} : s = 217;
	{8'd179,8'd179} : s = 214;
	{8'd179,8'd180} : s = 373;
	{8'd179,8'd181} : s = 89;
	{8'd179,8'd182} : s = 213;
	{8'd179,8'd183} : s = 211;
	{8'd179,8'd184} : s = 371;
	{8'd179,8'd185} : s = 206;
	{8'd179,8'd186} : s = 366;
	{8'd179,8'd187} : s = 365;
	{8'd179,8'd188} : s = 478;
	{8'd179,8'd189} : s = 86;
	{8'd179,8'd190} : s = 205;
	{8'd179,8'd191} : s = 203;
	{8'd179,8'd192} : s = 363;
	{8'd179,8'd193} : s = 199;
	{8'd179,8'd194} : s = 359;
	{8'd179,8'd195} : s = 350;
	{8'd179,8'd196} : s = 477;
	{8'd179,8'd197} : s = 188;
	{8'd179,8'd198} : s = 349;
	{8'd179,8'd199} : s = 347;
	{8'd179,8'd200} : s = 475;
	{8'd179,8'd201} : s = 343;
	{8'd179,8'd202} : s = 471;
	{8'd179,8'd203} : s = 463;
	{8'd179,8'd204} : s = 509;
	{8'd179,8'd205} : s = 3;
	{8'd179,8'd206} : s = 22;
	{8'd179,8'd207} : s = 21;
	{8'd179,8'd208} : s = 85;
	{8'd179,8'd209} : s = 19;
	{8'd179,8'd210} : s = 83;
	{8'd179,8'd211} : s = 78;
	{8'd179,8'd212} : s = 186;
	{8'd179,8'd213} : s = 14;
	{8'd179,8'd214} : s = 77;
	{8'd179,8'd215} : s = 75;
	{8'd179,8'd216} : s = 185;
	{8'd179,8'd217} : s = 71;
	{8'd179,8'd218} : s = 182;
	{8'd179,8'd219} : s = 181;
	{8'd179,8'd220} : s = 335;
	{8'd179,8'd221} : s = 13;
	{8'd179,8'd222} : s = 60;
	{8'd179,8'd223} : s = 58;
	{8'd179,8'd224} : s = 179;
	{8'd179,8'd225} : s = 57;
	{8'd179,8'd226} : s = 174;
	{8'd179,8'd227} : s = 173;
	{8'd179,8'd228} : s = 318;
	{8'd179,8'd229} : s = 54;
	{8'd179,8'd230} : s = 171;
	{8'd179,8'd231} : s = 167;
	{8'd179,8'd232} : s = 317;
	{8'd179,8'd233} : s = 158;
	{8'd179,8'd234} : s = 315;
	{8'd179,8'd235} : s = 311;
	{8'd179,8'd236} : s = 446;
	{8'd179,8'd237} : s = 11;
	{8'd179,8'd238} : s = 53;
	{8'd179,8'd239} : s = 51;
	{8'd179,8'd240} : s = 157;
	{8'd179,8'd241} : s = 46;
	{8'd179,8'd242} : s = 155;
	{8'd179,8'd243} : s = 151;
	{8'd179,8'd244} : s = 303;
	{8'd179,8'd245} : s = 45;
	{8'd179,8'd246} : s = 143;
	{8'd179,8'd247} : s = 124;
	{8'd179,8'd248} : s = 287;
	{8'd179,8'd249} : s = 122;
	{8'd179,8'd250} : s = 252;
	{8'd179,8'd251} : s = 250;
	{8'd179,8'd252} : s = 445;
	{8'd179,8'd253} : s = 43;
	{8'd179,8'd254} : s = 121;
	{8'd179,8'd255} : s = 118;
	{8'd180,8'd0} : s = 269;
	{8'd180,8'd1} : s = 398;
	{8'd180,8'd2} : s = 397;
	{8'd180,8'd3} : s = 483;
	{8'd180,8'd4} : s = 267;
	{8'd180,8'd5} : s = 395;
	{8'd180,8'd6} : s = 391;
	{8'd180,8'd7} : s = 476;
	{8'd180,8'd8} : s = 376;
	{8'd180,8'd9} : s = 474;
	{8'd180,8'd10} : s = 473;
	{8'd180,8'd11} : s = 506;
	{8'd180,8'd12} : s = 20;
	{8'd180,8'd13} : s = 104;
	{8'd180,8'd14} : s = 100;
	{8'd180,8'd15} : s = 263;
	{8'd180,8'd16} : s = 98;
	{8'd180,8'd17} : s = 240;
	{8'd180,8'd18} : s = 232;
	{8'd180,8'd19} : s = 372;
	{8'd180,8'd20} : s = 97;
	{8'd180,8'd21} : s = 228;
	{8'd180,8'd22} : s = 226;
	{8'd180,8'd23} : s = 370;
	{8'd180,8'd24} : s = 225;
	{8'd180,8'd25} : s = 369;
	{8'd180,8'd26} : s = 364;
	{8'd180,8'd27} : s = 470;
	{8'd180,8'd28} : s = 88;
	{8'd180,8'd29} : s = 216;
	{8'd180,8'd30} : s = 212;
	{8'd180,8'd31} : s = 362;
	{8'd180,8'd32} : s = 210;
	{8'd180,8'd33} : s = 361;
	{8'd180,8'd34} : s = 358;
	{8'd180,8'd35} : s = 469;
	{8'd180,8'd36} : s = 209;
	{8'd180,8'd37} : s = 357;
	{8'd180,8'd38} : s = 355;
	{8'd180,8'd39} : s = 467;
	{8'd180,8'd40} : s = 348;
	{8'd180,8'd41} : s = 462;
	{8'd180,8'd42} : s = 461;
	{8'd180,8'd43} : s = 505;
	{8'd180,8'd44} : s = 84;
	{8'd180,8'd45} : s = 204;
	{8'd180,8'd46} : s = 202;
	{8'd180,8'd47} : s = 346;
	{8'd180,8'd48} : s = 201;
	{8'd180,8'd49} : s = 345;
	{8'd180,8'd50} : s = 342;
	{8'd180,8'd51} : s = 459;
	{8'd180,8'd52} : s = 198;
	{8'd180,8'd53} : s = 341;
	{8'd180,8'd54} : s = 339;
	{8'd180,8'd55} : s = 455;
	{8'd180,8'd56} : s = 334;
	{8'd180,8'd57} : s = 444;
	{8'd180,8'd58} : s = 442;
	{8'd180,8'd59} : s = 502;
	{8'd180,8'd60} : s = 197;
	{8'd180,8'd61} : s = 333;
	{8'd180,8'd62} : s = 331;
	{8'd180,8'd63} : s = 441;
	{8'd180,8'd64} : s = 327;
	{8'd180,8'd65} : s = 438;
	{8'd180,8'd66} : s = 437;
	{8'd180,8'd67} : s = 501;
	{8'd180,8'd68} : s = 316;
	{8'd180,8'd69} : s = 435;
	{8'd180,8'd70} : s = 430;
	{8'd180,8'd71} : s = 499;
	{8'd180,8'd72} : s = 429;
	{8'd180,8'd73} : s = 494;
	{8'd180,8'd74} : s = 493;
	{8'd180,8'd75} : s = 510;
	{8'd180,8'd76} : s = 1;
	{8'd180,8'd77} : s = 18;
	{8'd180,8'd78} : s = 17;
	{8'd180,8'd79} : s = 82;
	{8'd180,8'd80} : s = 12;
	{8'd180,8'd81} : s = 81;
	{8'd180,8'd82} : s = 76;
	{8'd180,8'd83} : s = 195;
	{8'd180,8'd84} : s = 10;
	{8'd180,8'd85} : s = 74;
	{8'd180,8'd86} : s = 73;
	{8'd180,8'd87} : s = 184;
	{8'd180,8'd88} : s = 70;
	{8'd180,8'd89} : s = 180;
	{8'd180,8'd90} : s = 178;
	{8'd180,8'd91} : s = 314;
	{8'd180,8'd92} : s = 9;
	{8'd180,8'd93} : s = 69;
	{8'd180,8'd94} : s = 67;
	{8'd180,8'd95} : s = 177;
	{8'd180,8'd96} : s = 56;
	{8'd180,8'd97} : s = 172;
	{8'd180,8'd98} : s = 170;
	{8'd180,8'd99} : s = 313;
	{8'd180,8'd100} : s = 52;
	{8'd180,8'd101} : s = 169;
	{8'd180,8'd102} : s = 166;
	{8'd180,8'd103} : s = 310;
	{8'd180,8'd104} : s = 165;
	{8'd180,8'd105} : s = 309;
	{8'd180,8'd106} : s = 307;
	{8'd180,8'd107} : s = 427;
	{8'd180,8'd108} : s = 6;
	{8'd180,8'd109} : s = 50;
	{8'd180,8'd110} : s = 49;
	{8'd180,8'd111} : s = 163;
	{8'd180,8'd112} : s = 44;
	{8'd180,8'd113} : s = 156;
	{8'd180,8'd114} : s = 154;
	{8'd180,8'd115} : s = 302;
	{8'd180,8'd116} : s = 42;
	{8'd180,8'd117} : s = 153;
	{8'd180,8'd118} : s = 150;
	{8'd180,8'd119} : s = 301;
	{8'd180,8'd120} : s = 149;
	{8'd180,8'd121} : s = 299;
	{8'd180,8'd122} : s = 295;
	{8'd180,8'd123} : s = 423;
	{8'd180,8'd124} : s = 41;
	{8'd180,8'd125} : s = 147;
	{8'd180,8'd126} : s = 142;
	{8'd180,8'd127} : s = 286;
	{8'd180,8'd128} : s = 141;
	{8'd180,8'd129} : s = 285;
	{8'd180,8'd130} : s = 283;
	{8'd180,8'd131} : s = 414;
	{8'd180,8'd132} : s = 139;
	{8'd180,8'd133} : s = 279;
	{8'd180,8'd134} : s = 271;
	{8'd180,8'd135} : s = 413;
	{8'd180,8'd136} : s = 248;
	{8'd180,8'd137} : s = 411;
	{8'd180,8'd138} : s = 407;
	{8'd180,8'd139} : s = 491;
	{8'd180,8'd140} : s = 5;
	{8'd180,8'd141} : s = 38;
	{8'd180,8'd142} : s = 37;
	{8'd180,8'd143} : s = 135;
	{8'd180,8'd144} : s = 35;
	{8'd180,8'd145} : s = 120;
	{8'd180,8'd146} : s = 116;
	{8'd180,8'd147} : s = 244;
	{8'd180,8'd148} : s = 28;
	{8'd180,8'd149} : s = 114;
	{8'd180,8'd150} : s = 113;
	{8'd180,8'd151} : s = 242;
	{8'd180,8'd152} : s = 108;
	{8'd180,8'd153} : s = 241;
	{8'd180,8'd154} : s = 236;
	{8'd180,8'd155} : s = 399;
	{8'd180,8'd156} : s = 26;
	{8'd180,8'd157} : s = 106;
	{8'd180,8'd158} : s = 105;
	{8'd180,8'd159} : s = 234;
	{8'd180,8'd160} : s = 102;
	{8'd180,8'd161} : s = 233;
	{8'd180,8'd162} : s = 230;
	{8'd180,8'd163} : s = 380;
	{8'd180,8'd164} : s = 101;
	{8'd180,8'd165} : s = 229;
	{8'd180,8'd166} : s = 227;
	{8'd180,8'd167} : s = 378;
	{8'd180,8'd168} : s = 220;
	{8'd180,8'd169} : s = 377;
	{8'd180,8'd170} : s = 374;
	{8'd180,8'd171} : s = 487;
	{8'd180,8'd172} : s = 25;
	{8'd180,8'd173} : s = 99;
	{8'd180,8'd174} : s = 92;
	{8'd180,8'd175} : s = 218;
	{8'd180,8'd176} : s = 90;
	{8'd180,8'd177} : s = 217;
	{8'd180,8'd178} : s = 214;
	{8'd180,8'd179} : s = 373;
	{8'd180,8'd180} : s = 89;
	{8'd180,8'd181} : s = 213;
	{8'd180,8'd182} : s = 211;
	{8'd180,8'd183} : s = 371;
	{8'd180,8'd184} : s = 206;
	{8'd180,8'd185} : s = 366;
	{8'd180,8'd186} : s = 365;
	{8'd180,8'd187} : s = 478;
	{8'd180,8'd188} : s = 86;
	{8'd180,8'd189} : s = 205;
	{8'd180,8'd190} : s = 203;
	{8'd180,8'd191} : s = 363;
	{8'd180,8'd192} : s = 199;
	{8'd180,8'd193} : s = 359;
	{8'd180,8'd194} : s = 350;
	{8'd180,8'd195} : s = 477;
	{8'd180,8'd196} : s = 188;
	{8'd180,8'd197} : s = 349;
	{8'd180,8'd198} : s = 347;
	{8'd180,8'd199} : s = 475;
	{8'd180,8'd200} : s = 343;
	{8'd180,8'd201} : s = 471;
	{8'd180,8'd202} : s = 463;
	{8'd180,8'd203} : s = 509;
	{8'd180,8'd204} : s = 3;
	{8'd180,8'd205} : s = 22;
	{8'd180,8'd206} : s = 21;
	{8'd180,8'd207} : s = 85;
	{8'd180,8'd208} : s = 19;
	{8'd180,8'd209} : s = 83;
	{8'd180,8'd210} : s = 78;
	{8'd180,8'd211} : s = 186;
	{8'd180,8'd212} : s = 14;
	{8'd180,8'd213} : s = 77;
	{8'd180,8'd214} : s = 75;
	{8'd180,8'd215} : s = 185;
	{8'd180,8'd216} : s = 71;
	{8'd180,8'd217} : s = 182;
	{8'd180,8'd218} : s = 181;
	{8'd180,8'd219} : s = 335;
	{8'd180,8'd220} : s = 13;
	{8'd180,8'd221} : s = 60;
	{8'd180,8'd222} : s = 58;
	{8'd180,8'd223} : s = 179;
	{8'd180,8'd224} : s = 57;
	{8'd180,8'd225} : s = 174;
	{8'd180,8'd226} : s = 173;
	{8'd180,8'd227} : s = 318;
	{8'd180,8'd228} : s = 54;
	{8'd180,8'd229} : s = 171;
	{8'd180,8'd230} : s = 167;
	{8'd180,8'd231} : s = 317;
	{8'd180,8'd232} : s = 158;
	{8'd180,8'd233} : s = 315;
	{8'd180,8'd234} : s = 311;
	{8'd180,8'd235} : s = 446;
	{8'd180,8'd236} : s = 11;
	{8'd180,8'd237} : s = 53;
	{8'd180,8'd238} : s = 51;
	{8'd180,8'd239} : s = 157;
	{8'd180,8'd240} : s = 46;
	{8'd180,8'd241} : s = 155;
	{8'd180,8'd242} : s = 151;
	{8'd180,8'd243} : s = 303;
	{8'd180,8'd244} : s = 45;
	{8'd180,8'd245} : s = 143;
	{8'd180,8'd246} : s = 124;
	{8'd180,8'd247} : s = 287;
	{8'd180,8'd248} : s = 122;
	{8'd180,8'd249} : s = 252;
	{8'd180,8'd250} : s = 250;
	{8'd180,8'd251} : s = 445;
	{8'd180,8'd252} : s = 43;
	{8'd180,8'd253} : s = 121;
	{8'd180,8'd254} : s = 118;
	{8'd180,8'd255} : s = 249;
	{8'd181,8'd0} : s = 398;
	{8'd181,8'd1} : s = 397;
	{8'd181,8'd2} : s = 483;
	{8'd181,8'd3} : s = 267;
	{8'd181,8'd4} : s = 395;
	{8'd181,8'd5} : s = 391;
	{8'd181,8'd6} : s = 476;
	{8'd181,8'd7} : s = 376;
	{8'd181,8'd8} : s = 474;
	{8'd181,8'd9} : s = 473;
	{8'd181,8'd10} : s = 506;
	{8'd181,8'd11} : s = 20;
	{8'd181,8'd12} : s = 104;
	{8'd181,8'd13} : s = 100;
	{8'd181,8'd14} : s = 263;
	{8'd181,8'd15} : s = 98;
	{8'd181,8'd16} : s = 240;
	{8'd181,8'd17} : s = 232;
	{8'd181,8'd18} : s = 372;
	{8'd181,8'd19} : s = 97;
	{8'd181,8'd20} : s = 228;
	{8'd181,8'd21} : s = 226;
	{8'd181,8'd22} : s = 370;
	{8'd181,8'd23} : s = 225;
	{8'd181,8'd24} : s = 369;
	{8'd181,8'd25} : s = 364;
	{8'd181,8'd26} : s = 470;
	{8'd181,8'd27} : s = 88;
	{8'd181,8'd28} : s = 216;
	{8'd181,8'd29} : s = 212;
	{8'd181,8'd30} : s = 362;
	{8'd181,8'd31} : s = 210;
	{8'd181,8'd32} : s = 361;
	{8'd181,8'd33} : s = 358;
	{8'd181,8'd34} : s = 469;
	{8'd181,8'd35} : s = 209;
	{8'd181,8'd36} : s = 357;
	{8'd181,8'd37} : s = 355;
	{8'd181,8'd38} : s = 467;
	{8'd181,8'd39} : s = 348;
	{8'd181,8'd40} : s = 462;
	{8'd181,8'd41} : s = 461;
	{8'd181,8'd42} : s = 505;
	{8'd181,8'd43} : s = 84;
	{8'd181,8'd44} : s = 204;
	{8'd181,8'd45} : s = 202;
	{8'd181,8'd46} : s = 346;
	{8'd181,8'd47} : s = 201;
	{8'd181,8'd48} : s = 345;
	{8'd181,8'd49} : s = 342;
	{8'd181,8'd50} : s = 459;
	{8'd181,8'd51} : s = 198;
	{8'd181,8'd52} : s = 341;
	{8'd181,8'd53} : s = 339;
	{8'd181,8'd54} : s = 455;
	{8'd181,8'd55} : s = 334;
	{8'd181,8'd56} : s = 444;
	{8'd181,8'd57} : s = 442;
	{8'd181,8'd58} : s = 502;
	{8'd181,8'd59} : s = 197;
	{8'd181,8'd60} : s = 333;
	{8'd181,8'd61} : s = 331;
	{8'd181,8'd62} : s = 441;
	{8'd181,8'd63} : s = 327;
	{8'd181,8'd64} : s = 438;
	{8'd181,8'd65} : s = 437;
	{8'd181,8'd66} : s = 501;
	{8'd181,8'd67} : s = 316;
	{8'd181,8'd68} : s = 435;
	{8'd181,8'd69} : s = 430;
	{8'd181,8'd70} : s = 499;
	{8'd181,8'd71} : s = 429;
	{8'd181,8'd72} : s = 494;
	{8'd181,8'd73} : s = 493;
	{8'd181,8'd74} : s = 510;
	{8'd181,8'd75} : s = 1;
	{8'd181,8'd76} : s = 18;
	{8'd181,8'd77} : s = 17;
	{8'd181,8'd78} : s = 82;
	{8'd181,8'd79} : s = 12;
	{8'd181,8'd80} : s = 81;
	{8'd181,8'd81} : s = 76;
	{8'd181,8'd82} : s = 195;
	{8'd181,8'd83} : s = 10;
	{8'd181,8'd84} : s = 74;
	{8'd181,8'd85} : s = 73;
	{8'd181,8'd86} : s = 184;
	{8'd181,8'd87} : s = 70;
	{8'd181,8'd88} : s = 180;
	{8'd181,8'd89} : s = 178;
	{8'd181,8'd90} : s = 314;
	{8'd181,8'd91} : s = 9;
	{8'd181,8'd92} : s = 69;
	{8'd181,8'd93} : s = 67;
	{8'd181,8'd94} : s = 177;
	{8'd181,8'd95} : s = 56;
	{8'd181,8'd96} : s = 172;
	{8'd181,8'd97} : s = 170;
	{8'd181,8'd98} : s = 313;
	{8'd181,8'd99} : s = 52;
	{8'd181,8'd100} : s = 169;
	{8'd181,8'd101} : s = 166;
	{8'd181,8'd102} : s = 310;
	{8'd181,8'd103} : s = 165;
	{8'd181,8'd104} : s = 309;
	{8'd181,8'd105} : s = 307;
	{8'd181,8'd106} : s = 427;
	{8'd181,8'd107} : s = 6;
	{8'd181,8'd108} : s = 50;
	{8'd181,8'd109} : s = 49;
	{8'd181,8'd110} : s = 163;
	{8'd181,8'd111} : s = 44;
	{8'd181,8'd112} : s = 156;
	{8'd181,8'd113} : s = 154;
	{8'd181,8'd114} : s = 302;
	{8'd181,8'd115} : s = 42;
	{8'd181,8'd116} : s = 153;
	{8'd181,8'd117} : s = 150;
	{8'd181,8'd118} : s = 301;
	{8'd181,8'd119} : s = 149;
	{8'd181,8'd120} : s = 299;
	{8'd181,8'd121} : s = 295;
	{8'd181,8'd122} : s = 423;
	{8'd181,8'd123} : s = 41;
	{8'd181,8'd124} : s = 147;
	{8'd181,8'd125} : s = 142;
	{8'd181,8'd126} : s = 286;
	{8'd181,8'd127} : s = 141;
	{8'd181,8'd128} : s = 285;
	{8'd181,8'd129} : s = 283;
	{8'd181,8'd130} : s = 414;
	{8'd181,8'd131} : s = 139;
	{8'd181,8'd132} : s = 279;
	{8'd181,8'd133} : s = 271;
	{8'd181,8'd134} : s = 413;
	{8'd181,8'd135} : s = 248;
	{8'd181,8'd136} : s = 411;
	{8'd181,8'd137} : s = 407;
	{8'd181,8'd138} : s = 491;
	{8'd181,8'd139} : s = 5;
	{8'd181,8'd140} : s = 38;
	{8'd181,8'd141} : s = 37;
	{8'd181,8'd142} : s = 135;
	{8'd181,8'd143} : s = 35;
	{8'd181,8'd144} : s = 120;
	{8'd181,8'd145} : s = 116;
	{8'd181,8'd146} : s = 244;
	{8'd181,8'd147} : s = 28;
	{8'd181,8'd148} : s = 114;
	{8'd181,8'd149} : s = 113;
	{8'd181,8'd150} : s = 242;
	{8'd181,8'd151} : s = 108;
	{8'd181,8'd152} : s = 241;
	{8'd181,8'd153} : s = 236;
	{8'd181,8'd154} : s = 399;
	{8'd181,8'd155} : s = 26;
	{8'd181,8'd156} : s = 106;
	{8'd181,8'd157} : s = 105;
	{8'd181,8'd158} : s = 234;
	{8'd181,8'd159} : s = 102;
	{8'd181,8'd160} : s = 233;
	{8'd181,8'd161} : s = 230;
	{8'd181,8'd162} : s = 380;
	{8'd181,8'd163} : s = 101;
	{8'd181,8'd164} : s = 229;
	{8'd181,8'd165} : s = 227;
	{8'd181,8'd166} : s = 378;
	{8'd181,8'd167} : s = 220;
	{8'd181,8'd168} : s = 377;
	{8'd181,8'd169} : s = 374;
	{8'd181,8'd170} : s = 487;
	{8'd181,8'd171} : s = 25;
	{8'd181,8'd172} : s = 99;
	{8'd181,8'd173} : s = 92;
	{8'd181,8'd174} : s = 218;
	{8'd181,8'd175} : s = 90;
	{8'd181,8'd176} : s = 217;
	{8'd181,8'd177} : s = 214;
	{8'd181,8'd178} : s = 373;
	{8'd181,8'd179} : s = 89;
	{8'd181,8'd180} : s = 213;
	{8'd181,8'd181} : s = 211;
	{8'd181,8'd182} : s = 371;
	{8'd181,8'd183} : s = 206;
	{8'd181,8'd184} : s = 366;
	{8'd181,8'd185} : s = 365;
	{8'd181,8'd186} : s = 478;
	{8'd181,8'd187} : s = 86;
	{8'd181,8'd188} : s = 205;
	{8'd181,8'd189} : s = 203;
	{8'd181,8'd190} : s = 363;
	{8'd181,8'd191} : s = 199;
	{8'd181,8'd192} : s = 359;
	{8'd181,8'd193} : s = 350;
	{8'd181,8'd194} : s = 477;
	{8'd181,8'd195} : s = 188;
	{8'd181,8'd196} : s = 349;
	{8'd181,8'd197} : s = 347;
	{8'd181,8'd198} : s = 475;
	{8'd181,8'd199} : s = 343;
	{8'd181,8'd200} : s = 471;
	{8'd181,8'd201} : s = 463;
	{8'd181,8'd202} : s = 509;
	{8'd181,8'd203} : s = 3;
	{8'd181,8'd204} : s = 22;
	{8'd181,8'd205} : s = 21;
	{8'd181,8'd206} : s = 85;
	{8'd181,8'd207} : s = 19;
	{8'd181,8'd208} : s = 83;
	{8'd181,8'd209} : s = 78;
	{8'd181,8'd210} : s = 186;
	{8'd181,8'd211} : s = 14;
	{8'd181,8'd212} : s = 77;
	{8'd181,8'd213} : s = 75;
	{8'd181,8'd214} : s = 185;
	{8'd181,8'd215} : s = 71;
	{8'd181,8'd216} : s = 182;
	{8'd181,8'd217} : s = 181;
	{8'd181,8'd218} : s = 335;
	{8'd181,8'd219} : s = 13;
	{8'd181,8'd220} : s = 60;
	{8'd181,8'd221} : s = 58;
	{8'd181,8'd222} : s = 179;
	{8'd181,8'd223} : s = 57;
	{8'd181,8'd224} : s = 174;
	{8'd181,8'd225} : s = 173;
	{8'd181,8'd226} : s = 318;
	{8'd181,8'd227} : s = 54;
	{8'd181,8'd228} : s = 171;
	{8'd181,8'd229} : s = 167;
	{8'd181,8'd230} : s = 317;
	{8'd181,8'd231} : s = 158;
	{8'd181,8'd232} : s = 315;
	{8'd181,8'd233} : s = 311;
	{8'd181,8'd234} : s = 446;
	{8'd181,8'd235} : s = 11;
	{8'd181,8'd236} : s = 53;
	{8'd181,8'd237} : s = 51;
	{8'd181,8'd238} : s = 157;
	{8'd181,8'd239} : s = 46;
	{8'd181,8'd240} : s = 155;
	{8'd181,8'd241} : s = 151;
	{8'd181,8'd242} : s = 303;
	{8'd181,8'd243} : s = 45;
	{8'd181,8'd244} : s = 143;
	{8'd181,8'd245} : s = 124;
	{8'd181,8'd246} : s = 287;
	{8'd181,8'd247} : s = 122;
	{8'd181,8'd248} : s = 252;
	{8'd181,8'd249} : s = 250;
	{8'd181,8'd250} : s = 445;
	{8'd181,8'd251} : s = 43;
	{8'd181,8'd252} : s = 121;
	{8'd181,8'd253} : s = 118;
	{8'd181,8'd254} : s = 249;
	{8'd181,8'd255} : s = 117;
	{8'd182,8'd0} : s = 397;
	{8'd182,8'd1} : s = 483;
	{8'd182,8'd2} : s = 267;
	{8'd182,8'd3} : s = 395;
	{8'd182,8'd4} : s = 391;
	{8'd182,8'd5} : s = 476;
	{8'd182,8'd6} : s = 376;
	{8'd182,8'd7} : s = 474;
	{8'd182,8'd8} : s = 473;
	{8'd182,8'd9} : s = 506;
	{8'd182,8'd10} : s = 20;
	{8'd182,8'd11} : s = 104;
	{8'd182,8'd12} : s = 100;
	{8'd182,8'd13} : s = 263;
	{8'd182,8'd14} : s = 98;
	{8'd182,8'd15} : s = 240;
	{8'd182,8'd16} : s = 232;
	{8'd182,8'd17} : s = 372;
	{8'd182,8'd18} : s = 97;
	{8'd182,8'd19} : s = 228;
	{8'd182,8'd20} : s = 226;
	{8'd182,8'd21} : s = 370;
	{8'd182,8'd22} : s = 225;
	{8'd182,8'd23} : s = 369;
	{8'd182,8'd24} : s = 364;
	{8'd182,8'd25} : s = 470;
	{8'd182,8'd26} : s = 88;
	{8'd182,8'd27} : s = 216;
	{8'd182,8'd28} : s = 212;
	{8'd182,8'd29} : s = 362;
	{8'd182,8'd30} : s = 210;
	{8'd182,8'd31} : s = 361;
	{8'd182,8'd32} : s = 358;
	{8'd182,8'd33} : s = 469;
	{8'd182,8'd34} : s = 209;
	{8'd182,8'd35} : s = 357;
	{8'd182,8'd36} : s = 355;
	{8'd182,8'd37} : s = 467;
	{8'd182,8'd38} : s = 348;
	{8'd182,8'd39} : s = 462;
	{8'd182,8'd40} : s = 461;
	{8'd182,8'd41} : s = 505;
	{8'd182,8'd42} : s = 84;
	{8'd182,8'd43} : s = 204;
	{8'd182,8'd44} : s = 202;
	{8'd182,8'd45} : s = 346;
	{8'd182,8'd46} : s = 201;
	{8'd182,8'd47} : s = 345;
	{8'd182,8'd48} : s = 342;
	{8'd182,8'd49} : s = 459;
	{8'd182,8'd50} : s = 198;
	{8'd182,8'd51} : s = 341;
	{8'd182,8'd52} : s = 339;
	{8'd182,8'd53} : s = 455;
	{8'd182,8'd54} : s = 334;
	{8'd182,8'd55} : s = 444;
	{8'd182,8'd56} : s = 442;
	{8'd182,8'd57} : s = 502;
	{8'd182,8'd58} : s = 197;
	{8'd182,8'd59} : s = 333;
	{8'd182,8'd60} : s = 331;
	{8'd182,8'd61} : s = 441;
	{8'd182,8'd62} : s = 327;
	{8'd182,8'd63} : s = 438;
	{8'd182,8'd64} : s = 437;
	{8'd182,8'd65} : s = 501;
	{8'd182,8'd66} : s = 316;
	{8'd182,8'd67} : s = 435;
	{8'd182,8'd68} : s = 430;
	{8'd182,8'd69} : s = 499;
	{8'd182,8'd70} : s = 429;
	{8'd182,8'd71} : s = 494;
	{8'd182,8'd72} : s = 493;
	{8'd182,8'd73} : s = 510;
	{8'd182,8'd74} : s = 1;
	{8'd182,8'd75} : s = 18;
	{8'd182,8'd76} : s = 17;
	{8'd182,8'd77} : s = 82;
	{8'd182,8'd78} : s = 12;
	{8'd182,8'd79} : s = 81;
	{8'd182,8'd80} : s = 76;
	{8'd182,8'd81} : s = 195;
	{8'd182,8'd82} : s = 10;
	{8'd182,8'd83} : s = 74;
	{8'd182,8'd84} : s = 73;
	{8'd182,8'd85} : s = 184;
	{8'd182,8'd86} : s = 70;
	{8'd182,8'd87} : s = 180;
	{8'd182,8'd88} : s = 178;
	{8'd182,8'd89} : s = 314;
	{8'd182,8'd90} : s = 9;
	{8'd182,8'd91} : s = 69;
	{8'd182,8'd92} : s = 67;
	{8'd182,8'd93} : s = 177;
	{8'd182,8'd94} : s = 56;
	{8'd182,8'd95} : s = 172;
	{8'd182,8'd96} : s = 170;
	{8'd182,8'd97} : s = 313;
	{8'd182,8'd98} : s = 52;
	{8'd182,8'd99} : s = 169;
	{8'd182,8'd100} : s = 166;
	{8'd182,8'd101} : s = 310;
	{8'd182,8'd102} : s = 165;
	{8'd182,8'd103} : s = 309;
	{8'd182,8'd104} : s = 307;
	{8'd182,8'd105} : s = 427;
	{8'd182,8'd106} : s = 6;
	{8'd182,8'd107} : s = 50;
	{8'd182,8'd108} : s = 49;
	{8'd182,8'd109} : s = 163;
	{8'd182,8'd110} : s = 44;
	{8'd182,8'd111} : s = 156;
	{8'd182,8'd112} : s = 154;
	{8'd182,8'd113} : s = 302;
	{8'd182,8'd114} : s = 42;
	{8'd182,8'd115} : s = 153;
	{8'd182,8'd116} : s = 150;
	{8'd182,8'd117} : s = 301;
	{8'd182,8'd118} : s = 149;
	{8'd182,8'd119} : s = 299;
	{8'd182,8'd120} : s = 295;
	{8'd182,8'd121} : s = 423;
	{8'd182,8'd122} : s = 41;
	{8'd182,8'd123} : s = 147;
	{8'd182,8'd124} : s = 142;
	{8'd182,8'd125} : s = 286;
	{8'd182,8'd126} : s = 141;
	{8'd182,8'd127} : s = 285;
	{8'd182,8'd128} : s = 283;
	{8'd182,8'd129} : s = 414;
	{8'd182,8'd130} : s = 139;
	{8'd182,8'd131} : s = 279;
	{8'd182,8'd132} : s = 271;
	{8'd182,8'd133} : s = 413;
	{8'd182,8'd134} : s = 248;
	{8'd182,8'd135} : s = 411;
	{8'd182,8'd136} : s = 407;
	{8'd182,8'd137} : s = 491;
	{8'd182,8'd138} : s = 5;
	{8'd182,8'd139} : s = 38;
	{8'd182,8'd140} : s = 37;
	{8'd182,8'd141} : s = 135;
	{8'd182,8'd142} : s = 35;
	{8'd182,8'd143} : s = 120;
	{8'd182,8'd144} : s = 116;
	{8'd182,8'd145} : s = 244;
	{8'd182,8'd146} : s = 28;
	{8'd182,8'd147} : s = 114;
	{8'd182,8'd148} : s = 113;
	{8'd182,8'd149} : s = 242;
	{8'd182,8'd150} : s = 108;
	{8'd182,8'd151} : s = 241;
	{8'd182,8'd152} : s = 236;
	{8'd182,8'd153} : s = 399;
	{8'd182,8'd154} : s = 26;
	{8'd182,8'd155} : s = 106;
	{8'd182,8'd156} : s = 105;
	{8'd182,8'd157} : s = 234;
	{8'd182,8'd158} : s = 102;
	{8'd182,8'd159} : s = 233;
	{8'd182,8'd160} : s = 230;
	{8'd182,8'd161} : s = 380;
	{8'd182,8'd162} : s = 101;
	{8'd182,8'd163} : s = 229;
	{8'd182,8'd164} : s = 227;
	{8'd182,8'd165} : s = 378;
	{8'd182,8'd166} : s = 220;
	{8'd182,8'd167} : s = 377;
	{8'd182,8'd168} : s = 374;
	{8'd182,8'd169} : s = 487;
	{8'd182,8'd170} : s = 25;
	{8'd182,8'd171} : s = 99;
	{8'd182,8'd172} : s = 92;
	{8'd182,8'd173} : s = 218;
	{8'd182,8'd174} : s = 90;
	{8'd182,8'd175} : s = 217;
	{8'd182,8'd176} : s = 214;
	{8'd182,8'd177} : s = 373;
	{8'd182,8'd178} : s = 89;
	{8'd182,8'd179} : s = 213;
	{8'd182,8'd180} : s = 211;
	{8'd182,8'd181} : s = 371;
	{8'd182,8'd182} : s = 206;
	{8'd182,8'd183} : s = 366;
	{8'd182,8'd184} : s = 365;
	{8'd182,8'd185} : s = 478;
	{8'd182,8'd186} : s = 86;
	{8'd182,8'd187} : s = 205;
	{8'd182,8'd188} : s = 203;
	{8'd182,8'd189} : s = 363;
	{8'd182,8'd190} : s = 199;
	{8'd182,8'd191} : s = 359;
	{8'd182,8'd192} : s = 350;
	{8'd182,8'd193} : s = 477;
	{8'd182,8'd194} : s = 188;
	{8'd182,8'd195} : s = 349;
	{8'd182,8'd196} : s = 347;
	{8'd182,8'd197} : s = 475;
	{8'd182,8'd198} : s = 343;
	{8'd182,8'd199} : s = 471;
	{8'd182,8'd200} : s = 463;
	{8'd182,8'd201} : s = 509;
	{8'd182,8'd202} : s = 3;
	{8'd182,8'd203} : s = 22;
	{8'd182,8'd204} : s = 21;
	{8'd182,8'd205} : s = 85;
	{8'd182,8'd206} : s = 19;
	{8'd182,8'd207} : s = 83;
	{8'd182,8'd208} : s = 78;
	{8'd182,8'd209} : s = 186;
	{8'd182,8'd210} : s = 14;
	{8'd182,8'd211} : s = 77;
	{8'd182,8'd212} : s = 75;
	{8'd182,8'd213} : s = 185;
	{8'd182,8'd214} : s = 71;
	{8'd182,8'd215} : s = 182;
	{8'd182,8'd216} : s = 181;
	{8'd182,8'd217} : s = 335;
	{8'd182,8'd218} : s = 13;
	{8'd182,8'd219} : s = 60;
	{8'd182,8'd220} : s = 58;
	{8'd182,8'd221} : s = 179;
	{8'd182,8'd222} : s = 57;
	{8'd182,8'd223} : s = 174;
	{8'd182,8'd224} : s = 173;
	{8'd182,8'd225} : s = 318;
	{8'd182,8'd226} : s = 54;
	{8'd182,8'd227} : s = 171;
	{8'd182,8'd228} : s = 167;
	{8'd182,8'd229} : s = 317;
	{8'd182,8'd230} : s = 158;
	{8'd182,8'd231} : s = 315;
	{8'd182,8'd232} : s = 311;
	{8'd182,8'd233} : s = 446;
	{8'd182,8'd234} : s = 11;
	{8'd182,8'd235} : s = 53;
	{8'd182,8'd236} : s = 51;
	{8'd182,8'd237} : s = 157;
	{8'd182,8'd238} : s = 46;
	{8'd182,8'd239} : s = 155;
	{8'd182,8'd240} : s = 151;
	{8'd182,8'd241} : s = 303;
	{8'd182,8'd242} : s = 45;
	{8'd182,8'd243} : s = 143;
	{8'd182,8'd244} : s = 124;
	{8'd182,8'd245} : s = 287;
	{8'd182,8'd246} : s = 122;
	{8'd182,8'd247} : s = 252;
	{8'd182,8'd248} : s = 250;
	{8'd182,8'd249} : s = 445;
	{8'd182,8'd250} : s = 43;
	{8'd182,8'd251} : s = 121;
	{8'd182,8'd252} : s = 118;
	{8'd182,8'd253} : s = 249;
	{8'd182,8'd254} : s = 117;
	{8'd182,8'd255} : s = 246;
	{8'd183,8'd0} : s = 483;
	{8'd183,8'd1} : s = 267;
	{8'd183,8'd2} : s = 395;
	{8'd183,8'd3} : s = 391;
	{8'd183,8'd4} : s = 476;
	{8'd183,8'd5} : s = 376;
	{8'd183,8'd6} : s = 474;
	{8'd183,8'd7} : s = 473;
	{8'd183,8'd8} : s = 506;
	{8'd183,8'd9} : s = 20;
	{8'd183,8'd10} : s = 104;
	{8'd183,8'd11} : s = 100;
	{8'd183,8'd12} : s = 263;
	{8'd183,8'd13} : s = 98;
	{8'd183,8'd14} : s = 240;
	{8'd183,8'd15} : s = 232;
	{8'd183,8'd16} : s = 372;
	{8'd183,8'd17} : s = 97;
	{8'd183,8'd18} : s = 228;
	{8'd183,8'd19} : s = 226;
	{8'd183,8'd20} : s = 370;
	{8'd183,8'd21} : s = 225;
	{8'd183,8'd22} : s = 369;
	{8'd183,8'd23} : s = 364;
	{8'd183,8'd24} : s = 470;
	{8'd183,8'd25} : s = 88;
	{8'd183,8'd26} : s = 216;
	{8'd183,8'd27} : s = 212;
	{8'd183,8'd28} : s = 362;
	{8'd183,8'd29} : s = 210;
	{8'd183,8'd30} : s = 361;
	{8'd183,8'd31} : s = 358;
	{8'd183,8'd32} : s = 469;
	{8'd183,8'd33} : s = 209;
	{8'd183,8'd34} : s = 357;
	{8'd183,8'd35} : s = 355;
	{8'd183,8'd36} : s = 467;
	{8'd183,8'd37} : s = 348;
	{8'd183,8'd38} : s = 462;
	{8'd183,8'd39} : s = 461;
	{8'd183,8'd40} : s = 505;
	{8'd183,8'd41} : s = 84;
	{8'd183,8'd42} : s = 204;
	{8'd183,8'd43} : s = 202;
	{8'd183,8'd44} : s = 346;
	{8'd183,8'd45} : s = 201;
	{8'd183,8'd46} : s = 345;
	{8'd183,8'd47} : s = 342;
	{8'd183,8'd48} : s = 459;
	{8'd183,8'd49} : s = 198;
	{8'd183,8'd50} : s = 341;
	{8'd183,8'd51} : s = 339;
	{8'd183,8'd52} : s = 455;
	{8'd183,8'd53} : s = 334;
	{8'd183,8'd54} : s = 444;
	{8'd183,8'd55} : s = 442;
	{8'd183,8'd56} : s = 502;
	{8'd183,8'd57} : s = 197;
	{8'd183,8'd58} : s = 333;
	{8'd183,8'd59} : s = 331;
	{8'd183,8'd60} : s = 441;
	{8'd183,8'd61} : s = 327;
	{8'd183,8'd62} : s = 438;
	{8'd183,8'd63} : s = 437;
	{8'd183,8'd64} : s = 501;
	{8'd183,8'd65} : s = 316;
	{8'd183,8'd66} : s = 435;
	{8'd183,8'd67} : s = 430;
	{8'd183,8'd68} : s = 499;
	{8'd183,8'd69} : s = 429;
	{8'd183,8'd70} : s = 494;
	{8'd183,8'd71} : s = 493;
	{8'd183,8'd72} : s = 510;
	{8'd183,8'd73} : s = 1;
	{8'd183,8'd74} : s = 18;
	{8'd183,8'd75} : s = 17;
	{8'd183,8'd76} : s = 82;
	{8'd183,8'd77} : s = 12;
	{8'd183,8'd78} : s = 81;
	{8'd183,8'd79} : s = 76;
	{8'd183,8'd80} : s = 195;
	{8'd183,8'd81} : s = 10;
	{8'd183,8'd82} : s = 74;
	{8'd183,8'd83} : s = 73;
	{8'd183,8'd84} : s = 184;
	{8'd183,8'd85} : s = 70;
	{8'd183,8'd86} : s = 180;
	{8'd183,8'd87} : s = 178;
	{8'd183,8'd88} : s = 314;
	{8'd183,8'd89} : s = 9;
	{8'd183,8'd90} : s = 69;
	{8'd183,8'd91} : s = 67;
	{8'd183,8'd92} : s = 177;
	{8'd183,8'd93} : s = 56;
	{8'd183,8'd94} : s = 172;
	{8'd183,8'd95} : s = 170;
	{8'd183,8'd96} : s = 313;
	{8'd183,8'd97} : s = 52;
	{8'd183,8'd98} : s = 169;
	{8'd183,8'd99} : s = 166;
	{8'd183,8'd100} : s = 310;
	{8'd183,8'd101} : s = 165;
	{8'd183,8'd102} : s = 309;
	{8'd183,8'd103} : s = 307;
	{8'd183,8'd104} : s = 427;
	{8'd183,8'd105} : s = 6;
	{8'd183,8'd106} : s = 50;
	{8'd183,8'd107} : s = 49;
	{8'd183,8'd108} : s = 163;
	{8'd183,8'd109} : s = 44;
	{8'd183,8'd110} : s = 156;
	{8'd183,8'd111} : s = 154;
	{8'd183,8'd112} : s = 302;
	{8'd183,8'd113} : s = 42;
	{8'd183,8'd114} : s = 153;
	{8'd183,8'd115} : s = 150;
	{8'd183,8'd116} : s = 301;
	{8'd183,8'd117} : s = 149;
	{8'd183,8'd118} : s = 299;
	{8'd183,8'd119} : s = 295;
	{8'd183,8'd120} : s = 423;
	{8'd183,8'd121} : s = 41;
	{8'd183,8'd122} : s = 147;
	{8'd183,8'd123} : s = 142;
	{8'd183,8'd124} : s = 286;
	{8'd183,8'd125} : s = 141;
	{8'd183,8'd126} : s = 285;
	{8'd183,8'd127} : s = 283;
	{8'd183,8'd128} : s = 414;
	{8'd183,8'd129} : s = 139;
	{8'd183,8'd130} : s = 279;
	{8'd183,8'd131} : s = 271;
	{8'd183,8'd132} : s = 413;
	{8'd183,8'd133} : s = 248;
	{8'd183,8'd134} : s = 411;
	{8'd183,8'd135} : s = 407;
	{8'd183,8'd136} : s = 491;
	{8'd183,8'd137} : s = 5;
	{8'd183,8'd138} : s = 38;
	{8'd183,8'd139} : s = 37;
	{8'd183,8'd140} : s = 135;
	{8'd183,8'd141} : s = 35;
	{8'd183,8'd142} : s = 120;
	{8'd183,8'd143} : s = 116;
	{8'd183,8'd144} : s = 244;
	{8'd183,8'd145} : s = 28;
	{8'd183,8'd146} : s = 114;
	{8'd183,8'd147} : s = 113;
	{8'd183,8'd148} : s = 242;
	{8'd183,8'd149} : s = 108;
	{8'd183,8'd150} : s = 241;
	{8'd183,8'd151} : s = 236;
	{8'd183,8'd152} : s = 399;
	{8'd183,8'd153} : s = 26;
	{8'd183,8'd154} : s = 106;
	{8'd183,8'd155} : s = 105;
	{8'd183,8'd156} : s = 234;
	{8'd183,8'd157} : s = 102;
	{8'd183,8'd158} : s = 233;
	{8'd183,8'd159} : s = 230;
	{8'd183,8'd160} : s = 380;
	{8'd183,8'd161} : s = 101;
	{8'd183,8'd162} : s = 229;
	{8'd183,8'd163} : s = 227;
	{8'd183,8'd164} : s = 378;
	{8'd183,8'd165} : s = 220;
	{8'd183,8'd166} : s = 377;
	{8'd183,8'd167} : s = 374;
	{8'd183,8'd168} : s = 487;
	{8'd183,8'd169} : s = 25;
	{8'd183,8'd170} : s = 99;
	{8'd183,8'd171} : s = 92;
	{8'd183,8'd172} : s = 218;
	{8'd183,8'd173} : s = 90;
	{8'd183,8'd174} : s = 217;
	{8'd183,8'd175} : s = 214;
	{8'd183,8'd176} : s = 373;
	{8'd183,8'd177} : s = 89;
	{8'd183,8'd178} : s = 213;
	{8'd183,8'd179} : s = 211;
	{8'd183,8'd180} : s = 371;
	{8'd183,8'd181} : s = 206;
	{8'd183,8'd182} : s = 366;
	{8'd183,8'd183} : s = 365;
	{8'd183,8'd184} : s = 478;
	{8'd183,8'd185} : s = 86;
	{8'd183,8'd186} : s = 205;
	{8'd183,8'd187} : s = 203;
	{8'd183,8'd188} : s = 363;
	{8'd183,8'd189} : s = 199;
	{8'd183,8'd190} : s = 359;
	{8'd183,8'd191} : s = 350;
	{8'd183,8'd192} : s = 477;
	{8'd183,8'd193} : s = 188;
	{8'd183,8'd194} : s = 349;
	{8'd183,8'd195} : s = 347;
	{8'd183,8'd196} : s = 475;
	{8'd183,8'd197} : s = 343;
	{8'd183,8'd198} : s = 471;
	{8'd183,8'd199} : s = 463;
	{8'd183,8'd200} : s = 509;
	{8'd183,8'd201} : s = 3;
	{8'd183,8'd202} : s = 22;
	{8'd183,8'd203} : s = 21;
	{8'd183,8'd204} : s = 85;
	{8'd183,8'd205} : s = 19;
	{8'd183,8'd206} : s = 83;
	{8'd183,8'd207} : s = 78;
	{8'd183,8'd208} : s = 186;
	{8'd183,8'd209} : s = 14;
	{8'd183,8'd210} : s = 77;
	{8'd183,8'd211} : s = 75;
	{8'd183,8'd212} : s = 185;
	{8'd183,8'd213} : s = 71;
	{8'd183,8'd214} : s = 182;
	{8'd183,8'd215} : s = 181;
	{8'd183,8'd216} : s = 335;
	{8'd183,8'd217} : s = 13;
	{8'd183,8'd218} : s = 60;
	{8'd183,8'd219} : s = 58;
	{8'd183,8'd220} : s = 179;
	{8'd183,8'd221} : s = 57;
	{8'd183,8'd222} : s = 174;
	{8'd183,8'd223} : s = 173;
	{8'd183,8'd224} : s = 318;
	{8'd183,8'd225} : s = 54;
	{8'd183,8'd226} : s = 171;
	{8'd183,8'd227} : s = 167;
	{8'd183,8'd228} : s = 317;
	{8'd183,8'd229} : s = 158;
	{8'd183,8'd230} : s = 315;
	{8'd183,8'd231} : s = 311;
	{8'd183,8'd232} : s = 446;
	{8'd183,8'd233} : s = 11;
	{8'd183,8'd234} : s = 53;
	{8'd183,8'd235} : s = 51;
	{8'd183,8'd236} : s = 157;
	{8'd183,8'd237} : s = 46;
	{8'd183,8'd238} : s = 155;
	{8'd183,8'd239} : s = 151;
	{8'd183,8'd240} : s = 303;
	{8'd183,8'd241} : s = 45;
	{8'd183,8'd242} : s = 143;
	{8'd183,8'd243} : s = 124;
	{8'd183,8'd244} : s = 287;
	{8'd183,8'd245} : s = 122;
	{8'd183,8'd246} : s = 252;
	{8'd183,8'd247} : s = 250;
	{8'd183,8'd248} : s = 445;
	{8'd183,8'd249} : s = 43;
	{8'd183,8'd250} : s = 121;
	{8'd183,8'd251} : s = 118;
	{8'd183,8'd252} : s = 249;
	{8'd183,8'd253} : s = 117;
	{8'd183,8'd254} : s = 246;
	{8'd183,8'd255} : s = 245;
	{8'd184,8'd0} : s = 267;
	{8'd184,8'd1} : s = 395;
	{8'd184,8'd2} : s = 391;
	{8'd184,8'd3} : s = 476;
	{8'd184,8'd4} : s = 376;
	{8'd184,8'd5} : s = 474;
	{8'd184,8'd6} : s = 473;
	{8'd184,8'd7} : s = 506;
	{8'd184,8'd8} : s = 20;
	{8'd184,8'd9} : s = 104;
	{8'd184,8'd10} : s = 100;
	{8'd184,8'd11} : s = 263;
	{8'd184,8'd12} : s = 98;
	{8'd184,8'd13} : s = 240;
	{8'd184,8'd14} : s = 232;
	{8'd184,8'd15} : s = 372;
	{8'd184,8'd16} : s = 97;
	{8'd184,8'd17} : s = 228;
	{8'd184,8'd18} : s = 226;
	{8'd184,8'd19} : s = 370;
	{8'd184,8'd20} : s = 225;
	{8'd184,8'd21} : s = 369;
	{8'd184,8'd22} : s = 364;
	{8'd184,8'd23} : s = 470;
	{8'd184,8'd24} : s = 88;
	{8'd184,8'd25} : s = 216;
	{8'd184,8'd26} : s = 212;
	{8'd184,8'd27} : s = 362;
	{8'd184,8'd28} : s = 210;
	{8'd184,8'd29} : s = 361;
	{8'd184,8'd30} : s = 358;
	{8'd184,8'd31} : s = 469;
	{8'd184,8'd32} : s = 209;
	{8'd184,8'd33} : s = 357;
	{8'd184,8'd34} : s = 355;
	{8'd184,8'd35} : s = 467;
	{8'd184,8'd36} : s = 348;
	{8'd184,8'd37} : s = 462;
	{8'd184,8'd38} : s = 461;
	{8'd184,8'd39} : s = 505;
	{8'd184,8'd40} : s = 84;
	{8'd184,8'd41} : s = 204;
	{8'd184,8'd42} : s = 202;
	{8'd184,8'd43} : s = 346;
	{8'd184,8'd44} : s = 201;
	{8'd184,8'd45} : s = 345;
	{8'd184,8'd46} : s = 342;
	{8'd184,8'd47} : s = 459;
	{8'd184,8'd48} : s = 198;
	{8'd184,8'd49} : s = 341;
	{8'd184,8'd50} : s = 339;
	{8'd184,8'd51} : s = 455;
	{8'd184,8'd52} : s = 334;
	{8'd184,8'd53} : s = 444;
	{8'd184,8'd54} : s = 442;
	{8'd184,8'd55} : s = 502;
	{8'd184,8'd56} : s = 197;
	{8'd184,8'd57} : s = 333;
	{8'd184,8'd58} : s = 331;
	{8'd184,8'd59} : s = 441;
	{8'd184,8'd60} : s = 327;
	{8'd184,8'd61} : s = 438;
	{8'd184,8'd62} : s = 437;
	{8'd184,8'd63} : s = 501;
	{8'd184,8'd64} : s = 316;
	{8'd184,8'd65} : s = 435;
	{8'd184,8'd66} : s = 430;
	{8'd184,8'd67} : s = 499;
	{8'd184,8'd68} : s = 429;
	{8'd184,8'd69} : s = 494;
	{8'd184,8'd70} : s = 493;
	{8'd184,8'd71} : s = 510;
	{8'd184,8'd72} : s = 1;
	{8'd184,8'd73} : s = 18;
	{8'd184,8'd74} : s = 17;
	{8'd184,8'd75} : s = 82;
	{8'd184,8'd76} : s = 12;
	{8'd184,8'd77} : s = 81;
	{8'd184,8'd78} : s = 76;
	{8'd184,8'd79} : s = 195;
	{8'd184,8'd80} : s = 10;
	{8'd184,8'd81} : s = 74;
	{8'd184,8'd82} : s = 73;
	{8'd184,8'd83} : s = 184;
	{8'd184,8'd84} : s = 70;
	{8'd184,8'd85} : s = 180;
	{8'd184,8'd86} : s = 178;
	{8'd184,8'd87} : s = 314;
	{8'd184,8'd88} : s = 9;
	{8'd184,8'd89} : s = 69;
	{8'd184,8'd90} : s = 67;
	{8'd184,8'd91} : s = 177;
	{8'd184,8'd92} : s = 56;
	{8'd184,8'd93} : s = 172;
	{8'd184,8'd94} : s = 170;
	{8'd184,8'd95} : s = 313;
	{8'd184,8'd96} : s = 52;
	{8'd184,8'd97} : s = 169;
	{8'd184,8'd98} : s = 166;
	{8'd184,8'd99} : s = 310;
	{8'd184,8'd100} : s = 165;
	{8'd184,8'd101} : s = 309;
	{8'd184,8'd102} : s = 307;
	{8'd184,8'd103} : s = 427;
	{8'd184,8'd104} : s = 6;
	{8'd184,8'd105} : s = 50;
	{8'd184,8'd106} : s = 49;
	{8'd184,8'd107} : s = 163;
	{8'd184,8'd108} : s = 44;
	{8'd184,8'd109} : s = 156;
	{8'd184,8'd110} : s = 154;
	{8'd184,8'd111} : s = 302;
	{8'd184,8'd112} : s = 42;
	{8'd184,8'd113} : s = 153;
	{8'd184,8'd114} : s = 150;
	{8'd184,8'd115} : s = 301;
	{8'd184,8'd116} : s = 149;
	{8'd184,8'd117} : s = 299;
	{8'd184,8'd118} : s = 295;
	{8'd184,8'd119} : s = 423;
	{8'd184,8'd120} : s = 41;
	{8'd184,8'd121} : s = 147;
	{8'd184,8'd122} : s = 142;
	{8'd184,8'd123} : s = 286;
	{8'd184,8'd124} : s = 141;
	{8'd184,8'd125} : s = 285;
	{8'd184,8'd126} : s = 283;
	{8'd184,8'd127} : s = 414;
	{8'd184,8'd128} : s = 139;
	{8'd184,8'd129} : s = 279;
	{8'd184,8'd130} : s = 271;
	{8'd184,8'd131} : s = 413;
	{8'd184,8'd132} : s = 248;
	{8'd184,8'd133} : s = 411;
	{8'd184,8'd134} : s = 407;
	{8'd184,8'd135} : s = 491;
	{8'd184,8'd136} : s = 5;
	{8'd184,8'd137} : s = 38;
	{8'd184,8'd138} : s = 37;
	{8'd184,8'd139} : s = 135;
	{8'd184,8'd140} : s = 35;
	{8'd184,8'd141} : s = 120;
	{8'd184,8'd142} : s = 116;
	{8'd184,8'd143} : s = 244;
	{8'd184,8'd144} : s = 28;
	{8'd184,8'd145} : s = 114;
	{8'd184,8'd146} : s = 113;
	{8'd184,8'd147} : s = 242;
	{8'd184,8'd148} : s = 108;
	{8'd184,8'd149} : s = 241;
	{8'd184,8'd150} : s = 236;
	{8'd184,8'd151} : s = 399;
	{8'd184,8'd152} : s = 26;
	{8'd184,8'd153} : s = 106;
	{8'd184,8'd154} : s = 105;
	{8'd184,8'd155} : s = 234;
	{8'd184,8'd156} : s = 102;
	{8'd184,8'd157} : s = 233;
	{8'd184,8'd158} : s = 230;
	{8'd184,8'd159} : s = 380;
	{8'd184,8'd160} : s = 101;
	{8'd184,8'd161} : s = 229;
	{8'd184,8'd162} : s = 227;
	{8'd184,8'd163} : s = 378;
	{8'd184,8'd164} : s = 220;
	{8'd184,8'd165} : s = 377;
	{8'd184,8'd166} : s = 374;
	{8'd184,8'd167} : s = 487;
	{8'd184,8'd168} : s = 25;
	{8'd184,8'd169} : s = 99;
	{8'd184,8'd170} : s = 92;
	{8'd184,8'd171} : s = 218;
	{8'd184,8'd172} : s = 90;
	{8'd184,8'd173} : s = 217;
	{8'd184,8'd174} : s = 214;
	{8'd184,8'd175} : s = 373;
	{8'd184,8'd176} : s = 89;
	{8'd184,8'd177} : s = 213;
	{8'd184,8'd178} : s = 211;
	{8'd184,8'd179} : s = 371;
	{8'd184,8'd180} : s = 206;
	{8'd184,8'd181} : s = 366;
	{8'd184,8'd182} : s = 365;
	{8'd184,8'd183} : s = 478;
	{8'd184,8'd184} : s = 86;
	{8'd184,8'd185} : s = 205;
	{8'd184,8'd186} : s = 203;
	{8'd184,8'd187} : s = 363;
	{8'd184,8'd188} : s = 199;
	{8'd184,8'd189} : s = 359;
	{8'd184,8'd190} : s = 350;
	{8'd184,8'd191} : s = 477;
	{8'd184,8'd192} : s = 188;
	{8'd184,8'd193} : s = 349;
	{8'd184,8'd194} : s = 347;
	{8'd184,8'd195} : s = 475;
	{8'd184,8'd196} : s = 343;
	{8'd184,8'd197} : s = 471;
	{8'd184,8'd198} : s = 463;
	{8'd184,8'd199} : s = 509;
	{8'd184,8'd200} : s = 3;
	{8'd184,8'd201} : s = 22;
	{8'd184,8'd202} : s = 21;
	{8'd184,8'd203} : s = 85;
	{8'd184,8'd204} : s = 19;
	{8'd184,8'd205} : s = 83;
	{8'd184,8'd206} : s = 78;
	{8'd184,8'd207} : s = 186;
	{8'd184,8'd208} : s = 14;
	{8'd184,8'd209} : s = 77;
	{8'd184,8'd210} : s = 75;
	{8'd184,8'd211} : s = 185;
	{8'd184,8'd212} : s = 71;
	{8'd184,8'd213} : s = 182;
	{8'd184,8'd214} : s = 181;
	{8'd184,8'd215} : s = 335;
	{8'd184,8'd216} : s = 13;
	{8'd184,8'd217} : s = 60;
	{8'd184,8'd218} : s = 58;
	{8'd184,8'd219} : s = 179;
	{8'd184,8'd220} : s = 57;
	{8'd184,8'd221} : s = 174;
	{8'd184,8'd222} : s = 173;
	{8'd184,8'd223} : s = 318;
	{8'd184,8'd224} : s = 54;
	{8'd184,8'd225} : s = 171;
	{8'd184,8'd226} : s = 167;
	{8'd184,8'd227} : s = 317;
	{8'd184,8'd228} : s = 158;
	{8'd184,8'd229} : s = 315;
	{8'd184,8'd230} : s = 311;
	{8'd184,8'd231} : s = 446;
	{8'd184,8'd232} : s = 11;
	{8'd184,8'd233} : s = 53;
	{8'd184,8'd234} : s = 51;
	{8'd184,8'd235} : s = 157;
	{8'd184,8'd236} : s = 46;
	{8'd184,8'd237} : s = 155;
	{8'd184,8'd238} : s = 151;
	{8'd184,8'd239} : s = 303;
	{8'd184,8'd240} : s = 45;
	{8'd184,8'd241} : s = 143;
	{8'd184,8'd242} : s = 124;
	{8'd184,8'd243} : s = 287;
	{8'd184,8'd244} : s = 122;
	{8'd184,8'd245} : s = 252;
	{8'd184,8'd246} : s = 250;
	{8'd184,8'd247} : s = 445;
	{8'd184,8'd248} : s = 43;
	{8'd184,8'd249} : s = 121;
	{8'd184,8'd250} : s = 118;
	{8'd184,8'd251} : s = 249;
	{8'd184,8'd252} : s = 117;
	{8'd184,8'd253} : s = 246;
	{8'd184,8'd254} : s = 245;
	{8'd184,8'd255} : s = 443;
	{8'd185,8'd0} : s = 395;
	{8'd185,8'd1} : s = 391;
	{8'd185,8'd2} : s = 476;
	{8'd185,8'd3} : s = 376;
	{8'd185,8'd4} : s = 474;
	{8'd185,8'd5} : s = 473;
	{8'd185,8'd6} : s = 506;
	{8'd185,8'd7} : s = 20;
	{8'd185,8'd8} : s = 104;
	{8'd185,8'd9} : s = 100;
	{8'd185,8'd10} : s = 263;
	{8'd185,8'd11} : s = 98;
	{8'd185,8'd12} : s = 240;
	{8'd185,8'd13} : s = 232;
	{8'd185,8'd14} : s = 372;
	{8'd185,8'd15} : s = 97;
	{8'd185,8'd16} : s = 228;
	{8'd185,8'd17} : s = 226;
	{8'd185,8'd18} : s = 370;
	{8'd185,8'd19} : s = 225;
	{8'd185,8'd20} : s = 369;
	{8'd185,8'd21} : s = 364;
	{8'd185,8'd22} : s = 470;
	{8'd185,8'd23} : s = 88;
	{8'd185,8'd24} : s = 216;
	{8'd185,8'd25} : s = 212;
	{8'd185,8'd26} : s = 362;
	{8'd185,8'd27} : s = 210;
	{8'd185,8'd28} : s = 361;
	{8'd185,8'd29} : s = 358;
	{8'd185,8'd30} : s = 469;
	{8'd185,8'd31} : s = 209;
	{8'd185,8'd32} : s = 357;
	{8'd185,8'd33} : s = 355;
	{8'd185,8'd34} : s = 467;
	{8'd185,8'd35} : s = 348;
	{8'd185,8'd36} : s = 462;
	{8'd185,8'd37} : s = 461;
	{8'd185,8'd38} : s = 505;
	{8'd185,8'd39} : s = 84;
	{8'd185,8'd40} : s = 204;
	{8'd185,8'd41} : s = 202;
	{8'd185,8'd42} : s = 346;
	{8'd185,8'd43} : s = 201;
	{8'd185,8'd44} : s = 345;
	{8'd185,8'd45} : s = 342;
	{8'd185,8'd46} : s = 459;
	{8'd185,8'd47} : s = 198;
	{8'd185,8'd48} : s = 341;
	{8'd185,8'd49} : s = 339;
	{8'd185,8'd50} : s = 455;
	{8'd185,8'd51} : s = 334;
	{8'd185,8'd52} : s = 444;
	{8'd185,8'd53} : s = 442;
	{8'd185,8'd54} : s = 502;
	{8'd185,8'd55} : s = 197;
	{8'd185,8'd56} : s = 333;
	{8'd185,8'd57} : s = 331;
	{8'd185,8'd58} : s = 441;
	{8'd185,8'd59} : s = 327;
	{8'd185,8'd60} : s = 438;
	{8'd185,8'd61} : s = 437;
	{8'd185,8'd62} : s = 501;
	{8'd185,8'd63} : s = 316;
	{8'd185,8'd64} : s = 435;
	{8'd185,8'd65} : s = 430;
	{8'd185,8'd66} : s = 499;
	{8'd185,8'd67} : s = 429;
	{8'd185,8'd68} : s = 494;
	{8'd185,8'd69} : s = 493;
	{8'd185,8'd70} : s = 510;
	{8'd185,8'd71} : s = 1;
	{8'd185,8'd72} : s = 18;
	{8'd185,8'd73} : s = 17;
	{8'd185,8'd74} : s = 82;
	{8'd185,8'd75} : s = 12;
	{8'd185,8'd76} : s = 81;
	{8'd185,8'd77} : s = 76;
	{8'd185,8'd78} : s = 195;
	{8'd185,8'd79} : s = 10;
	{8'd185,8'd80} : s = 74;
	{8'd185,8'd81} : s = 73;
	{8'd185,8'd82} : s = 184;
	{8'd185,8'd83} : s = 70;
	{8'd185,8'd84} : s = 180;
	{8'd185,8'd85} : s = 178;
	{8'd185,8'd86} : s = 314;
	{8'd185,8'd87} : s = 9;
	{8'd185,8'd88} : s = 69;
	{8'd185,8'd89} : s = 67;
	{8'd185,8'd90} : s = 177;
	{8'd185,8'd91} : s = 56;
	{8'd185,8'd92} : s = 172;
	{8'd185,8'd93} : s = 170;
	{8'd185,8'd94} : s = 313;
	{8'd185,8'd95} : s = 52;
	{8'd185,8'd96} : s = 169;
	{8'd185,8'd97} : s = 166;
	{8'd185,8'd98} : s = 310;
	{8'd185,8'd99} : s = 165;
	{8'd185,8'd100} : s = 309;
	{8'd185,8'd101} : s = 307;
	{8'd185,8'd102} : s = 427;
	{8'd185,8'd103} : s = 6;
	{8'd185,8'd104} : s = 50;
	{8'd185,8'd105} : s = 49;
	{8'd185,8'd106} : s = 163;
	{8'd185,8'd107} : s = 44;
	{8'd185,8'd108} : s = 156;
	{8'd185,8'd109} : s = 154;
	{8'd185,8'd110} : s = 302;
	{8'd185,8'd111} : s = 42;
	{8'd185,8'd112} : s = 153;
	{8'd185,8'd113} : s = 150;
	{8'd185,8'd114} : s = 301;
	{8'd185,8'd115} : s = 149;
	{8'd185,8'd116} : s = 299;
	{8'd185,8'd117} : s = 295;
	{8'd185,8'd118} : s = 423;
	{8'd185,8'd119} : s = 41;
	{8'd185,8'd120} : s = 147;
	{8'd185,8'd121} : s = 142;
	{8'd185,8'd122} : s = 286;
	{8'd185,8'd123} : s = 141;
	{8'd185,8'd124} : s = 285;
	{8'd185,8'd125} : s = 283;
	{8'd185,8'd126} : s = 414;
	{8'd185,8'd127} : s = 139;
	{8'd185,8'd128} : s = 279;
	{8'd185,8'd129} : s = 271;
	{8'd185,8'd130} : s = 413;
	{8'd185,8'd131} : s = 248;
	{8'd185,8'd132} : s = 411;
	{8'd185,8'd133} : s = 407;
	{8'd185,8'd134} : s = 491;
	{8'd185,8'd135} : s = 5;
	{8'd185,8'd136} : s = 38;
	{8'd185,8'd137} : s = 37;
	{8'd185,8'd138} : s = 135;
	{8'd185,8'd139} : s = 35;
	{8'd185,8'd140} : s = 120;
	{8'd185,8'd141} : s = 116;
	{8'd185,8'd142} : s = 244;
	{8'd185,8'd143} : s = 28;
	{8'd185,8'd144} : s = 114;
	{8'd185,8'd145} : s = 113;
	{8'd185,8'd146} : s = 242;
	{8'd185,8'd147} : s = 108;
	{8'd185,8'd148} : s = 241;
	{8'd185,8'd149} : s = 236;
	{8'd185,8'd150} : s = 399;
	{8'd185,8'd151} : s = 26;
	{8'd185,8'd152} : s = 106;
	{8'd185,8'd153} : s = 105;
	{8'd185,8'd154} : s = 234;
	{8'd185,8'd155} : s = 102;
	{8'd185,8'd156} : s = 233;
	{8'd185,8'd157} : s = 230;
	{8'd185,8'd158} : s = 380;
	{8'd185,8'd159} : s = 101;
	{8'd185,8'd160} : s = 229;
	{8'd185,8'd161} : s = 227;
	{8'd185,8'd162} : s = 378;
	{8'd185,8'd163} : s = 220;
	{8'd185,8'd164} : s = 377;
	{8'd185,8'd165} : s = 374;
	{8'd185,8'd166} : s = 487;
	{8'd185,8'd167} : s = 25;
	{8'd185,8'd168} : s = 99;
	{8'd185,8'd169} : s = 92;
	{8'd185,8'd170} : s = 218;
	{8'd185,8'd171} : s = 90;
	{8'd185,8'd172} : s = 217;
	{8'd185,8'd173} : s = 214;
	{8'd185,8'd174} : s = 373;
	{8'd185,8'd175} : s = 89;
	{8'd185,8'd176} : s = 213;
	{8'd185,8'd177} : s = 211;
	{8'd185,8'd178} : s = 371;
	{8'd185,8'd179} : s = 206;
	{8'd185,8'd180} : s = 366;
	{8'd185,8'd181} : s = 365;
	{8'd185,8'd182} : s = 478;
	{8'd185,8'd183} : s = 86;
	{8'd185,8'd184} : s = 205;
	{8'd185,8'd185} : s = 203;
	{8'd185,8'd186} : s = 363;
	{8'd185,8'd187} : s = 199;
	{8'd185,8'd188} : s = 359;
	{8'd185,8'd189} : s = 350;
	{8'd185,8'd190} : s = 477;
	{8'd185,8'd191} : s = 188;
	{8'd185,8'd192} : s = 349;
	{8'd185,8'd193} : s = 347;
	{8'd185,8'd194} : s = 475;
	{8'd185,8'd195} : s = 343;
	{8'd185,8'd196} : s = 471;
	{8'd185,8'd197} : s = 463;
	{8'd185,8'd198} : s = 509;
	{8'd185,8'd199} : s = 3;
	{8'd185,8'd200} : s = 22;
	{8'd185,8'd201} : s = 21;
	{8'd185,8'd202} : s = 85;
	{8'd185,8'd203} : s = 19;
	{8'd185,8'd204} : s = 83;
	{8'd185,8'd205} : s = 78;
	{8'd185,8'd206} : s = 186;
	{8'd185,8'd207} : s = 14;
	{8'd185,8'd208} : s = 77;
	{8'd185,8'd209} : s = 75;
	{8'd185,8'd210} : s = 185;
	{8'd185,8'd211} : s = 71;
	{8'd185,8'd212} : s = 182;
	{8'd185,8'd213} : s = 181;
	{8'd185,8'd214} : s = 335;
	{8'd185,8'd215} : s = 13;
	{8'd185,8'd216} : s = 60;
	{8'd185,8'd217} : s = 58;
	{8'd185,8'd218} : s = 179;
	{8'd185,8'd219} : s = 57;
	{8'd185,8'd220} : s = 174;
	{8'd185,8'd221} : s = 173;
	{8'd185,8'd222} : s = 318;
	{8'd185,8'd223} : s = 54;
	{8'd185,8'd224} : s = 171;
	{8'd185,8'd225} : s = 167;
	{8'd185,8'd226} : s = 317;
	{8'd185,8'd227} : s = 158;
	{8'd185,8'd228} : s = 315;
	{8'd185,8'd229} : s = 311;
	{8'd185,8'd230} : s = 446;
	{8'd185,8'd231} : s = 11;
	{8'd185,8'd232} : s = 53;
	{8'd185,8'd233} : s = 51;
	{8'd185,8'd234} : s = 157;
	{8'd185,8'd235} : s = 46;
	{8'd185,8'd236} : s = 155;
	{8'd185,8'd237} : s = 151;
	{8'd185,8'd238} : s = 303;
	{8'd185,8'd239} : s = 45;
	{8'd185,8'd240} : s = 143;
	{8'd185,8'd241} : s = 124;
	{8'd185,8'd242} : s = 287;
	{8'd185,8'd243} : s = 122;
	{8'd185,8'd244} : s = 252;
	{8'd185,8'd245} : s = 250;
	{8'd185,8'd246} : s = 445;
	{8'd185,8'd247} : s = 43;
	{8'd185,8'd248} : s = 121;
	{8'd185,8'd249} : s = 118;
	{8'd185,8'd250} : s = 249;
	{8'd185,8'd251} : s = 117;
	{8'd185,8'd252} : s = 246;
	{8'd185,8'd253} : s = 245;
	{8'd185,8'd254} : s = 443;
	{8'd185,8'd255} : s = 115;
	{8'd186,8'd0} : s = 391;
	{8'd186,8'd1} : s = 476;
	{8'd186,8'd2} : s = 376;
	{8'd186,8'd3} : s = 474;
	{8'd186,8'd4} : s = 473;
	{8'd186,8'd5} : s = 506;
	{8'd186,8'd6} : s = 20;
	{8'd186,8'd7} : s = 104;
	{8'd186,8'd8} : s = 100;
	{8'd186,8'd9} : s = 263;
	{8'd186,8'd10} : s = 98;
	{8'd186,8'd11} : s = 240;
	{8'd186,8'd12} : s = 232;
	{8'd186,8'd13} : s = 372;
	{8'd186,8'd14} : s = 97;
	{8'd186,8'd15} : s = 228;
	{8'd186,8'd16} : s = 226;
	{8'd186,8'd17} : s = 370;
	{8'd186,8'd18} : s = 225;
	{8'd186,8'd19} : s = 369;
	{8'd186,8'd20} : s = 364;
	{8'd186,8'd21} : s = 470;
	{8'd186,8'd22} : s = 88;
	{8'd186,8'd23} : s = 216;
	{8'd186,8'd24} : s = 212;
	{8'd186,8'd25} : s = 362;
	{8'd186,8'd26} : s = 210;
	{8'd186,8'd27} : s = 361;
	{8'd186,8'd28} : s = 358;
	{8'd186,8'd29} : s = 469;
	{8'd186,8'd30} : s = 209;
	{8'd186,8'd31} : s = 357;
	{8'd186,8'd32} : s = 355;
	{8'd186,8'd33} : s = 467;
	{8'd186,8'd34} : s = 348;
	{8'd186,8'd35} : s = 462;
	{8'd186,8'd36} : s = 461;
	{8'd186,8'd37} : s = 505;
	{8'd186,8'd38} : s = 84;
	{8'd186,8'd39} : s = 204;
	{8'd186,8'd40} : s = 202;
	{8'd186,8'd41} : s = 346;
	{8'd186,8'd42} : s = 201;
	{8'd186,8'd43} : s = 345;
	{8'd186,8'd44} : s = 342;
	{8'd186,8'd45} : s = 459;
	{8'd186,8'd46} : s = 198;
	{8'd186,8'd47} : s = 341;
	{8'd186,8'd48} : s = 339;
	{8'd186,8'd49} : s = 455;
	{8'd186,8'd50} : s = 334;
	{8'd186,8'd51} : s = 444;
	{8'd186,8'd52} : s = 442;
	{8'd186,8'd53} : s = 502;
	{8'd186,8'd54} : s = 197;
	{8'd186,8'd55} : s = 333;
	{8'd186,8'd56} : s = 331;
	{8'd186,8'd57} : s = 441;
	{8'd186,8'd58} : s = 327;
	{8'd186,8'd59} : s = 438;
	{8'd186,8'd60} : s = 437;
	{8'd186,8'd61} : s = 501;
	{8'd186,8'd62} : s = 316;
	{8'd186,8'd63} : s = 435;
	{8'd186,8'd64} : s = 430;
	{8'd186,8'd65} : s = 499;
	{8'd186,8'd66} : s = 429;
	{8'd186,8'd67} : s = 494;
	{8'd186,8'd68} : s = 493;
	{8'd186,8'd69} : s = 510;
	{8'd186,8'd70} : s = 1;
	{8'd186,8'd71} : s = 18;
	{8'd186,8'd72} : s = 17;
	{8'd186,8'd73} : s = 82;
	{8'd186,8'd74} : s = 12;
	{8'd186,8'd75} : s = 81;
	{8'd186,8'd76} : s = 76;
	{8'd186,8'd77} : s = 195;
	{8'd186,8'd78} : s = 10;
	{8'd186,8'd79} : s = 74;
	{8'd186,8'd80} : s = 73;
	{8'd186,8'd81} : s = 184;
	{8'd186,8'd82} : s = 70;
	{8'd186,8'd83} : s = 180;
	{8'd186,8'd84} : s = 178;
	{8'd186,8'd85} : s = 314;
	{8'd186,8'd86} : s = 9;
	{8'd186,8'd87} : s = 69;
	{8'd186,8'd88} : s = 67;
	{8'd186,8'd89} : s = 177;
	{8'd186,8'd90} : s = 56;
	{8'd186,8'd91} : s = 172;
	{8'd186,8'd92} : s = 170;
	{8'd186,8'd93} : s = 313;
	{8'd186,8'd94} : s = 52;
	{8'd186,8'd95} : s = 169;
	{8'd186,8'd96} : s = 166;
	{8'd186,8'd97} : s = 310;
	{8'd186,8'd98} : s = 165;
	{8'd186,8'd99} : s = 309;
	{8'd186,8'd100} : s = 307;
	{8'd186,8'd101} : s = 427;
	{8'd186,8'd102} : s = 6;
	{8'd186,8'd103} : s = 50;
	{8'd186,8'd104} : s = 49;
	{8'd186,8'd105} : s = 163;
	{8'd186,8'd106} : s = 44;
	{8'd186,8'd107} : s = 156;
	{8'd186,8'd108} : s = 154;
	{8'd186,8'd109} : s = 302;
	{8'd186,8'd110} : s = 42;
	{8'd186,8'd111} : s = 153;
	{8'd186,8'd112} : s = 150;
	{8'd186,8'd113} : s = 301;
	{8'd186,8'd114} : s = 149;
	{8'd186,8'd115} : s = 299;
	{8'd186,8'd116} : s = 295;
	{8'd186,8'd117} : s = 423;
	{8'd186,8'd118} : s = 41;
	{8'd186,8'd119} : s = 147;
	{8'd186,8'd120} : s = 142;
	{8'd186,8'd121} : s = 286;
	{8'd186,8'd122} : s = 141;
	{8'd186,8'd123} : s = 285;
	{8'd186,8'd124} : s = 283;
	{8'd186,8'd125} : s = 414;
	{8'd186,8'd126} : s = 139;
	{8'd186,8'd127} : s = 279;
	{8'd186,8'd128} : s = 271;
	{8'd186,8'd129} : s = 413;
	{8'd186,8'd130} : s = 248;
	{8'd186,8'd131} : s = 411;
	{8'd186,8'd132} : s = 407;
	{8'd186,8'd133} : s = 491;
	{8'd186,8'd134} : s = 5;
	{8'd186,8'd135} : s = 38;
	{8'd186,8'd136} : s = 37;
	{8'd186,8'd137} : s = 135;
	{8'd186,8'd138} : s = 35;
	{8'd186,8'd139} : s = 120;
	{8'd186,8'd140} : s = 116;
	{8'd186,8'd141} : s = 244;
	{8'd186,8'd142} : s = 28;
	{8'd186,8'd143} : s = 114;
	{8'd186,8'd144} : s = 113;
	{8'd186,8'd145} : s = 242;
	{8'd186,8'd146} : s = 108;
	{8'd186,8'd147} : s = 241;
	{8'd186,8'd148} : s = 236;
	{8'd186,8'd149} : s = 399;
	{8'd186,8'd150} : s = 26;
	{8'd186,8'd151} : s = 106;
	{8'd186,8'd152} : s = 105;
	{8'd186,8'd153} : s = 234;
	{8'd186,8'd154} : s = 102;
	{8'd186,8'd155} : s = 233;
	{8'd186,8'd156} : s = 230;
	{8'd186,8'd157} : s = 380;
	{8'd186,8'd158} : s = 101;
	{8'd186,8'd159} : s = 229;
	{8'd186,8'd160} : s = 227;
	{8'd186,8'd161} : s = 378;
	{8'd186,8'd162} : s = 220;
	{8'd186,8'd163} : s = 377;
	{8'd186,8'd164} : s = 374;
	{8'd186,8'd165} : s = 487;
	{8'd186,8'd166} : s = 25;
	{8'd186,8'd167} : s = 99;
	{8'd186,8'd168} : s = 92;
	{8'd186,8'd169} : s = 218;
	{8'd186,8'd170} : s = 90;
	{8'd186,8'd171} : s = 217;
	{8'd186,8'd172} : s = 214;
	{8'd186,8'd173} : s = 373;
	{8'd186,8'd174} : s = 89;
	{8'd186,8'd175} : s = 213;
	{8'd186,8'd176} : s = 211;
	{8'd186,8'd177} : s = 371;
	{8'd186,8'd178} : s = 206;
	{8'd186,8'd179} : s = 366;
	{8'd186,8'd180} : s = 365;
	{8'd186,8'd181} : s = 478;
	{8'd186,8'd182} : s = 86;
	{8'd186,8'd183} : s = 205;
	{8'd186,8'd184} : s = 203;
	{8'd186,8'd185} : s = 363;
	{8'd186,8'd186} : s = 199;
	{8'd186,8'd187} : s = 359;
	{8'd186,8'd188} : s = 350;
	{8'd186,8'd189} : s = 477;
	{8'd186,8'd190} : s = 188;
	{8'd186,8'd191} : s = 349;
	{8'd186,8'd192} : s = 347;
	{8'd186,8'd193} : s = 475;
	{8'd186,8'd194} : s = 343;
	{8'd186,8'd195} : s = 471;
	{8'd186,8'd196} : s = 463;
	{8'd186,8'd197} : s = 509;
	{8'd186,8'd198} : s = 3;
	{8'd186,8'd199} : s = 22;
	{8'd186,8'd200} : s = 21;
	{8'd186,8'd201} : s = 85;
	{8'd186,8'd202} : s = 19;
	{8'd186,8'd203} : s = 83;
	{8'd186,8'd204} : s = 78;
	{8'd186,8'd205} : s = 186;
	{8'd186,8'd206} : s = 14;
	{8'd186,8'd207} : s = 77;
	{8'd186,8'd208} : s = 75;
	{8'd186,8'd209} : s = 185;
	{8'd186,8'd210} : s = 71;
	{8'd186,8'd211} : s = 182;
	{8'd186,8'd212} : s = 181;
	{8'd186,8'd213} : s = 335;
	{8'd186,8'd214} : s = 13;
	{8'd186,8'd215} : s = 60;
	{8'd186,8'd216} : s = 58;
	{8'd186,8'd217} : s = 179;
	{8'd186,8'd218} : s = 57;
	{8'd186,8'd219} : s = 174;
	{8'd186,8'd220} : s = 173;
	{8'd186,8'd221} : s = 318;
	{8'd186,8'd222} : s = 54;
	{8'd186,8'd223} : s = 171;
	{8'd186,8'd224} : s = 167;
	{8'd186,8'd225} : s = 317;
	{8'd186,8'd226} : s = 158;
	{8'd186,8'd227} : s = 315;
	{8'd186,8'd228} : s = 311;
	{8'd186,8'd229} : s = 446;
	{8'd186,8'd230} : s = 11;
	{8'd186,8'd231} : s = 53;
	{8'd186,8'd232} : s = 51;
	{8'd186,8'd233} : s = 157;
	{8'd186,8'd234} : s = 46;
	{8'd186,8'd235} : s = 155;
	{8'd186,8'd236} : s = 151;
	{8'd186,8'd237} : s = 303;
	{8'd186,8'd238} : s = 45;
	{8'd186,8'd239} : s = 143;
	{8'd186,8'd240} : s = 124;
	{8'd186,8'd241} : s = 287;
	{8'd186,8'd242} : s = 122;
	{8'd186,8'd243} : s = 252;
	{8'd186,8'd244} : s = 250;
	{8'd186,8'd245} : s = 445;
	{8'd186,8'd246} : s = 43;
	{8'd186,8'd247} : s = 121;
	{8'd186,8'd248} : s = 118;
	{8'd186,8'd249} : s = 249;
	{8'd186,8'd250} : s = 117;
	{8'd186,8'd251} : s = 246;
	{8'd186,8'd252} : s = 245;
	{8'd186,8'd253} : s = 443;
	{8'd186,8'd254} : s = 115;
	{8'd186,8'd255} : s = 243;
	{8'd187,8'd0} : s = 476;
	{8'd187,8'd1} : s = 376;
	{8'd187,8'd2} : s = 474;
	{8'd187,8'd3} : s = 473;
	{8'd187,8'd4} : s = 506;
	{8'd187,8'd5} : s = 20;
	{8'd187,8'd6} : s = 104;
	{8'd187,8'd7} : s = 100;
	{8'd187,8'd8} : s = 263;
	{8'd187,8'd9} : s = 98;
	{8'd187,8'd10} : s = 240;
	{8'd187,8'd11} : s = 232;
	{8'd187,8'd12} : s = 372;
	{8'd187,8'd13} : s = 97;
	{8'd187,8'd14} : s = 228;
	{8'd187,8'd15} : s = 226;
	{8'd187,8'd16} : s = 370;
	{8'd187,8'd17} : s = 225;
	{8'd187,8'd18} : s = 369;
	{8'd187,8'd19} : s = 364;
	{8'd187,8'd20} : s = 470;
	{8'd187,8'd21} : s = 88;
	{8'd187,8'd22} : s = 216;
	{8'd187,8'd23} : s = 212;
	{8'd187,8'd24} : s = 362;
	{8'd187,8'd25} : s = 210;
	{8'd187,8'd26} : s = 361;
	{8'd187,8'd27} : s = 358;
	{8'd187,8'd28} : s = 469;
	{8'd187,8'd29} : s = 209;
	{8'd187,8'd30} : s = 357;
	{8'd187,8'd31} : s = 355;
	{8'd187,8'd32} : s = 467;
	{8'd187,8'd33} : s = 348;
	{8'd187,8'd34} : s = 462;
	{8'd187,8'd35} : s = 461;
	{8'd187,8'd36} : s = 505;
	{8'd187,8'd37} : s = 84;
	{8'd187,8'd38} : s = 204;
	{8'd187,8'd39} : s = 202;
	{8'd187,8'd40} : s = 346;
	{8'd187,8'd41} : s = 201;
	{8'd187,8'd42} : s = 345;
	{8'd187,8'd43} : s = 342;
	{8'd187,8'd44} : s = 459;
	{8'd187,8'd45} : s = 198;
	{8'd187,8'd46} : s = 341;
	{8'd187,8'd47} : s = 339;
	{8'd187,8'd48} : s = 455;
	{8'd187,8'd49} : s = 334;
	{8'd187,8'd50} : s = 444;
	{8'd187,8'd51} : s = 442;
	{8'd187,8'd52} : s = 502;
	{8'd187,8'd53} : s = 197;
	{8'd187,8'd54} : s = 333;
	{8'd187,8'd55} : s = 331;
	{8'd187,8'd56} : s = 441;
	{8'd187,8'd57} : s = 327;
	{8'd187,8'd58} : s = 438;
	{8'd187,8'd59} : s = 437;
	{8'd187,8'd60} : s = 501;
	{8'd187,8'd61} : s = 316;
	{8'd187,8'd62} : s = 435;
	{8'd187,8'd63} : s = 430;
	{8'd187,8'd64} : s = 499;
	{8'd187,8'd65} : s = 429;
	{8'd187,8'd66} : s = 494;
	{8'd187,8'd67} : s = 493;
	{8'd187,8'd68} : s = 510;
	{8'd187,8'd69} : s = 1;
	{8'd187,8'd70} : s = 18;
	{8'd187,8'd71} : s = 17;
	{8'd187,8'd72} : s = 82;
	{8'd187,8'd73} : s = 12;
	{8'd187,8'd74} : s = 81;
	{8'd187,8'd75} : s = 76;
	{8'd187,8'd76} : s = 195;
	{8'd187,8'd77} : s = 10;
	{8'd187,8'd78} : s = 74;
	{8'd187,8'd79} : s = 73;
	{8'd187,8'd80} : s = 184;
	{8'd187,8'd81} : s = 70;
	{8'd187,8'd82} : s = 180;
	{8'd187,8'd83} : s = 178;
	{8'd187,8'd84} : s = 314;
	{8'd187,8'd85} : s = 9;
	{8'd187,8'd86} : s = 69;
	{8'd187,8'd87} : s = 67;
	{8'd187,8'd88} : s = 177;
	{8'd187,8'd89} : s = 56;
	{8'd187,8'd90} : s = 172;
	{8'd187,8'd91} : s = 170;
	{8'd187,8'd92} : s = 313;
	{8'd187,8'd93} : s = 52;
	{8'd187,8'd94} : s = 169;
	{8'd187,8'd95} : s = 166;
	{8'd187,8'd96} : s = 310;
	{8'd187,8'd97} : s = 165;
	{8'd187,8'd98} : s = 309;
	{8'd187,8'd99} : s = 307;
	{8'd187,8'd100} : s = 427;
	{8'd187,8'd101} : s = 6;
	{8'd187,8'd102} : s = 50;
	{8'd187,8'd103} : s = 49;
	{8'd187,8'd104} : s = 163;
	{8'd187,8'd105} : s = 44;
	{8'd187,8'd106} : s = 156;
	{8'd187,8'd107} : s = 154;
	{8'd187,8'd108} : s = 302;
	{8'd187,8'd109} : s = 42;
	{8'd187,8'd110} : s = 153;
	{8'd187,8'd111} : s = 150;
	{8'd187,8'd112} : s = 301;
	{8'd187,8'd113} : s = 149;
	{8'd187,8'd114} : s = 299;
	{8'd187,8'd115} : s = 295;
	{8'd187,8'd116} : s = 423;
	{8'd187,8'd117} : s = 41;
	{8'd187,8'd118} : s = 147;
	{8'd187,8'd119} : s = 142;
	{8'd187,8'd120} : s = 286;
	{8'd187,8'd121} : s = 141;
	{8'd187,8'd122} : s = 285;
	{8'd187,8'd123} : s = 283;
	{8'd187,8'd124} : s = 414;
	{8'd187,8'd125} : s = 139;
	{8'd187,8'd126} : s = 279;
	{8'd187,8'd127} : s = 271;
	{8'd187,8'd128} : s = 413;
	{8'd187,8'd129} : s = 248;
	{8'd187,8'd130} : s = 411;
	{8'd187,8'd131} : s = 407;
	{8'd187,8'd132} : s = 491;
	{8'd187,8'd133} : s = 5;
	{8'd187,8'd134} : s = 38;
	{8'd187,8'd135} : s = 37;
	{8'd187,8'd136} : s = 135;
	{8'd187,8'd137} : s = 35;
	{8'd187,8'd138} : s = 120;
	{8'd187,8'd139} : s = 116;
	{8'd187,8'd140} : s = 244;
	{8'd187,8'd141} : s = 28;
	{8'd187,8'd142} : s = 114;
	{8'd187,8'd143} : s = 113;
	{8'd187,8'd144} : s = 242;
	{8'd187,8'd145} : s = 108;
	{8'd187,8'd146} : s = 241;
	{8'd187,8'd147} : s = 236;
	{8'd187,8'd148} : s = 399;
	{8'd187,8'd149} : s = 26;
	{8'd187,8'd150} : s = 106;
	{8'd187,8'd151} : s = 105;
	{8'd187,8'd152} : s = 234;
	{8'd187,8'd153} : s = 102;
	{8'd187,8'd154} : s = 233;
	{8'd187,8'd155} : s = 230;
	{8'd187,8'd156} : s = 380;
	{8'd187,8'd157} : s = 101;
	{8'd187,8'd158} : s = 229;
	{8'd187,8'd159} : s = 227;
	{8'd187,8'd160} : s = 378;
	{8'd187,8'd161} : s = 220;
	{8'd187,8'd162} : s = 377;
	{8'd187,8'd163} : s = 374;
	{8'd187,8'd164} : s = 487;
	{8'd187,8'd165} : s = 25;
	{8'd187,8'd166} : s = 99;
	{8'd187,8'd167} : s = 92;
	{8'd187,8'd168} : s = 218;
	{8'd187,8'd169} : s = 90;
	{8'd187,8'd170} : s = 217;
	{8'd187,8'd171} : s = 214;
	{8'd187,8'd172} : s = 373;
	{8'd187,8'd173} : s = 89;
	{8'd187,8'd174} : s = 213;
	{8'd187,8'd175} : s = 211;
	{8'd187,8'd176} : s = 371;
	{8'd187,8'd177} : s = 206;
	{8'd187,8'd178} : s = 366;
	{8'd187,8'd179} : s = 365;
	{8'd187,8'd180} : s = 478;
	{8'd187,8'd181} : s = 86;
	{8'd187,8'd182} : s = 205;
	{8'd187,8'd183} : s = 203;
	{8'd187,8'd184} : s = 363;
	{8'd187,8'd185} : s = 199;
	{8'd187,8'd186} : s = 359;
	{8'd187,8'd187} : s = 350;
	{8'd187,8'd188} : s = 477;
	{8'd187,8'd189} : s = 188;
	{8'd187,8'd190} : s = 349;
	{8'd187,8'd191} : s = 347;
	{8'd187,8'd192} : s = 475;
	{8'd187,8'd193} : s = 343;
	{8'd187,8'd194} : s = 471;
	{8'd187,8'd195} : s = 463;
	{8'd187,8'd196} : s = 509;
	{8'd187,8'd197} : s = 3;
	{8'd187,8'd198} : s = 22;
	{8'd187,8'd199} : s = 21;
	{8'd187,8'd200} : s = 85;
	{8'd187,8'd201} : s = 19;
	{8'd187,8'd202} : s = 83;
	{8'd187,8'd203} : s = 78;
	{8'd187,8'd204} : s = 186;
	{8'd187,8'd205} : s = 14;
	{8'd187,8'd206} : s = 77;
	{8'd187,8'd207} : s = 75;
	{8'd187,8'd208} : s = 185;
	{8'd187,8'd209} : s = 71;
	{8'd187,8'd210} : s = 182;
	{8'd187,8'd211} : s = 181;
	{8'd187,8'd212} : s = 335;
	{8'd187,8'd213} : s = 13;
	{8'd187,8'd214} : s = 60;
	{8'd187,8'd215} : s = 58;
	{8'd187,8'd216} : s = 179;
	{8'd187,8'd217} : s = 57;
	{8'd187,8'd218} : s = 174;
	{8'd187,8'd219} : s = 173;
	{8'd187,8'd220} : s = 318;
	{8'd187,8'd221} : s = 54;
	{8'd187,8'd222} : s = 171;
	{8'd187,8'd223} : s = 167;
	{8'd187,8'd224} : s = 317;
	{8'd187,8'd225} : s = 158;
	{8'd187,8'd226} : s = 315;
	{8'd187,8'd227} : s = 311;
	{8'd187,8'd228} : s = 446;
	{8'd187,8'd229} : s = 11;
	{8'd187,8'd230} : s = 53;
	{8'd187,8'd231} : s = 51;
	{8'd187,8'd232} : s = 157;
	{8'd187,8'd233} : s = 46;
	{8'd187,8'd234} : s = 155;
	{8'd187,8'd235} : s = 151;
	{8'd187,8'd236} : s = 303;
	{8'd187,8'd237} : s = 45;
	{8'd187,8'd238} : s = 143;
	{8'd187,8'd239} : s = 124;
	{8'd187,8'd240} : s = 287;
	{8'd187,8'd241} : s = 122;
	{8'd187,8'd242} : s = 252;
	{8'd187,8'd243} : s = 250;
	{8'd187,8'd244} : s = 445;
	{8'd187,8'd245} : s = 43;
	{8'd187,8'd246} : s = 121;
	{8'd187,8'd247} : s = 118;
	{8'd187,8'd248} : s = 249;
	{8'd187,8'd249} : s = 117;
	{8'd187,8'd250} : s = 246;
	{8'd187,8'd251} : s = 245;
	{8'd187,8'd252} : s = 443;
	{8'd187,8'd253} : s = 115;
	{8'd187,8'd254} : s = 243;
	{8'd187,8'd255} : s = 238;
	{8'd188,8'd0} : s = 376;
	{8'd188,8'd1} : s = 474;
	{8'd188,8'd2} : s = 473;
	{8'd188,8'd3} : s = 506;
	{8'd188,8'd4} : s = 20;
	{8'd188,8'd5} : s = 104;
	{8'd188,8'd6} : s = 100;
	{8'd188,8'd7} : s = 263;
	{8'd188,8'd8} : s = 98;
	{8'd188,8'd9} : s = 240;
	{8'd188,8'd10} : s = 232;
	{8'd188,8'd11} : s = 372;
	{8'd188,8'd12} : s = 97;
	{8'd188,8'd13} : s = 228;
	{8'd188,8'd14} : s = 226;
	{8'd188,8'd15} : s = 370;
	{8'd188,8'd16} : s = 225;
	{8'd188,8'd17} : s = 369;
	{8'd188,8'd18} : s = 364;
	{8'd188,8'd19} : s = 470;
	{8'd188,8'd20} : s = 88;
	{8'd188,8'd21} : s = 216;
	{8'd188,8'd22} : s = 212;
	{8'd188,8'd23} : s = 362;
	{8'd188,8'd24} : s = 210;
	{8'd188,8'd25} : s = 361;
	{8'd188,8'd26} : s = 358;
	{8'd188,8'd27} : s = 469;
	{8'd188,8'd28} : s = 209;
	{8'd188,8'd29} : s = 357;
	{8'd188,8'd30} : s = 355;
	{8'd188,8'd31} : s = 467;
	{8'd188,8'd32} : s = 348;
	{8'd188,8'd33} : s = 462;
	{8'd188,8'd34} : s = 461;
	{8'd188,8'd35} : s = 505;
	{8'd188,8'd36} : s = 84;
	{8'd188,8'd37} : s = 204;
	{8'd188,8'd38} : s = 202;
	{8'd188,8'd39} : s = 346;
	{8'd188,8'd40} : s = 201;
	{8'd188,8'd41} : s = 345;
	{8'd188,8'd42} : s = 342;
	{8'd188,8'd43} : s = 459;
	{8'd188,8'd44} : s = 198;
	{8'd188,8'd45} : s = 341;
	{8'd188,8'd46} : s = 339;
	{8'd188,8'd47} : s = 455;
	{8'd188,8'd48} : s = 334;
	{8'd188,8'd49} : s = 444;
	{8'd188,8'd50} : s = 442;
	{8'd188,8'd51} : s = 502;
	{8'd188,8'd52} : s = 197;
	{8'd188,8'd53} : s = 333;
	{8'd188,8'd54} : s = 331;
	{8'd188,8'd55} : s = 441;
	{8'd188,8'd56} : s = 327;
	{8'd188,8'd57} : s = 438;
	{8'd188,8'd58} : s = 437;
	{8'd188,8'd59} : s = 501;
	{8'd188,8'd60} : s = 316;
	{8'd188,8'd61} : s = 435;
	{8'd188,8'd62} : s = 430;
	{8'd188,8'd63} : s = 499;
	{8'd188,8'd64} : s = 429;
	{8'd188,8'd65} : s = 494;
	{8'd188,8'd66} : s = 493;
	{8'd188,8'd67} : s = 510;
	{8'd188,8'd68} : s = 1;
	{8'd188,8'd69} : s = 18;
	{8'd188,8'd70} : s = 17;
	{8'd188,8'd71} : s = 82;
	{8'd188,8'd72} : s = 12;
	{8'd188,8'd73} : s = 81;
	{8'd188,8'd74} : s = 76;
	{8'd188,8'd75} : s = 195;
	{8'd188,8'd76} : s = 10;
	{8'd188,8'd77} : s = 74;
	{8'd188,8'd78} : s = 73;
	{8'd188,8'd79} : s = 184;
	{8'd188,8'd80} : s = 70;
	{8'd188,8'd81} : s = 180;
	{8'd188,8'd82} : s = 178;
	{8'd188,8'd83} : s = 314;
	{8'd188,8'd84} : s = 9;
	{8'd188,8'd85} : s = 69;
	{8'd188,8'd86} : s = 67;
	{8'd188,8'd87} : s = 177;
	{8'd188,8'd88} : s = 56;
	{8'd188,8'd89} : s = 172;
	{8'd188,8'd90} : s = 170;
	{8'd188,8'd91} : s = 313;
	{8'd188,8'd92} : s = 52;
	{8'd188,8'd93} : s = 169;
	{8'd188,8'd94} : s = 166;
	{8'd188,8'd95} : s = 310;
	{8'd188,8'd96} : s = 165;
	{8'd188,8'd97} : s = 309;
	{8'd188,8'd98} : s = 307;
	{8'd188,8'd99} : s = 427;
	{8'd188,8'd100} : s = 6;
	{8'd188,8'd101} : s = 50;
	{8'd188,8'd102} : s = 49;
	{8'd188,8'd103} : s = 163;
	{8'd188,8'd104} : s = 44;
	{8'd188,8'd105} : s = 156;
	{8'd188,8'd106} : s = 154;
	{8'd188,8'd107} : s = 302;
	{8'd188,8'd108} : s = 42;
	{8'd188,8'd109} : s = 153;
	{8'd188,8'd110} : s = 150;
	{8'd188,8'd111} : s = 301;
	{8'd188,8'd112} : s = 149;
	{8'd188,8'd113} : s = 299;
	{8'd188,8'd114} : s = 295;
	{8'd188,8'd115} : s = 423;
	{8'd188,8'd116} : s = 41;
	{8'd188,8'd117} : s = 147;
	{8'd188,8'd118} : s = 142;
	{8'd188,8'd119} : s = 286;
	{8'd188,8'd120} : s = 141;
	{8'd188,8'd121} : s = 285;
	{8'd188,8'd122} : s = 283;
	{8'd188,8'd123} : s = 414;
	{8'd188,8'd124} : s = 139;
	{8'd188,8'd125} : s = 279;
	{8'd188,8'd126} : s = 271;
	{8'd188,8'd127} : s = 413;
	{8'd188,8'd128} : s = 248;
	{8'd188,8'd129} : s = 411;
	{8'd188,8'd130} : s = 407;
	{8'd188,8'd131} : s = 491;
	{8'd188,8'd132} : s = 5;
	{8'd188,8'd133} : s = 38;
	{8'd188,8'd134} : s = 37;
	{8'd188,8'd135} : s = 135;
	{8'd188,8'd136} : s = 35;
	{8'd188,8'd137} : s = 120;
	{8'd188,8'd138} : s = 116;
	{8'd188,8'd139} : s = 244;
	{8'd188,8'd140} : s = 28;
	{8'd188,8'd141} : s = 114;
	{8'd188,8'd142} : s = 113;
	{8'd188,8'd143} : s = 242;
	{8'd188,8'd144} : s = 108;
	{8'd188,8'd145} : s = 241;
	{8'd188,8'd146} : s = 236;
	{8'd188,8'd147} : s = 399;
	{8'd188,8'd148} : s = 26;
	{8'd188,8'd149} : s = 106;
	{8'd188,8'd150} : s = 105;
	{8'd188,8'd151} : s = 234;
	{8'd188,8'd152} : s = 102;
	{8'd188,8'd153} : s = 233;
	{8'd188,8'd154} : s = 230;
	{8'd188,8'd155} : s = 380;
	{8'd188,8'd156} : s = 101;
	{8'd188,8'd157} : s = 229;
	{8'd188,8'd158} : s = 227;
	{8'd188,8'd159} : s = 378;
	{8'd188,8'd160} : s = 220;
	{8'd188,8'd161} : s = 377;
	{8'd188,8'd162} : s = 374;
	{8'd188,8'd163} : s = 487;
	{8'd188,8'd164} : s = 25;
	{8'd188,8'd165} : s = 99;
	{8'd188,8'd166} : s = 92;
	{8'd188,8'd167} : s = 218;
	{8'd188,8'd168} : s = 90;
	{8'd188,8'd169} : s = 217;
	{8'd188,8'd170} : s = 214;
	{8'd188,8'd171} : s = 373;
	{8'd188,8'd172} : s = 89;
	{8'd188,8'd173} : s = 213;
	{8'd188,8'd174} : s = 211;
	{8'd188,8'd175} : s = 371;
	{8'd188,8'd176} : s = 206;
	{8'd188,8'd177} : s = 366;
	{8'd188,8'd178} : s = 365;
	{8'd188,8'd179} : s = 478;
	{8'd188,8'd180} : s = 86;
	{8'd188,8'd181} : s = 205;
	{8'd188,8'd182} : s = 203;
	{8'd188,8'd183} : s = 363;
	{8'd188,8'd184} : s = 199;
	{8'd188,8'd185} : s = 359;
	{8'd188,8'd186} : s = 350;
	{8'd188,8'd187} : s = 477;
	{8'd188,8'd188} : s = 188;
	{8'd188,8'd189} : s = 349;
	{8'd188,8'd190} : s = 347;
	{8'd188,8'd191} : s = 475;
	{8'd188,8'd192} : s = 343;
	{8'd188,8'd193} : s = 471;
	{8'd188,8'd194} : s = 463;
	{8'd188,8'd195} : s = 509;
	{8'd188,8'd196} : s = 3;
	{8'd188,8'd197} : s = 22;
	{8'd188,8'd198} : s = 21;
	{8'd188,8'd199} : s = 85;
	{8'd188,8'd200} : s = 19;
	{8'd188,8'd201} : s = 83;
	{8'd188,8'd202} : s = 78;
	{8'd188,8'd203} : s = 186;
	{8'd188,8'd204} : s = 14;
	{8'd188,8'd205} : s = 77;
	{8'd188,8'd206} : s = 75;
	{8'd188,8'd207} : s = 185;
	{8'd188,8'd208} : s = 71;
	{8'd188,8'd209} : s = 182;
	{8'd188,8'd210} : s = 181;
	{8'd188,8'd211} : s = 335;
	{8'd188,8'd212} : s = 13;
	{8'd188,8'd213} : s = 60;
	{8'd188,8'd214} : s = 58;
	{8'd188,8'd215} : s = 179;
	{8'd188,8'd216} : s = 57;
	{8'd188,8'd217} : s = 174;
	{8'd188,8'd218} : s = 173;
	{8'd188,8'd219} : s = 318;
	{8'd188,8'd220} : s = 54;
	{8'd188,8'd221} : s = 171;
	{8'd188,8'd222} : s = 167;
	{8'd188,8'd223} : s = 317;
	{8'd188,8'd224} : s = 158;
	{8'd188,8'd225} : s = 315;
	{8'd188,8'd226} : s = 311;
	{8'd188,8'd227} : s = 446;
	{8'd188,8'd228} : s = 11;
	{8'd188,8'd229} : s = 53;
	{8'd188,8'd230} : s = 51;
	{8'd188,8'd231} : s = 157;
	{8'd188,8'd232} : s = 46;
	{8'd188,8'd233} : s = 155;
	{8'd188,8'd234} : s = 151;
	{8'd188,8'd235} : s = 303;
	{8'd188,8'd236} : s = 45;
	{8'd188,8'd237} : s = 143;
	{8'd188,8'd238} : s = 124;
	{8'd188,8'd239} : s = 287;
	{8'd188,8'd240} : s = 122;
	{8'd188,8'd241} : s = 252;
	{8'd188,8'd242} : s = 250;
	{8'd188,8'd243} : s = 445;
	{8'd188,8'd244} : s = 43;
	{8'd188,8'd245} : s = 121;
	{8'd188,8'd246} : s = 118;
	{8'd188,8'd247} : s = 249;
	{8'd188,8'd248} : s = 117;
	{8'd188,8'd249} : s = 246;
	{8'd188,8'd250} : s = 245;
	{8'd188,8'd251} : s = 443;
	{8'd188,8'd252} : s = 115;
	{8'd188,8'd253} : s = 243;
	{8'd188,8'd254} : s = 238;
	{8'd188,8'd255} : s = 439;
	{8'd189,8'd0} : s = 474;
	{8'd189,8'd1} : s = 473;
	{8'd189,8'd2} : s = 506;
	{8'd189,8'd3} : s = 20;
	{8'd189,8'd4} : s = 104;
	{8'd189,8'd5} : s = 100;
	{8'd189,8'd6} : s = 263;
	{8'd189,8'd7} : s = 98;
	{8'd189,8'd8} : s = 240;
	{8'd189,8'd9} : s = 232;
	{8'd189,8'd10} : s = 372;
	{8'd189,8'd11} : s = 97;
	{8'd189,8'd12} : s = 228;
	{8'd189,8'd13} : s = 226;
	{8'd189,8'd14} : s = 370;
	{8'd189,8'd15} : s = 225;
	{8'd189,8'd16} : s = 369;
	{8'd189,8'd17} : s = 364;
	{8'd189,8'd18} : s = 470;
	{8'd189,8'd19} : s = 88;
	{8'd189,8'd20} : s = 216;
	{8'd189,8'd21} : s = 212;
	{8'd189,8'd22} : s = 362;
	{8'd189,8'd23} : s = 210;
	{8'd189,8'd24} : s = 361;
	{8'd189,8'd25} : s = 358;
	{8'd189,8'd26} : s = 469;
	{8'd189,8'd27} : s = 209;
	{8'd189,8'd28} : s = 357;
	{8'd189,8'd29} : s = 355;
	{8'd189,8'd30} : s = 467;
	{8'd189,8'd31} : s = 348;
	{8'd189,8'd32} : s = 462;
	{8'd189,8'd33} : s = 461;
	{8'd189,8'd34} : s = 505;
	{8'd189,8'd35} : s = 84;
	{8'd189,8'd36} : s = 204;
	{8'd189,8'd37} : s = 202;
	{8'd189,8'd38} : s = 346;
	{8'd189,8'd39} : s = 201;
	{8'd189,8'd40} : s = 345;
	{8'd189,8'd41} : s = 342;
	{8'd189,8'd42} : s = 459;
	{8'd189,8'd43} : s = 198;
	{8'd189,8'd44} : s = 341;
	{8'd189,8'd45} : s = 339;
	{8'd189,8'd46} : s = 455;
	{8'd189,8'd47} : s = 334;
	{8'd189,8'd48} : s = 444;
	{8'd189,8'd49} : s = 442;
	{8'd189,8'd50} : s = 502;
	{8'd189,8'd51} : s = 197;
	{8'd189,8'd52} : s = 333;
	{8'd189,8'd53} : s = 331;
	{8'd189,8'd54} : s = 441;
	{8'd189,8'd55} : s = 327;
	{8'd189,8'd56} : s = 438;
	{8'd189,8'd57} : s = 437;
	{8'd189,8'd58} : s = 501;
	{8'd189,8'd59} : s = 316;
	{8'd189,8'd60} : s = 435;
	{8'd189,8'd61} : s = 430;
	{8'd189,8'd62} : s = 499;
	{8'd189,8'd63} : s = 429;
	{8'd189,8'd64} : s = 494;
	{8'd189,8'd65} : s = 493;
	{8'd189,8'd66} : s = 510;
	{8'd189,8'd67} : s = 1;
	{8'd189,8'd68} : s = 18;
	{8'd189,8'd69} : s = 17;
	{8'd189,8'd70} : s = 82;
	{8'd189,8'd71} : s = 12;
	{8'd189,8'd72} : s = 81;
	{8'd189,8'd73} : s = 76;
	{8'd189,8'd74} : s = 195;
	{8'd189,8'd75} : s = 10;
	{8'd189,8'd76} : s = 74;
	{8'd189,8'd77} : s = 73;
	{8'd189,8'd78} : s = 184;
	{8'd189,8'd79} : s = 70;
	{8'd189,8'd80} : s = 180;
	{8'd189,8'd81} : s = 178;
	{8'd189,8'd82} : s = 314;
	{8'd189,8'd83} : s = 9;
	{8'd189,8'd84} : s = 69;
	{8'd189,8'd85} : s = 67;
	{8'd189,8'd86} : s = 177;
	{8'd189,8'd87} : s = 56;
	{8'd189,8'd88} : s = 172;
	{8'd189,8'd89} : s = 170;
	{8'd189,8'd90} : s = 313;
	{8'd189,8'd91} : s = 52;
	{8'd189,8'd92} : s = 169;
	{8'd189,8'd93} : s = 166;
	{8'd189,8'd94} : s = 310;
	{8'd189,8'd95} : s = 165;
	{8'd189,8'd96} : s = 309;
	{8'd189,8'd97} : s = 307;
	{8'd189,8'd98} : s = 427;
	{8'd189,8'd99} : s = 6;
	{8'd189,8'd100} : s = 50;
	{8'd189,8'd101} : s = 49;
	{8'd189,8'd102} : s = 163;
	{8'd189,8'd103} : s = 44;
	{8'd189,8'd104} : s = 156;
	{8'd189,8'd105} : s = 154;
	{8'd189,8'd106} : s = 302;
	{8'd189,8'd107} : s = 42;
	{8'd189,8'd108} : s = 153;
	{8'd189,8'd109} : s = 150;
	{8'd189,8'd110} : s = 301;
	{8'd189,8'd111} : s = 149;
	{8'd189,8'd112} : s = 299;
	{8'd189,8'd113} : s = 295;
	{8'd189,8'd114} : s = 423;
	{8'd189,8'd115} : s = 41;
	{8'd189,8'd116} : s = 147;
	{8'd189,8'd117} : s = 142;
	{8'd189,8'd118} : s = 286;
	{8'd189,8'd119} : s = 141;
	{8'd189,8'd120} : s = 285;
	{8'd189,8'd121} : s = 283;
	{8'd189,8'd122} : s = 414;
	{8'd189,8'd123} : s = 139;
	{8'd189,8'd124} : s = 279;
	{8'd189,8'd125} : s = 271;
	{8'd189,8'd126} : s = 413;
	{8'd189,8'd127} : s = 248;
	{8'd189,8'd128} : s = 411;
	{8'd189,8'd129} : s = 407;
	{8'd189,8'd130} : s = 491;
	{8'd189,8'd131} : s = 5;
	{8'd189,8'd132} : s = 38;
	{8'd189,8'd133} : s = 37;
	{8'd189,8'd134} : s = 135;
	{8'd189,8'd135} : s = 35;
	{8'd189,8'd136} : s = 120;
	{8'd189,8'd137} : s = 116;
	{8'd189,8'd138} : s = 244;
	{8'd189,8'd139} : s = 28;
	{8'd189,8'd140} : s = 114;
	{8'd189,8'd141} : s = 113;
	{8'd189,8'd142} : s = 242;
	{8'd189,8'd143} : s = 108;
	{8'd189,8'd144} : s = 241;
	{8'd189,8'd145} : s = 236;
	{8'd189,8'd146} : s = 399;
	{8'd189,8'd147} : s = 26;
	{8'd189,8'd148} : s = 106;
	{8'd189,8'd149} : s = 105;
	{8'd189,8'd150} : s = 234;
	{8'd189,8'd151} : s = 102;
	{8'd189,8'd152} : s = 233;
	{8'd189,8'd153} : s = 230;
	{8'd189,8'd154} : s = 380;
	{8'd189,8'd155} : s = 101;
	{8'd189,8'd156} : s = 229;
	{8'd189,8'd157} : s = 227;
	{8'd189,8'd158} : s = 378;
	{8'd189,8'd159} : s = 220;
	{8'd189,8'd160} : s = 377;
	{8'd189,8'd161} : s = 374;
	{8'd189,8'd162} : s = 487;
	{8'd189,8'd163} : s = 25;
	{8'd189,8'd164} : s = 99;
	{8'd189,8'd165} : s = 92;
	{8'd189,8'd166} : s = 218;
	{8'd189,8'd167} : s = 90;
	{8'd189,8'd168} : s = 217;
	{8'd189,8'd169} : s = 214;
	{8'd189,8'd170} : s = 373;
	{8'd189,8'd171} : s = 89;
	{8'd189,8'd172} : s = 213;
	{8'd189,8'd173} : s = 211;
	{8'd189,8'd174} : s = 371;
	{8'd189,8'd175} : s = 206;
	{8'd189,8'd176} : s = 366;
	{8'd189,8'd177} : s = 365;
	{8'd189,8'd178} : s = 478;
	{8'd189,8'd179} : s = 86;
	{8'd189,8'd180} : s = 205;
	{8'd189,8'd181} : s = 203;
	{8'd189,8'd182} : s = 363;
	{8'd189,8'd183} : s = 199;
	{8'd189,8'd184} : s = 359;
	{8'd189,8'd185} : s = 350;
	{8'd189,8'd186} : s = 477;
	{8'd189,8'd187} : s = 188;
	{8'd189,8'd188} : s = 349;
	{8'd189,8'd189} : s = 347;
	{8'd189,8'd190} : s = 475;
	{8'd189,8'd191} : s = 343;
	{8'd189,8'd192} : s = 471;
	{8'd189,8'd193} : s = 463;
	{8'd189,8'd194} : s = 509;
	{8'd189,8'd195} : s = 3;
	{8'd189,8'd196} : s = 22;
	{8'd189,8'd197} : s = 21;
	{8'd189,8'd198} : s = 85;
	{8'd189,8'd199} : s = 19;
	{8'd189,8'd200} : s = 83;
	{8'd189,8'd201} : s = 78;
	{8'd189,8'd202} : s = 186;
	{8'd189,8'd203} : s = 14;
	{8'd189,8'd204} : s = 77;
	{8'd189,8'd205} : s = 75;
	{8'd189,8'd206} : s = 185;
	{8'd189,8'd207} : s = 71;
	{8'd189,8'd208} : s = 182;
	{8'd189,8'd209} : s = 181;
	{8'd189,8'd210} : s = 335;
	{8'd189,8'd211} : s = 13;
	{8'd189,8'd212} : s = 60;
	{8'd189,8'd213} : s = 58;
	{8'd189,8'd214} : s = 179;
	{8'd189,8'd215} : s = 57;
	{8'd189,8'd216} : s = 174;
	{8'd189,8'd217} : s = 173;
	{8'd189,8'd218} : s = 318;
	{8'd189,8'd219} : s = 54;
	{8'd189,8'd220} : s = 171;
	{8'd189,8'd221} : s = 167;
	{8'd189,8'd222} : s = 317;
	{8'd189,8'd223} : s = 158;
	{8'd189,8'd224} : s = 315;
	{8'd189,8'd225} : s = 311;
	{8'd189,8'd226} : s = 446;
	{8'd189,8'd227} : s = 11;
	{8'd189,8'd228} : s = 53;
	{8'd189,8'd229} : s = 51;
	{8'd189,8'd230} : s = 157;
	{8'd189,8'd231} : s = 46;
	{8'd189,8'd232} : s = 155;
	{8'd189,8'd233} : s = 151;
	{8'd189,8'd234} : s = 303;
	{8'd189,8'd235} : s = 45;
	{8'd189,8'd236} : s = 143;
	{8'd189,8'd237} : s = 124;
	{8'd189,8'd238} : s = 287;
	{8'd189,8'd239} : s = 122;
	{8'd189,8'd240} : s = 252;
	{8'd189,8'd241} : s = 250;
	{8'd189,8'd242} : s = 445;
	{8'd189,8'd243} : s = 43;
	{8'd189,8'd244} : s = 121;
	{8'd189,8'd245} : s = 118;
	{8'd189,8'd246} : s = 249;
	{8'd189,8'd247} : s = 117;
	{8'd189,8'd248} : s = 246;
	{8'd189,8'd249} : s = 245;
	{8'd189,8'd250} : s = 443;
	{8'd189,8'd251} : s = 115;
	{8'd189,8'd252} : s = 243;
	{8'd189,8'd253} : s = 238;
	{8'd189,8'd254} : s = 439;
	{8'd189,8'd255} : s = 237;
	{8'd190,8'd0} : s = 473;
	{8'd190,8'd1} : s = 506;
	{8'd190,8'd2} : s = 20;
	{8'd190,8'd3} : s = 104;
	{8'd190,8'd4} : s = 100;
	{8'd190,8'd5} : s = 263;
	{8'd190,8'd6} : s = 98;
	{8'd190,8'd7} : s = 240;
	{8'd190,8'd8} : s = 232;
	{8'd190,8'd9} : s = 372;
	{8'd190,8'd10} : s = 97;
	{8'd190,8'd11} : s = 228;
	{8'd190,8'd12} : s = 226;
	{8'd190,8'd13} : s = 370;
	{8'd190,8'd14} : s = 225;
	{8'd190,8'd15} : s = 369;
	{8'd190,8'd16} : s = 364;
	{8'd190,8'd17} : s = 470;
	{8'd190,8'd18} : s = 88;
	{8'd190,8'd19} : s = 216;
	{8'd190,8'd20} : s = 212;
	{8'd190,8'd21} : s = 362;
	{8'd190,8'd22} : s = 210;
	{8'd190,8'd23} : s = 361;
	{8'd190,8'd24} : s = 358;
	{8'd190,8'd25} : s = 469;
	{8'd190,8'd26} : s = 209;
	{8'd190,8'd27} : s = 357;
	{8'd190,8'd28} : s = 355;
	{8'd190,8'd29} : s = 467;
	{8'd190,8'd30} : s = 348;
	{8'd190,8'd31} : s = 462;
	{8'd190,8'd32} : s = 461;
	{8'd190,8'd33} : s = 505;
	{8'd190,8'd34} : s = 84;
	{8'd190,8'd35} : s = 204;
	{8'd190,8'd36} : s = 202;
	{8'd190,8'd37} : s = 346;
	{8'd190,8'd38} : s = 201;
	{8'd190,8'd39} : s = 345;
	{8'd190,8'd40} : s = 342;
	{8'd190,8'd41} : s = 459;
	{8'd190,8'd42} : s = 198;
	{8'd190,8'd43} : s = 341;
	{8'd190,8'd44} : s = 339;
	{8'd190,8'd45} : s = 455;
	{8'd190,8'd46} : s = 334;
	{8'd190,8'd47} : s = 444;
	{8'd190,8'd48} : s = 442;
	{8'd190,8'd49} : s = 502;
	{8'd190,8'd50} : s = 197;
	{8'd190,8'd51} : s = 333;
	{8'd190,8'd52} : s = 331;
	{8'd190,8'd53} : s = 441;
	{8'd190,8'd54} : s = 327;
	{8'd190,8'd55} : s = 438;
	{8'd190,8'd56} : s = 437;
	{8'd190,8'd57} : s = 501;
	{8'd190,8'd58} : s = 316;
	{8'd190,8'd59} : s = 435;
	{8'd190,8'd60} : s = 430;
	{8'd190,8'd61} : s = 499;
	{8'd190,8'd62} : s = 429;
	{8'd190,8'd63} : s = 494;
	{8'd190,8'd64} : s = 493;
	{8'd190,8'd65} : s = 510;
	{8'd190,8'd66} : s = 1;
	{8'd190,8'd67} : s = 18;
	{8'd190,8'd68} : s = 17;
	{8'd190,8'd69} : s = 82;
	{8'd190,8'd70} : s = 12;
	{8'd190,8'd71} : s = 81;
	{8'd190,8'd72} : s = 76;
	{8'd190,8'd73} : s = 195;
	{8'd190,8'd74} : s = 10;
	{8'd190,8'd75} : s = 74;
	{8'd190,8'd76} : s = 73;
	{8'd190,8'd77} : s = 184;
	{8'd190,8'd78} : s = 70;
	{8'd190,8'd79} : s = 180;
	{8'd190,8'd80} : s = 178;
	{8'd190,8'd81} : s = 314;
	{8'd190,8'd82} : s = 9;
	{8'd190,8'd83} : s = 69;
	{8'd190,8'd84} : s = 67;
	{8'd190,8'd85} : s = 177;
	{8'd190,8'd86} : s = 56;
	{8'd190,8'd87} : s = 172;
	{8'd190,8'd88} : s = 170;
	{8'd190,8'd89} : s = 313;
	{8'd190,8'd90} : s = 52;
	{8'd190,8'd91} : s = 169;
	{8'd190,8'd92} : s = 166;
	{8'd190,8'd93} : s = 310;
	{8'd190,8'd94} : s = 165;
	{8'd190,8'd95} : s = 309;
	{8'd190,8'd96} : s = 307;
	{8'd190,8'd97} : s = 427;
	{8'd190,8'd98} : s = 6;
	{8'd190,8'd99} : s = 50;
	{8'd190,8'd100} : s = 49;
	{8'd190,8'd101} : s = 163;
	{8'd190,8'd102} : s = 44;
	{8'd190,8'd103} : s = 156;
	{8'd190,8'd104} : s = 154;
	{8'd190,8'd105} : s = 302;
	{8'd190,8'd106} : s = 42;
	{8'd190,8'd107} : s = 153;
	{8'd190,8'd108} : s = 150;
	{8'd190,8'd109} : s = 301;
	{8'd190,8'd110} : s = 149;
	{8'd190,8'd111} : s = 299;
	{8'd190,8'd112} : s = 295;
	{8'd190,8'd113} : s = 423;
	{8'd190,8'd114} : s = 41;
	{8'd190,8'd115} : s = 147;
	{8'd190,8'd116} : s = 142;
	{8'd190,8'd117} : s = 286;
	{8'd190,8'd118} : s = 141;
	{8'd190,8'd119} : s = 285;
	{8'd190,8'd120} : s = 283;
	{8'd190,8'd121} : s = 414;
	{8'd190,8'd122} : s = 139;
	{8'd190,8'd123} : s = 279;
	{8'd190,8'd124} : s = 271;
	{8'd190,8'd125} : s = 413;
	{8'd190,8'd126} : s = 248;
	{8'd190,8'd127} : s = 411;
	{8'd190,8'd128} : s = 407;
	{8'd190,8'd129} : s = 491;
	{8'd190,8'd130} : s = 5;
	{8'd190,8'd131} : s = 38;
	{8'd190,8'd132} : s = 37;
	{8'd190,8'd133} : s = 135;
	{8'd190,8'd134} : s = 35;
	{8'd190,8'd135} : s = 120;
	{8'd190,8'd136} : s = 116;
	{8'd190,8'd137} : s = 244;
	{8'd190,8'd138} : s = 28;
	{8'd190,8'd139} : s = 114;
	{8'd190,8'd140} : s = 113;
	{8'd190,8'd141} : s = 242;
	{8'd190,8'd142} : s = 108;
	{8'd190,8'd143} : s = 241;
	{8'd190,8'd144} : s = 236;
	{8'd190,8'd145} : s = 399;
	{8'd190,8'd146} : s = 26;
	{8'd190,8'd147} : s = 106;
	{8'd190,8'd148} : s = 105;
	{8'd190,8'd149} : s = 234;
	{8'd190,8'd150} : s = 102;
	{8'd190,8'd151} : s = 233;
	{8'd190,8'd152} : s = 230;
	{8'd190,8'd153} : s = 380;
	{8'd190,8'd154} : s = 101;
	{8'd190,8'd155} : s = 229;
	{8'd190,8'd156} : s = 227;
	{8'd190,8'd157} : s = 378;
	{8'd190,8'd158} : s = 220;
	{8'd190,8'd159} : s = 377;
	{8'd190,8'd160} : s = 374;
	{8'd190,8'd161} : s = 487;
	{8'd190,8'd162} : s = 25;
	{8'd190,8'd163} : s = 99;
	{8'd190,8'd164} : s = 92;
	{8'd190,8'd165} : s = 218;
	{8'd190,8'd166} : s = 90;
	{8'd190,8'd167} : s = 217;
	{8'd190,8'd168} : s = 214;
	{8'd190,8'd169} : s = 373;
	{8'd190,8'd170} : s = 89;
	{8'd190,8'd171} : s = 213;
	{8'd190,8'd172} : s = 211;
	{8'd190,8'd173} : s = 371;
	{8'd190,8'd174} : s = 206;
	{8'd190,8'd175} : s = 366;
	{8'd190,8'd176} : s = 365;
	{8'd190,8'd177} : s = 478;
	{8'd190,8'd178} : s = 86;
	{8'd190,8'd179} : s = 205;
	{8'd190,8'd180} : s = 203;
	{8'd190,8'd181} : s = 363;
	{8'd190,8'd182} : s = 199;
	{8'd190,8'd183} : s = 359;
	{8'd190,8'd184} : s = 350;
	{8'd190,8'd185} : s = 477;
	{8'd190,8'd186} : s = 188;
	{8'd190,8'd187} : s = 349;
	{8'd190,8'd188} : s = 347;
	{8'd190,8'd189} : s = 475;
	{8'd190,8'd190} : s = 343;
	{8'd190,8'd191} : s = 471;
	{8'd190,8'd192} : s = 463;
	{8'd190,8'd193} : s = 509;
	{8'd190,8'd194} : s = 3;
	{8'd190,8'd195} : s = 22;
	{8'd190,8'd196} : s = 21;
	{8'd190,8'd197} : s = 85;
	{8'd190,8'd198} : s = 19;
	{8'd190,8'd199} : s = 83;
	{8'd190,8'd200} : s = 78;
	{8'd190,8'd201} : s = 186;
	{8'd190,8'd202} : s = 14;
	{8'd190,8'd203} : s = 77;
	{8'd190,8'd204} : s = 75;
	{8'd190,8'd205} : s = 185;
	{8'd190,8'd206} : s = 71;
	{8'd190,8'd207} : s = 182;
	{8'd190,8'd208} : s = 181;
	{8'd190,8'd209} : s = 335;
	{8'd190,8'd210} : s = 13;
	{8'd190,8'd211} : s = 60;
	{8'd190,8'd212} : s = 58;
	{8'd190,8'd213} : s = 179;
	{8'd190,8'd214} : s = 57;
	{8'd190,8'd215} : s = 174;
	{8'd190,8'd216} : s = 173;
	{8'd190,8'd217} : s = 318;
	{8'd190,8'd218} : s = 54;
	{8'd190,8'd219} : s = 171;
	{8'd190,8'd220} : s = 167;
	{8'd190,8'd221} : s = 317;
	{8'd190,8'd222} : s = 158;
	{8'd190,8'd223} : s = 315;
	{8'd190,8'd224} : s = 311;
	{8'd190,8'd225} : s = 446;
	{8'd190,8'd226} : s = 11;
	{8'd190,8'd227} : s = 53;
	{8'd190,8'd228} : s = 51;
	{8'd190,8'd229} : s = 157;
	{8'd190,8'd230} : s = 46;
	{8'd190,8'd231} : s = 155;
	{8'd190,8'd232} : s = 151;
	{8'd190,8'd233} : s = 303;
	{8'd190,8'd234} : s = 45;
	{8'd190,8'd235} : s = 143;
	{8'd190,8'd236} : s = 124;
	{8'd190,8'd237} : s = 287;
	{8'd190,8'd238} : s = 122;
	{8'd190,8'd239} : s = 252;
	{8'd190,8'd240} : s = 250;
	{8'd190,8'd241} : s = 445;
	{8'd190,8'd242} : s = 43;
	{8'd190,8'd243} : s = 121;
	{8'd190,8'd244} : s = 118;
	{8'd190,8'd245} : s = 249;
	{8'd190,8'd246} : s = 117;
	{8'd190,8'd247} : s = 246;
	{8'd190,8'd248} : s = 245;
	{8'd190,8'd249} : s = 443;
	{8'd190,8'd250} : s = 115;
	{8'd190,8'd251} : s = 243;
	{8'd190,8'd252} : s = 238;
	{8'd190,8'd253} : s = 439;
	{8'd190,8'd254} : s = 237;
	{8'd190,8'd255} : s = 431;
	{8'd191,8'd0} : s = 506;
	{8'd191,8'd1} : s = 20;
	{8'd191,8'd2} : s = 104;
	{8'd191,8'd3} : s = 100;
	{8'd191,8'd4} : s = 263;
	{8'd191,8'd5} : s = 98;
	{8'd191,8'd6} : s = 240;
	{8'd191,8'd7} : s = 232;
	{8'd191,8'd8} : s = 372;
	{8'd191,8'd9} : s = 97;
	{8'd191,8'd10} : s = 228;
	{8'd191,8'd11} : s = 226;
	{8'd191,8'd12} : s = 370;
	{8'd191,8'd13} : s = 225;
	{8'd191,8'd14} : s = 369;
	{8'd191,8'd15} : s = 364;
	{8'd191,8'd16} : s = 470;
	{8'd191,8'd17} : s = 88;
	{8'd191,8'd18} : s = 216;
	{8'd191,8'd19} : s = 212;
	{8'd191,8'd20} : s = 362;
	{8'd191,8'd21} : s = 210;
	{8'd191,8'd22} : s = 361;
	{8'd191,8'd23} : s = 358;
	{8'd191,8'd24} : s = 469;
	{8'd191,8'd25} : s = 209;
	{8'd191,8'd26} : s = 357;
	{8'd191,8'd27} : s = 355;
	{8'd191,8'd28} : s = 467;
	{8'd191,8'd29} : s = 348;
	{8'd191,8'd30} : s = 462;
	{8'd191,8'd31} : s = 461;
	{8'd191,8'd32} : s = 505;
	{8'd191,8'd33} : s = 84;
	{8'd191,8'd34} : s = 204;
	{8'd191,8'd35} : s = 202;
	{8'd191,8'd36} : s = 346;
	{8'd191,8'd37} : s = 201;
	{8'd191,8'd38} : s = 345;
	{8'd191,8'd39} : s = 342;
	{8'd191,8'd40} : s = 459;
	{8'd191,8'd41} : s = 198;
	{8'd191,8'd42} : s = 341;
	{8'd191,8'd43} : s = 339;
	{8'd191,8'd44} : s = 455;
	{8'd191,8'd45} : s = 334;
	{8'd191,8'd46} : s = 444;
	{8'd191,8'd47} : s = 442;
	{8'd191,8'd48} : s = 502;
	{8'd191,8'd49} : s = 197;
	{8'd191,8'd50} : s = 333;
	{8'd191,8'd51} : s = 331;
	{8'd191,8'd52} : s = 441;
	{8'd191,8'd53} : s = 327;
	{8'd191,8'd54} : s = 438;
	{8'd191,8'd55} : s = 437;
	{8'd191,8'd56} : s = 501;
	{8'd191,8'd57} : s = 316;
	{8'd191,8'd58} : s = 435;
	{8'd191,8'd59} : s = 430;
	{8'd191,8'd60} : s = 499;
	{8'd191,8'd61} : s = 429;
	{8'd191,8'd62} : s = 494;
	{8'd191,8'd63} : s = 493;
	{8'd191,8'd64} : s = 510;
	{8'd191,8'd65} : s = 1;
	{8'd191,8'd66} : s = 18;
	{8'd191,8'd67} : s = 17;
	{8'd191,8'd68} : s = 82;
	{8'd191,8'd69} : s = 12;
	{8'd191,8'd70} : s = 81;
	{8'd191,8'd71} : s = 76;
	{8'd191,8'd72} : s = 195;
	{8'd191,8'd73} : s = 10;
	{8'd191,8'd74} : s = 74;
	{8'd191,8'd75} : s = 73;
	{8'd191,8'd76} : s = 184;
	{8'd191,8'd77} : s = 70;
	{8'd191,8'd78} : s = 180;
	{8'd191,8'd79} : s = 178;
	{8'd191,8'd80} : s = 314;
	{8'd191,8'd81} : s = 9;
	{8'd191,8'd82} : s = 69;
	{8'd191,8'd83} : s = 67;
	{8'd191,8'd84} : s = 177;
	{8'd191,8'd85} : s = 56;
	{8'd191,8'd86} : s = 172;
	{8'd191,8'd87} : s = 170;
	{8'd191,8'd88} : s = 313;
	{8'd191,8'd89} : s = 52;
	{8'd191,8'd90} : s = 169;
	{8'd191,8'd91} : s = 166;
	{8'd191,8'd92} : s = 310;
	{8'd191,8'd93} : s = 165;
	{8'd191,8'd94} : s = 309;
	{8'd191,8'd95} : s = 307;
	{8'd191,8'd96} : s = 427;
	{8'd191,8'd97} : s = 6;
	{8'd191,8'd98} : s = 50;
	{8'd191,8'd99} : s = 49;
	{8'd191,8'd100} : s = 163;
	{8'd191,8'd101} : s = 44;
	{8'd191,8'd102} : s = 156;
	{8'd191,8'd103} : s = 154;
	{8'd191,8'd104} : s = 302;
	{8'd191,8'd105} : s = 42;
	{8'd191,8'd106} : s = 153;
	{8'd191,8'd107} : s = 150;
	{8'd191,8'd108} : s = 301;
	{8'd191,8'd109} : s = 149;
	{8'd191,8'd110} : s = 299;
	{8'd191,8'd111} : s = 295;
	{8'd191,8'd112} : s = 423;
	{8'd191,8'd113} : s = 41;
	{8'd191,8'd114} : s = 147;
	{8'd191,8'd115} : s = 142;
	{8'd191,8'd116} : s = 286;
	{8'd191,8'd117} : s = 141;
	{8'd191,8'd118} : s = 285;
	{8'd191,8'd119} : s = 283;
	{8'd191,8'd120} : s = 414;
	{8'd191,8'd121} : s = 139;
	{8'd191,8'd122} : s = 279;
	{8'd191,8'd123} : s = 271;
	{8'd191,8'd124} : s = 413;
	{8'd191,8'd125} : s = 248;
	{8'd191,8'd126} : s = 411;
	{8'd191,8'd127} : s = 407;
	{8'd191,8'd128} : s = 491;
	{8'd191,8'd129} : s = 5;
	{8'd191,8'd130} : s = 38;
	{8'd191,8'd131} : s = 37;
	{8'd191,8'd132} : s = 135;
	{8'd191,8'd133} : s = 35;
	{8'd191,8'd134} : s = 120;
	{8'd191,8'd135} : s = 116;
	{8'd191,8'd136} : s = 244;
	{8'd191,8'd137} : s = 28;
	{8'd191,8'd138} : s = 114;
	{8'd191,8'd139} : s = 113;
	{8'd191,8'd140} : s = 242;
	{8'd191,8'd141} : s = 108;
	{8'd191,8'd142} : s = 241;
	{8'd191,8'd143} : s = 236;
	{8'd191,8'd144} : s = 399;
	{8'd191,8'd145} : s = 26;
	{8'd191,8'd146} : s = 106;
	{8'd191,8'd147} : s = 105;
	{8'd191,8'd148} : s = 234;
	{8'd191,8'd149} : s = 102;
	{8'd191,8'd150} : s = 233;
	{8'd191,8'd151} : s = 230;
	{8'd191,8'd152} : s = 380;
	{8'd191,8'd153} : s = 101;
	{8'd191,8'd154} : s = 229;
	{8'd191,8'd155} : s = 227;
	{8'd191,8'd156} : s = 378;
	{8'd191,8'd157} : s = 220;
	{8'd191,8'd158} : s = 377;
	{8'd191,8'd159} : s = 374;
	{8'd191,8'd160} : s = 487;
	{8'd191,8'd161} : s = 25;
	{8'd191,8'd162} : s = 99;
	{8'd191,8'd163} : s = 92;
	{8'd191,8'd164} : s = 218;
	{8'd191,8'd165} : s = 90;
	{8'd191,8'd166} : s = 217;
	{8'd191,8'd167} : s = 214;
	{8'd191,8'd168} : s = 373;
	{8'd191,8'd169} : s = 89;
	{8'd191,8'd170} : s = 213;
	{8'd191,8'd171} : s = 211;
	{8'd191,8'd172} : s = 371;
	{8'd191,8'd173} : s = 206;
	{8'd191,8'd174} : s = 366;
	{8'd191,8'd175} : s = 365;
	{8'd191,8'd176} : s = 478;
	{8'd191,8'd177} : s = 86;
	{8'd191,8'd178} : s = 205;
	{8'd191,8'd179} : s = 203;
	{8'd191,8'd180} : s = 363;
	{8'd191,8'd181} : s = 199;
	{8'd191,8'd182} : s = 359;
	{8'd191,8'd183} : s = 350;
	{8'd191,8'd184} : s = 477;
	{8'd191,8'd185} : s = 188;
	{8'd191,8'd186} : s = 349;
	{8'd191,8'd187} : s = 347;
	{8'd191,8'd188} : s = 475;
	{8'd191,8'd189} : s = 343;
	{8'd191,8'd190} : s = 471;
	{8'd191,8'd191} : s = 463;
	{8'd191,8'd192} : s = 509;
	{8'd191,8'd193} : s = 3;
	{8'd191,8'd194} : s = 22;
	{8'd191,8'd195} : s = 21;
	{8'd191,8'd196} : s = 85;
	{8'd191,8'd197} : s = 19;
	{8'd191,8'd198} : s = 83;
	{8'd191,8'd199} : s = 78;
	{8'd191,8'd200} : s = 186;
	{8'd191,8'd201} : s = 14;
	{8'd191,8'd202} : s = 77;
	{8'd191,8'd203} : s = 75;
	{8'd191,8'd204} : s = 185;
	{8'd191,8'd205} : s = 71;
	{8'd191,8'd206} : s = 182;
	{8'd191,8'd207} : s = 181;
	{8'd191,8'd208} : s = 335;
	{8'd191,8'd209} : s = 13;
	{8'd191,8'd210} : s = 60;
	{8'd191,8'd211} : s = 58;
	{8'd191,8'd212} : s = 179;
	{8'd191,8'd213} : s = 57;
	{8'd191,8'd214} : s = 174;
	{8'd191,8'd215} : s = 173;
	{8'd191,8'd216} : s = 318;
	{8'd191,8'd217} : s = 54;
	{8'd191,8'd218} : s = 171;
	{8'd191,8'd219} : s = 167;
	{8'd191,8'd220} : s = 317;
	{8'd191,8'd221} : s = 158;
	{8'd191,8'd222} : s = 315;
	{8'd191,8'd223} : s = 311;
	{8'd191,8'd224} : s = 446;
	{8'd191,8'd225} : s = 11;
	{8'd191,8'd226} : s = 53;
	{8'd191,8'd227} : s = 51;
	{8'd191,8'd228} : s = 157;
	{8'd191,8'd229} : s = 46;
	{8'd191,8'd230} : s = 155;
	{8'd191,8'd231} : s = 151;
	{8'd191,8'd232} : s = 303;
	{8'd191,8'd233} : s = 45;
	{8'd191,8'd234} : s = 143;
	{8'd191,8'd235} : s = 124;
	{8'd191,8'd236} : s = 287;
	{8'd191,8'd237} : s = 122;
	{8'd191,8'd238} : s = 252;
	{8'd191,8'd239} : s = 250;
	{8'd191,8'd240} : s = 445;
	{8'd191,8'd241} : s = 43;
	{8'd191,8'd242} : s = 121;
	{8'd191,8'd243} : s = 118;
	{8'd191,8'd244} : s = 249;
	{8'd191,8'd245} : s = 117;
	{8'd191,8'd246} : s = 246;
	{8'd191,8'd247} : s = 245;
	{8'd191,8'd248} : s = 443;
	{8'd191,8'd249} : s = 115;
	{8'd191,8'd250} : s = 243;
	{8'd191,8'd251} : s = 238;
	{8'd191,8'd252} : s = 439;
	{8'd191,8'd253} : s = 237;
	{8'd191,8'd254} : s = 431;
	{8'd191,8'd255} : s = 415;
	{8'd192,8'd0} : s = 20;
	{8'd192,8'd1} : s = 104;
	{8'd192,8'd2} : s = 100;
	{8'd192,8'd3} : s = 263;
	{8'd192,8'd4} : s = 98;
	{8'd192,8'd5} : s = 240;
	{8'd192,8'd6} : s = 232;
	{8'd192,8'd7} : s = 372;
	{8'd192,8'd8} : s = 97;
	{8'd192,8'd9} : s = 228;
	{8'd192,8'd10} : s = 226;
	{8'd192,8'd11} : s = 370;
	{8'd192,8'd12} : s = 225;
	{8'd192,8'd13} : s = 369;
	{8'd192,8'd14} : s = 364;
	{8'd192,8'd15} : s = 470;
	{8'd192,8'd16} : s = 88;
	{8'd192,8'd17} : s = 216;
	{8'd192,8'd18} : s = 212;
	{8'd192,8'd19} : s = 362;
	{8'd192,8'd20} : s = 210;
	{8'd192,8'd21} : s = 361;
	{8'd192,8'd22} : s = 358;
	{8'd192,8'd23} : s = 469;
	{8'd192,8'd24} : s = 209;
	{8'd192,8'd25} : s = 357;
	{8'd192,8'd26} : s = 355;
	{8'd192,8'd27} : s = 467;
	{8'd192,8'd28} : s = 348;
	{8'd192,8'd29} : s = 462;
	{8'd192,8'd30} : s = 461;
	{8'd192,8'd31} : s = 505;
	{8'd192,8'd32} : s = 84;
	{8'd192,8'd33} : s = 204;
	{8'd192,8'd34} : s = 202;
	{8'd192,8'd35} : s = 346;
	{8'd192,8'd36} : s = 201;
	{8'd192,8'd37} : s = 345;
	{8'd192,8'd38} : s = 342;
	{8'd192,8'd39} : s = 459;
	{8'd192,8'd40} : s = 198;
	{8'd192,8'd41} : s = 341;
	{8'd192,8'd42} : s = 339;
	{8'd192,8'd43} : s = 455;
	{8'd192,8'd44} : s = 334;
	{8'd192,8'd45} : s = 444;
	{8'd192,8'd46} : s = 442;
	{8'd192,8'd47} : s = 502;
	{8'd192,8'd48} : s = 197;
	{8'd192,8'd49} : s = 333;
	{8'd192,8'd50} : s = 331;
	{8'd192,8'd51} : s = 441;
	{8'd192,8'd52} : s = 327;
	{8'd192,8'd53} : s = 438;
	{8'd192,8'd54} : s = 437;
	{8'd192,8'd55} : s = 501;
	{8'd192,8'd56} : s = 316;
	{8'd192,8'd57} : s = 435;
	{8'd192,8'd58} : s = 430;
	{8'd192,8'd59} : s = 499;
	{8'd192,8'd60} : s = 429;
	{8'd192,8'd61} : s = 494;
	{8'd192,8'd62} : s = 493;
	{8'd192,8'd63} : s = 510;
	{8'd192,8'd64} : s = 1;
	{8'd192,8'd65} : s = 18;
	{8'd192,8'd66} : s = 17;
	{8'd192,8'd67} : s = 82;
	{8'd192,8'd68} : s = 12;
	{8'd192,8'd69} : s = 81;
	{8'd192,8'd70} : s = 76;
	{8'd192,8'd71} : s = 195;
	{8'd192,8'd72} : s = 10;
	{8'd192,8'd73} : s = 74;
	{8'd192,8'd74} : s = 73;
	{8'd192,8'd75} : s = 184;
	{8'd192,8'd76} : s = 70;
	{8'd192,8'd77} : s = 180;
	{8'd192,8'd78} : s = 178;
	{8'd192,8'd79} : s = 314;
	{8'd192,8'd80} : s = 9;
	{8'd192,8'd81} : s = 69;
	{8'd192,8'd82} : s = 67;
	{8'd192,8'd83} : s = 177;
	{8'd192,8'd84} : s = 56;
	{8'd192,8'd85} : s = 172;
	{8'd192,8'd86} : s = 170;
	{8'd192,8'd87} : s = 313;
	{8'd192,8'd88} : s = 52;
	{8'd192,8'd89} : s = 169;
	{8'd192,8'd90} : s = 166;
	{8'd192,8'd91} : s = 310;
	{8'd192,8'd92} : s = 165;
	{8'd192,8'd93} : s = 309;
	{8'd192,8'd94} : s = 307;
	{8'd192,8'd95} : s = 427;
	{8'd192,8'd96} : s = 6;
	{8'd192,8'd97} : s = 50;
	{8'd192,8'd98} : s = 49;
	{8'd192,8'd99} : s = 163;
	{8'd192,8'd100} : s = 44;
	{8'd192,8'd101} : s = 156;
	{8'd192,8'd102} : s = 154;
	{8'd192,8'd103} : s = 302;
	{8'd192,8'd104} : s = 42;
	{8'd192,8'd105} : s = 153;
	{8'd192,8'd106} : s = 150;
	{8'd192,8'd107} : s = 301;
	{8'd192,8'd108} : s = 149;
	{8'd192,8'd109} : s = 299;
	{8'd192,8'd110} : s = 295;
	{8'd192,8'd111} : s = 423;
	{8'd192,8'd112} : s = 41;
	{8'd192,8'd113} : s = 147;
	{8'd192,8'd114} : s = 142;
	{8'd192,8'd115} : s = 286;
	{8'd192,8'd116} : s = 141;
	{8'd192,8'd117} : s = 285;
	{8'd192,8'd118} : s = 283;
	{8'd192,8'd119} : s = 414;
	{8'd192,8'd120} : s = 139;
	{8'd192,8'd121} : s = 279;
	{8'd192,8'd122} : s = 271;
	{8'd192,8'd123} : s = 413;
	{8'd192,8'd124} : s = 248;
	{8'd192,8'd125} : s = 411;
	{8'd192,8'd126} : s = 407;
	{8'd192,8'd127} : s = 491;
	{8'd192,8'd128} : s = 5;
	{8'd192,8'd129} : s = 38;
	{8'd192,8'd130} : s = 37;
	{8'd192,8'd131} : s = 135;
	{8'd192,8'd132} : s = 35;
	{8'd192,8'd133} : s = 120;
	{8'd192,8'd134} : s = 116;
	{8'd192,8'd135} : s = 244;
	{8'd192,8'd136} : s = 28;
	{8'd192,8'd137} : s = 114;
	{8'd192,8'd138} : s = 113;
	{8'd192,8'd139} : s = 242;
	{8'd192,8'd140} : s = 108;
	{8'd192,8'd141} : s = 241;
	{8'd192,8'd142} : s = 236;
	{8'd192,8'd143} : s = 399;
	{8'd192,8'd144} : s = 26;
	{8'd192,8'd145} : s = 106;
	{8'd192,8'd146} : s = 105;
	{8'd192,8'd147} : s = 234;
	{8'd192,8'd148} : s = 102;
	{8'd192,8'd149} : s = 233;
	{8'd192,8'd150} : s = 230;
	{8'd192,8'd151} : s = 380;
	{8'd192,8'd152} : s = 101;
	{8'd192,8'd153} : s = 229;
	{8'd192,8'd154} : s = 227;
	{8'd192,8'd155} : s = 378;
	{8'd192,8'd156} : s = 220;
	{8'd192,8'd157} : s = 377;
	{8'd192,8'd158} : s = 374;
	{8'd192,8'd159} : s = 487;
	{8'd192,8'd160} : s = 25;
	{8'd192,8'd161} : s = 99;
	{8'd192,8'd162} : s = 92;
	{8'd192,8'd163} : s = 218;
	{8'd192,8'd164} : s = 90;
	{8'd192,8'd165} : s = 217;
	{8'd192,8'd166} : s = 214;
	{8'd192,8'd167} : s = 373;
	{8'd192,8'd168} : s = 89;
	{8'd192,8'd169} : s = 213;
	{8'd192,8'd170} : s = 211;
	{8'd192,8'd171} : s = 371;
	{8'd192,8'd172} : s = 206;
	{8'd192,8'd173} : s = 366;
	{8'd192,8'd174} : s = 365;
	{8'd192,8'd175} : s = 478;
	{8'd192,8'd176} : s = 86;
	{8'd192,8'd177} : s = 205;
	{8'd192,8'd178} : s = 203;
	{8'd192,8'd179} : s = 363;
	{8'd192,8'd180} : s = 199;
	{8'd192,8'd181} : s = 359;
	{8'd192,8'd182} : s = 350;
	{8'd192,8'd183} : s = 477;
	{8'd192,8'd184} : s = 188;
	{8'd192,8'd185} : s = 349;
	{8'd192,8'd186} : s = 347;
	{8'd192,8'd187} : s = 475;
	{8'd192,8'd188} : s = 343;
	{8'd192,8'd189} : s = 471;
	{8'd192,8'd190} : s = 463;
	{8'd192,8'd191} : s = 509;
	{8'd192,8'd192} : s = 3;
	{8'd192,8'd193} : s = 22;
	{8'd192,8'd194} : s = 21;
	{8'd192,8'd195} : s = 85;
	{8'd192,8'd196} : s = 19;
	{8'd192,8'd197} : s = 83;
	{8'd192,8'd198} : s = 78;
	{8'd192,8'd199} : s = 186;
	{8'd192,8'd200} : s = 14;
	{8'd192,8'd201} : s = 77;
	{8'd192,8'd202} : s = 75;
	{8'd192,8'd203} : s = 185;
	{8'd192,8'd204} : s = 71;
	{8'd192,8'd205} : s = 182;
	{8'd192,8'd206} : s = 181;
	{8'd192,8'd207} : s = 335;
	{8'd192,8'd208} : s = 13;
	{8'd192,8'd209} : s = 60;
	{8'd192,8'd210} : s = 58;
	{8'd192,8'd211} : s = 179;
	{8'd192,8'd212} : s = 57;
	{8'd192,8'd213} : s = 174;
	{8'd192,8'd214} : s = 173;
	{8'd192,8'd215} : s = 318;
	{8'd192,8'd216} : s = 54;
	{8'd192,8'd217} : s = 171;
	{8'd192,8'd218} : s = 167;
	{8'd192,8'd219} : s = 317;
	{8'd192,8'd220} : s = 158;
	{8'd192,8'd221} : s = 315;
	{8'd192,8'd222} : s = 311;
	{8'd192,8'd223} : s = 446;
	{8'd192,8'd224} : s = 11;
	{8'd192,8'd225} : s = 53;
	{8'd192,8'd226} : s = 51;
	{8'd192,8'd227} : s = 157;
	{8'd192,8'd228} : s = 46;
	{8'd192,8'd229} : s = 155;
	{8'd192,8'd230} : s = 151;
	{8'd192,8'd231} : s = 303;
	{8'd192,8'd232} : s = 45;
	{8'd192,8'd233} : s = 143;
	{8'd192,8'd234} : s = 124;
	{8'd192,8'd235} : s = 287;
	{8'd192,8'd236} : s = 122;
	{8'd192,8'd237} : s = 252;
	{8'd192,8'd238} : s = 250;
	{8'd192,8'd239} : s = 445;
	{8'd192,8'd240} : s = 43;
	{8'd192,8'd241} : s = 121;
	{8'd192,8'd242} : s = 118;
	{8'd192,8'd243} : s = 249;
	{8'd192,8'd244} : s = 117;
	{8'd192,8'd245} : s = 246;
	{8'd192,8'd246} : s = 245;
	{8'd192,8'd247} : s = 443;
	{8'd192,8'd248} : s = 115;
	{8'd192,8'd249} : s = 243;
	{8'd192,8'd250} : s = 238;
	{8'd192,8'd251} : s = 439;
	{8'd192,8'd252} : s = 237;
	{8'd192,8'd253} : s = 431;
	{8'd192,8'd254} : s = 415;
	{8'd192,8'd255} : s = 507;
	{8'd193,8'd0} : s = 104;
	{8'd193,8'd1} : s = 100;
	{8'd193,8'd2} : s = 263;
	{8'd193,8'd3} : s = 98;
	{8'd193,8'd4} : s = 240;
	{8'd193,8'd5} : s = 232;
	{8'd193,8'd6} : s = 372;
	{8'd193,8'd7} : s = 97;
	{8'd193,8'd8} : s = 228;
	{8'd193,8'd9} : s = 226;
	{8'd193,8'd10} : s = 370;
	{8'd193,8'd11} : s = 225;
	{8'd193,8'd12} : s = 369;
	{8'd193,8'd13} : s = 364;
	{8'd193,8'd14} : s = 470;
	{8'd193,8'd15} : s = 88;
	{8'd193,8'd16} : s = 216;
	{8'd193,8'd17} : s = 212;
	{8'd193,8'd18} : s = 362;
	{8'd193,8'd19} : s = 210;
	{8'd193,8'd20} : s = 361;
	{8'd193,8'd21} : s = 358;
	{8'd193,8'd22} : s = 469;
	{8'd193,8'd23} : s = 209;
	{8'd193,8'd24} : s = 357;
	{8'd193,8'd25} : s = 355;
	{8'd193,8'd26} : s = 467;
	{8'd193,8'd27} : s = 348;
	{8'd193,8'd28} : s = 462;
	{8'd193,8'd29} : s = 461;
	{8'd193,8'd30} : s = 505;
	{8'd193,8'd31} : s = 84;
	{8'd193,8'd32} : s = 204;
	{8'd193,8'd33} : s = 202;
	{8'd193,8'd34} : s = 346;
	{8'd193,8'd35} : s = 201;
	{8'd193,8'd36} : s = 345;
	{8'd193,8'd37} : s = 342;
	{8'd193,8'd38} : s = 459;
	{8'd193,8'd39} : s = 198;
	{8'd193,8'd40} : s = 341;
	{8'd193,8'd41} : s = 339;
	{8'd193,8'd42} : s = 455;
	{8'd193,8'd43} : s = 334;
	{8'd193,8'd44} : s = 444;
	{8'd193,8'd45} : s = 442;
	{8'd193,8'd46} : s = 502;
	{8'd193,8'd47} : s = 197;
	{8'd193,8'd48} : s = 333;
	{8'd193,8'd49} : s = 331;
	{8'd193,8'd50} : s = 441;
	{8'd193,8'd51} : s = 327;
	{8'd193,8'd52} : s = 438;
	{8'd193,8'd53} : s = 437;
	{8'd193,8'd54} : s = 501;
	{8'd193,8'd55} : s = 316;
	{8'd193,8'd56} : s = 435;
	{8'd193,8'd57} : s = 430;
	{8'd193,8'd58} : s = 499;
	{8'd193,8'd59} : s = 429;
	{8'd193,8'd60} : s = 494;
	{8'd193,8'd61} : s = 493;
	{8'd193,8'd62} : s = 510;
	{8'd193,8'd63} : s = 1;
	{8'd193,8'd64} : s = 18;
	{8'd193,8'd65} : s = 17;
	{8'd193,8'd66} : s = 82;
	{8'd193,8'd67} : s = 12;
	{8'd193,8'd68} : s = 81;
	{8'd193,8'd69} : s = 76;
	{8'd193,8'd70} : s = 195;
	{8'd193,8'd71} : s = 10;
	{8'd193,8'd72} : s = 74;
	{8'd193,8'd73} : s = 73;
	{8'd193,8'd74} : s = 184;
	{8'd193,8'd75} : s = 70;
	{8'd193,8'd76} : s = 180;
	{8'd193,8'd77} : s = 178;
	{8'd193,8'd78} : s = 314;
	{8'd193,8'd79} : s = 9;
	{8'd193,8'd80} : s = 69;
	{8'd193,8'd81} : s = 67;
	{8'd193,8'd82} : s = 177;
	{8'd193,8'd83} : s = 56;
	{8'd193,8'd84} : s = 172;
	{8'd193,8'd85} : s = 170;
	{8'd193,8'd86} : s = 313;
	{8'd193,8'd87} : s = 52;
	{8'd193,8'd88} : s = 169;
	{8'd193,8'd89} : s = 166;
	{8'd193,8'd90} : s = 310;
	{8'd193,8'd91} : s = 165;
	{8'd193,8'd92} : s = 309;
	{8'd193,8'd93} : s = 307;
	{8'd193,8'd94} : s = 427;
	{8'd193,8'd95} : s = 6;
	{8'd193,8'd96} : s = 50;
	{8'd193,8'd97} : s = 49;
	{8'd193,8'd98} : s = 163;
	{8'd193,8'd99} : s = 44;
	{8'd193,8'd100} : s = 156;
	{8'd193,8'd101} : s = 154;
	{8'd193,8'd102} : s = 302;
	{8'd193,8'd103} : s = 42;
	{8'd193,8'd104} : s = 153;
	{8'd193,8'd105} : s = 150;
	{8'd193,8'd106} : s = 301;
	{8'd193,8'd107} : s = 149;
	{8'd193,8'd108} : s = 299;
	{8'd193,8'd109} : s = 295;
	{8'd193,8'd110} : s = 423;
	{8'd193,8'd111} : s = 41;
	{8'd193,8'd112} : s = 147;
	{8'd193,8'd113} : s = 142;
	{8'd193,8'd114} : s = 286;
	{8'd193,8'd115} : s = 141;
	{8'd193,8'd116} : s = 285;
	{8'd193,8'd117} : s = 283;
	{8'd193,8'd118} : s = 414;
	{8'd193,8'd119} : s = 139;
	{8'd193,8'd120} : s = 279;
	{8'd193,8'd121} : s = 271;
	{8'd193,8'd122} : s = 413;
	{8'd193,8'd123} : s = 248;
	{8'd193,8'd124} : s = 411;
	{8'd193,8'd125} : s = 407;
	{8'd193,8'd126} : s = 491;
	{8'd193,8'd127} : s = 5;
	{8'd193,8'd128} : s = 38;
	{8'd193,8'd129} : s = 37;
	{8'd193,8'd130} : s = 135;
	{8'd193,8'd131} : s = 35;
	{8'd193,8'd132} : s = 120;
	{8'd193,8'd133} : s = 116;
	{8'd193,8'd134} : s = 244;
	{8'd193,8'd135} : s = 28;
	{8'd193,8'd136} : s = 114;
	{8'd193,8'd137} : s = 113;
	{8'd193,8'd138} : s = 242;
	{8'd193,8'd139} : s = 108;
	{8'd193,8'd140} : s = 241;
	{8'd193,8'd141} : s = 236;
	{8'd193,8'd142} : s = 399;
	{8'd193,8'd143} : s = 26;
	{8'd193,8'd144} : s = 106;
	{8'd193,8'd145} : s = 105;
	{8'd193,8'd146} : s = 234;
	{8'd193,8'd147} : s = 102;
	{8'd193,8'd148} : s = 233;
	{8'd193,8'd149} : s = 230;
	{8'd193,8'd150} : s = 380;
	{8'd193,8'd151} : s = 101;
	{8'd193,8'd152} : s = 229;
	{8'd193,8'd153} : s = 227;
	{8'd193,8'd154} : s = 378;
	{8'd193,8'd155} : s = 220;
	{8'd193,8'd156} : s = 377;
	{8'd193,8'd157} : s = 374;
	{8'd193,8'd158} : s = 487;
	{8'd193,8'd159} : s = 25;
	{8'd193,8'd160} : s = 99;
	{8'd193,8'd161} : s = 92;
	{8'd193,8'd162} : s = 218;
	{8'd193,8'd163} : s = 90;
	{8'd193,8'd164} : s = 217;
	{8'd193,8'd165} : s = 214;
	{8'd193,8'd166} : s = 373;
	{8'd193,8'd167} : s = 89;
	{8'd193,8'd168} : s = 213;
	{8'd193,8'd169} : s = 211;
	{8'd193,8'd170} : s = 371;
	{8'd193,8'd171} : s = 206;
	{8'd193,8'd172} : s = 366;
	{8'd193,8'd173} : s = 365;
	{8'd193,8'd174} : s = 478;
	{8'd193,8'd175} : s = 86;
	{8'd193,8'd176} : s = 205;
	{8'd193,8'd177} : s = 203;
	{8'd193,8'd178} : s = 363;
	{8'd193,8'd179} : s = 199;
	{8'd193,8'd180} : s = 359;
	{8'd193,8'd181} : s = 350;
	{8'd193,8'd182} : s = 477;
	{8'd193,8'd183} : s = 188;
	{8'd193,8'd184} : s = 349;
	{8'd193,8'd185} : s = 347;
	{8'd193,8'd186} : s = 475;
	{8'd193,8'd187} : s = 343;
	{8'd193,8'd188} : s = 471;
	{8'd193,8'd189} : s = 463;
	{8'd193,8'd190} : s = 509;
	{8'd193,8'd191} : s = 3;
	{8'd193,8'd192} : s = 22;
	{8'd193,8'd193} : s = 21;
	{8'd193,8'd194} : s = 85;
	{8'd193,8'd195} : s = 19;
	{8'd193,8'd196} : s = 83;
	{8'd193,8'd197} : s = 78;
	{8'd193,8'd198} : s = 186;
	{8'd193,8'd199} : s = 14;
	{8'd193,8'd200} : s = 77;
	{8'd193,8'd201} : s = 75;
	{8'd193,8'd202} : s = 185;
	{8'd193,8'd203} : s = 71;
	{8'd193,8'd204} : s = 182;
	{8'd193,8'd205} : s = 181;
	{8'd193,8'd206} : s = 335;
	{8'd193,8'd207} : s = 13;
	{8'd193,8'd208} : s = 60;
	{8'd193,8'd209} : s = 58;
	{8'd193,8'd210} : s = 179;
	{8'd193,8'd211} : s = 57;
	{8'd193,8'd212} : s = 174;
	{8'd193,8'd213} : s = 173;
	{8'd193,8'd214} : s = 318;
	{8'd193,8'd215} : s = 54;
	{8'd193,8'd216} : s = 171;
	{8'd193,8'd217} : s = 167;
	{8'd193,8'd218} : s = 317;
	{8'd193,8'd219} : s = 158;
	{8'd193,8'd220} : s = 315;
	{8'd193,8'd221} : s = 311;
	{8'd193,8'd222} : s = 446;
	{8'd193,8'd223} : s = 11;
	{8'd193,8'd224} : s = 53;
	{8'd193,8'd225} : s = 51;
	{8'd193,8'd226} : s = 157;
	{8'd193,8'd227} : s = 46;
	{8'd193,8'd228} : s = 155;
	{8'd193,8'd229} : s = 151;
	{8'd193,8'd230} : s = 303;
	{8'd193,8'd231} : s = 45;
	{8'd193,8'd232} : s = 143;
	{8'd193,8'd233} : s = 124;
	{8'd193,8'd234} : s = 287;
	{8'd193,8'd235} : s = 122;
	{8'd193,8'd236} : s = 252;
	{8'd193,8'd237} : s = 250;
	{8'd193,8'd238} : s = 445;
	{8'd193,8'd239} : s = 43;
	{8'd193,8'd240} : s = 121;
	{8'd193,8'd241} : s = 118;
	{8'd193,8'd242} : s = 249;
	{8'd193,8'd243} : s = 117;
	{8'd193,8'd244} : s = 246;
	{8'd193,8'd245} : s = 245;
	{8'd193,8'd246} : s = 443;
	{8'd193,8'd247} : s = 115;
	{8'd193,8'd248} : s = 243;
	{8'd193,8'd249} : s = 238;
	{8'd193,8'd250} : s = 439;
	{8'd193,8'd251} : s = 237;
	{8'd193,8'd252} : s = 431;
	{8'd193,8'd253} : s = 415;
	{8'd193,8'd254} : s = 507;
	{8'd193,8'd255} : s = 7;
	{8'd194,8'd0} : s = 100;
	{8'd194,8'd1} : s = 263;
	{8'd194,8'd2} : s = 98;
	{8'd194,8'd3} : s = 240;
	{8'd194,8'd4} : s = 232;
	{8'd194,8'd5} : s = 372;
	{8'd194,8'd6} : s = 97;
	{8'd194,8'd7} : s = 228;
	{8'd194,8'd8} : s = 226;
	{8'd194,8'd9} : s = 370;
	{8'd194,8'd10} : s = 225;
	{8'd194,8'd11} : s = 369;
	{8'd194,8'd12} : s = 364;
	{8'd194,8'd13} : s = 470;
	{8'd194,8'd14} : s = 88;
	{8'd194,8'd15} : s = 216;
	{8'd194,8'd16} : s = 212;
	{8'd194,8'd17} : s = 362;
	{8'd194,8'd18} : s = 210;
	{8'd194,8'd19} : s = 361;
	{8'd194,8'd20} : s = 358;
	{8'd194,8'd21} : s = 469;
	{8'd194,8'd22} : s = 209;
	{8'd194,8'd23} : s = 357;
	{8'd194,8'd24} : s = 355;
	{8'd194,8'd25} : s = 467;
	{8'd194,8'd26} : s = 348;
	{8'd194,8'd27} : s = 462;
	{8'd194,8'd28} : s = 461;
	{8'd194,8'd29} : s = 505;
	{8'd194,8'd30} : s = 84;
	{8'd194,8'd31} : s = 204;
	{8'd194,8'd32} : s = 202;
	{8'd194,8'd33} : s = 346;
	{8'd194,8'd34} : s = 201;
	{8'd194,8'd35} : s = 345;
	{8'd194,8'd36} : s = 342;
	{8'd194,8'd37} : s = 459;
	{8'd194,8'd38} : s = 198;
	{8'd194,8'd39} : s = 341;
	{8'd194,8'd40} : s = 339;
	{8'd194,8'd41} : s = 455;
	{8'd194,8'd42} : s = 334;
	{8'd194,8'd43} : s = 444;
	{8'd194,8'd44} : s = 442;
	{8'd194,8'd45} : s = 502;
	{8'd194,8'd46} : s = 197;
	{8'd194,8'd47} : s = 333;
	{8'd194,8'd48} : s = 331;
	{8'd194,8'd49} : s = 441;
	{8'd194,8'd50} : s = 327;
	{8'd194,8'd51} : s = 438;
	{8'd194,8'd52} : s = 437;
	{8'd194,8'd53} : s = 501;
	{8'd194,8'd54} : s = 316;
	{8'd194,8'd55} : s = 435;
	{8'd194,8'd56} : s = 430;
	{8'd194,8'd57} : s = 499;
	{8'd194,8'd58} : s = 429;
	{8'd194,8'd59} : s = 494;
	{8'd194,8'd60} : s = 493;
	{8'd194,8'd61} : s = 510;
	{8'd194,8'd62} : s = 1;
	{8'd194,8'd63} : s = 18;
	{8'd194,8'd64} : s = 17;
	{8'd194,8'd65} : s = 82;
	{8'd194,8'd66} : s = 12;
	{8'd194,8'd67} : s = 81;
	{8'd194,8'd68} : s = 76;
	{8'd194,8'd69} : s = 195;
	{8'd194,8'd70} : s = 10;
	{8'd194,8'd71} : s = 74;
	{8'd194,8'd72} : s = 73;
	{8'd194,8'd73} : s = 184;
	{8'd194,8'd74} : s = 70;
	{8'd194,8'd75} : s = 180;
	{8'd194,8'd76} : s = 178;
	{8'd194,8'd77} : s = 314;
	{8'd194,8'd78} : s = 9;
	{8'd194,8'd79} : s = 69;
	{8'd194,8'd80} : s = 67;
	{8'd194,8'd81} : s = 177;
	{8'd194,8'd82} : s = 56;
	{8'd194,8'd83} : s = 172;
	{8'd194,8'd84} : s = 170;
	{8'd194,8'd85} : s = 313;
	{8'd194,8'd86} : s = 52;
	{8'd194,8'd87} : s = 169;
	{8'd194,8'd88} : s = 166;
	{8'd194,8'd89} : s = 310;
	{8'd194,8'd90} : s = 165;
	{8'd194,8'd91} : s = 309;
	{8'd194,8'd92} : s = 307;
	{8'd194,8'd93} : s = 427;
	{8'd194,8'd94} : s = 6;
	{8'd194,8'd95} : s = 50;
	{8'd194,8'd96} : s = 49;
	{8'd194,8'd97} : s = 163;
	{8'd194,8'd98} : s = 44;
	{8'd194,8'd99} : s = 156;
	{8'd194,8'd100} : s = 154;
	{8'd194,8'd101} : s = 302;
	{8'd194,8'd102} : s = 42;
	{8'd194,8'd103} : s = 153;
	{8'd194,8'd104} : s = 150;
	{8'd194,8'd105} : s = 301;
	{8'd194,8'd106} : s = 149;
	{8'd194,8'd107} : s = 299;
	{8'd194,8'd108} : s = 295;
	{8'd194,8'd109} : s = 423;
	{8'd194,8'd110} : s = 41;
	{8'd194,8'd111} : s = 147;
	{8'd194,8'd112} : s = 142;
	{8'd194,8'd113} : s = 286;
	{8'd194,8'd114} : s = 141;
	{8'd194,8'd115} : s = 285;
	{8'd194,8'd116} : s = 283;
	{8'd194,8'd117} : s = 414;
	{8'd194,8'd118} : s = 139;
	{8'd194,8'd119} : s = 279;
	{8'd194,8'd120} : s = 271;
	{8'd194,8'd121} : s = 413;
	{8'd194,8'd122} : s = 248;
	{8'd194,8'd123} : s = 411;
	{8'd194,8'd124} : s = 407;
	{8'd194,8'd125} : s = 491;
	{8'd194,8'd126} : s = 5;
	{8'd194,8'd127} : s = 38;
	{8'd194,8'd128} : s = 37;
	{8'd194,8'd129} : s = 135;
	{8'd194,8'd130} : s = 35;
	{8'd194,8'd131} : s = 120;
	{8'd194,8'd132} : s = 116;
	{8'd194,8'd133} : s = 244;
	{8'd194,8'd134} : s = 28;
	{8'd194,8'd135} : s = 114;
	{8'd194,8'd136} : s = 113;
	{8'd194,8'd137} : s = 242;
	{8'd194,8'd138} : s = 108;
	{8'd194,8'd139} : s = 241;
	{8'd194,8'd140} : s = 236;
	{8'd194,8'd141} : s = 399;
	{8'd194,8'd142} : s = 26;
	{8'd194,8'd143} : s = 106;
	{8'd194,8'd144} : s = 105;
	{8'd194,8'd145} : s = 234;
	{8'd194,8'd146} : s = 102;
	{8'd194,8'd147} : s = 233;
	{8'd194,8'd148} : s = 230;
	{8'd194,8'd149} : s = 380;
	{8'd194,8'd150} : s = 101;
	{8'd194,8'd151} : s = 229;
	{8'd194,8'd152} : s = 227;
	{8'd194,8'd153} : s = 378;
	{8'd194,8'd154} : s = 220;
	{8'd194,8'd155} : s = 377;
	{8'd194,8'd156} : s = 374;
	{8'd194,8'd157} : s = 487;
	{8'd194,8'd158} : s = 25;
	{8'd194,8'd159} : s = 99;
	{8'd194,8'd160} : s = 92;
	{8'd194,8'd161} : s = 218;
	{8'd194,8'd162} : s = 90;
	{8'd194,8'd163} : s = 217;
	{8'd194,8'd164} : s = 214;
	{8'd194,8'd165} : s = 373;
	{8'd194,8'd166} : s = 89;
	{8'd194,8'd167} : s = 213;
	{8'd194,8'd168} : s = 211;
	{8'd194,8'd169} : s = 371;
	{8'd194,8'd170} : s = 206;
	{8'd194,8'd171} : s = 366;
	{8'd194,8'd172} : s = 365;
	{8'd194,8'd173} : s = 478;
	{8'd194,8'd174} : s = 86;
	{8'd194,8'd175} : s = 205;
	{8'd194,8'd176} : s = 203;
	{8'd194,8'd177} : s = 363;
	{8'd194,8'd178} : s = 199;
	{8'd194,8'd179} : s = 359;
	{8'd194,8'd180} : s = 350;
	{8'd194,8'd181} : s = 477;
	{8'd194,8'd182} : s = 188;
	{8'd194,8'd183} : s = 349;
	{8'd194,8'd184} : s = 347;
	{8'd194,8'd185} : s = 475;
	{8'd194,8'd186} : s = 343;
	{8'd194,8'd187} : s = 471;
	{8'd194,8'd188} : s = 463;
	{8'd194,8'd189} : s = 509;
	{8'd194,8'd190} : s = 3;
	{8'd194,8'd191} : s = 22;
	{8'd194,8'd192} : s = 21;
	{8'd194,8'd193} : s = 85;
	{8'd194,8'd194} : s = 19;
	{8'd194,8'd195} : s = 83;
	{8'd194,8'd196} : s = 78;
	{8'd194,8'd197} : s = 186;
	{8'd194,8'd198} : s = 14;
	{8'd194,8'd199} : s = 77;
	{8'd194,8'd200} : s = 75;
	{8'd194,8'd201} : s = 185;
	{8'd194,8'd202} : s = 71;
	{8'd194,8'd203} : s = 182;
	{8'd194,8'd204} : s = 181;
	{8'd194,8'd205} : s = 335;
	{8'd194,8'd206} : s = 13;
	{8'd194,8'd207} : s = 60;
	{8'd194,8'd208} : s = 58;
	{8'd194,8'd209} : s = 179;
	{8'd194,8'd210} : s = 57;
	{8'd194,8'd211} : s = 174;
	{8'd194,8'd212} : s = 173;
	{8'd194,8'd213} : s = 318;
	{8'd194,8'd214} : s = 54;
	{8'd194,8'd215} : s = 171;
	{8'd194,8'd216} : s = 167;
	{8'd194,8'd217} : s = 317;
	{8'd194,8'd218} : s = 158;
	{8'd194,8'd219} : s = 315;
	{8'd194,8'd220} : s = 311;
	{8'd194,8'd221} : s = 446;
	{8'd194,8'd222} : s = 11;
	{8'd194,8'd223} : s = 53;
	{8'd194,8'd224} : s = 51;
	{8'd194,8'd225} : s = 157;
	{8'd194,8'd226} : s = 46;
	{8'd194,8'd227} : s = 155;
	{8'd194,8'd228} : s = 151;
	{8'd194,8'd229} : s = 303;
	{8'd194,8'd230} : s = 45;
	{8'd194,8'd231} : s = 143;
	{8'd194,8'd232} : s = 124;
	{8'd194,8'd233} : s = 287;
	{8'd194,8'd234} : s = 122;
	{8'd194,8'd235} : s = 252;
	{8'd194,8'd236} : s = 250;
	{8'd194,8'd237} : s = 445;
	{8'd194,8'd238} : s = 43;
	{8'd194,8'd239} : s = 121;
	{8'd194,8'd240} : s = 118;
	{8'd194,8'd241} : s = 249;
	{8'd194,8'd242} : s = 117;
	{8'd194,8'd243} : s = 246;
	{8'd194,8'd244} : s = 245;
	{8'd194,8'd245} : s = 443;
	{8'd194,8'd246} : s = 115;
	{8'd194,8'd247} : s = 243;
	{8'd194,8'd248} : s = 238;
	{8'd194,8'd249} : s = 439;
	{8'd194,8'd250} : s = 237;
	{8'd194,8'd251} : s = 431;
	{8'd194,8'd252} : s = 415;
	{8'd194,8'd253} : s = 507;
	{8'd194,8'd254} : s = 7;
	{8'd194,8'd255} : s = 39;
	{8'd195,8'd0} : s = 263;
	{8'd195,8'd1} : s = 98;
	{8'd195,8'd2} : s = 240;
	{8'd195,8'd3} : s = 232;
	{8'd195,8'd4} : s = 372;
	{8'd195,8'd5} : s = 97;
	{8'd195,8'd6} : s = 228;
	{8'd195,8'd7} : s = 226;
	{8'd195,8'd8} : s = 370;
	{8'd195,8'd9} : s = 225;
	{8'd195,8'd10} : s = 369;
	{8'd195,8'd11} : s = 364;
	{8'd195,8'd12} : s = 470;
	{8'd195,8'd13} : s = 88;
	{8'd195,8'd14} : s = 216;
	{8'd195,8'd15} : s = 212;
	{8'd195,8'd16} : s = 362;
	{8'd195,8'd17} : s = 210;
	{8'd195,8'd18} : s = 361;
	{8'd195,8'd19} : s = 358;
	{8'd195,8'd20} : s = 469;
	{8'd195,8'd21} : s = 209;
	{8'd195,8'd22} : s = 357;
	{8'd195,8'd23} : s = 355;
	{8'd195,8'd24} : s = 467;
	{8'd195,8'd25} : s = 348;
	{8'd195,8'd26} : s = 462;
	{8'd195,8'd27} : s = 461;
	{8'd195,8'd28} : s = 505;
	{8'd195,8'd29} : s = 84;
	{8'd195,8'd30} : s = 204;
	{8'd195,8'd31} : s = 202;
	{8'd195,8'd32} : s = 346;
	{8'd195,8'd33} : s = 201;
	{8'd195,8'd34} : s = 345;
	{8'd195,8'd35} : s = 342;
	{8'd195,8'd36} : s = 459;
	{8'd195,8'd37} : s = 198;
	{8'd195,8'd38} : s = 341;
	{8'd195,8'd39} : s = 339;
	{8'd195,8'd40} : s = 455;
	{8'd195,8'd41} : s = 334;
	{8'd195,8'd42} : s = 444;
	{8'd195,8'd43} : s = 442;
	{8'd195,8'd44} : s = 502;
	{8'd195,8'd45} : s = 197;
	{8'd195,8'd46} : s = 333;
	{8'd195,8'd47} : s = 331;
	{8'd195,8'd48} : s = 441;
	{8'd195,8'd49} : s = 327;
	{8'd195,8'd50} : s = 438;
	{8'd195,8'd51} : s = 437;
	{8'd195,8'd52} : s = 501;
	{8'd195,8'd53} : s = 316;
	{8'd195,8'd54} : s = 435;
	{8'd195,8'd55} : s = 430;
	{8'd195,8'd56} : s = 499;
	{8'd195,8'd57} : s = 429;
	{8'd195,8'd58} : s = 494;
	{8'd195,8'd59} : s = 493;
	{8'd195,8'd60} : s = 510;
	{8'd195,8'd61} : s = 1;
	{8'd195,8'd62} : s = 18;
	{8'd195,8'd63} : s = 17;
	{8'd195,8'd64} : s = 82;
	{8'd195,8'd65} : s = 12;
	{8'd195,8'd66} : s = 81;
	{8'd195,8'd67} : s = 76;
	{8'd195,8'd68} : s = 195;
	{8'd195,8'd69} : s = 10;
	{8'd195,8'd70} : s = 74;
	{8'd195,8'd71} : s = 73;
	{8'd195,8'd72} : s = 184;
	{8'd195,8'd73} : s = 70;
	{8'd195,8'd74} : s = 180;
	{8'd195,8'd75} : s = 178;
	{8'd195,8'd76} : s = 314;
	{8'd195,8'd77} : s = 9;
	{8'd195,8'd78} : s = 69;
	{8'd195,8'd79} : s = 67;
	{8'd195,8'd80} : s = 177;
	{8'd195,8'd81} : s = 56;
	{8'd195,8'd82} : s = 172;
	{8'd195,8'd83} : s = 170;
	{8'd195,8'd84} : s = 313;
	{8'd195,8'd85} : s = 52;
	{8'd195,8'd86} : s = 169;
	{8'd195,8'd87} : s = 166;
	{8'd195,8'd88} : s = 310;
	{8'd195,8'd89} : s = 165;
	{8'd195,8'd90} : s = 309;
	{8'd195,8'd91} : s = 307;
	{8'd195,8'd92} : s = 427;
	{8'd195,8'd93} : s = 6;
	{8'd195,8'd94} : s = 50;
	{8'd195,8'd95} : s = 49;
	{8'd195,8'd96} : s = 163;
	{8'd195,8'd97} : s = 44;
	{8'd195,8'd98} : s = 156;
	{8'd195,8'd99} : s = 154;
	{8'd195,8'd100} : s = 302;
	{8'd195,8'd101} : s = 42;
	{8'd195,8'd102} : s = 153;
	{8'd195,8'd103} : s = 150;
	{8'd195,8'd104} : s = 301;
	{8'd195,8'd105} : s = 149;
	{8'd195,8'd106} : s = 299;
	{8'd195,8'd107} : s = 295;
	{8'd195,8'd108} : s = 423;
	{8'd195,8'd109} : s = 41;
	{8'd195,8'd110} : s = 147;
	{8'd195,8'd111} : s = 142;
	{8'd195,8'd112} : s = 286;
	{8'd195,8'd113} : s = 141;
	{8'd195,8'd114} : s = 285;
	{8'd195,8'd115} : s = 283;
	{8'd195,8'd116} : s = 414;
	{8'd195,8'd117} : s = 139;
	{8'd195,8'd118} : s = 279;
	{8'd195,8'd119} : s = 271;
	{8'd195,8'd120} : s = 413;
	{8'd195,8'd121} : s = 248;
	{8'd195,8'd122} : s = 411;
	{8'd195,8'd123} : s = 407;
	{8'd195,8'd124} : s = 491;
	{8'd195,8'd125} : s = 5;
	{8'd195,8'd126} : s = 38;
	{8'd195,8'd127} : s = 37;
	{8'd195,8'd128} : s = 135;
	{8'd195,8'd129} : s = 35;
	{8'd195,8'd130} : s = 120;
	{8'd195,8'd131} : s = 116;
	{8'd195,8'd132} : s = 244;
	{8'd195,8'd133} : s = 28;
	{8'd195,8'd134} : s = 114;
	{8'd195,8'd135} : s = 113;
	{8'd195,8'd136} : s = 242;
	{8'd195,8'd137} : s = 108;
	{8'd195,8'd138} : s = 241;
	{8'd195,8'd139} : s = 236;
	{8'd195,8'd140} : s = 399;
	{8'd195,8'd141} : s = 26;
	{8'd195,8'd142} : s = 106;
	{8'd195,8'd143} : s = 105;
	{8'd195,8'd144} : s = 234;
	{8'd195,8'd145} : s = 102;
	{8'd195,8'd146} : s = 233;
	{8'd195,8'd147} : s = 230;
	{8'd195,8'd148} : s = 380;
	{8'd195,8'd149} : s = 101;
	{8'd195,8'd150} : s = 229;
	{8'd195,8'd151} : s = 227;
	{8'd195,8'd152} : s = 378;
	{8'd195,8'd153} : s = 220;
	{8'd195,8'd154} : s = 377;
	{8'd195,8'd155} : s = 374;
	{8'd195,8'd156} : s = 487;
	{8'd195,8'd157} : s = 25;
	{8'd195,8'd158} : s = 99;
	{8'd195,8'd159} : s = 92;
	{8'd195,8'd160} : s = 218;
	{8'd195,8'd161} : s = 90;
	{8'd195,8'd162} : s = 217;
	{8'd195,8'd163} : s = 214;
	{8'd195,8'd164} : s = 373;
	{8'd195,8'd165} : s = 89;
	{8'd195,8'd166} : s = 213;
	{8'd195,8'd167} : s = 211;
	{8'd195,8'd168} : s = 371;
	{8'd195,8'd169} : s = 206;
	{8'd195,8'd170} : s = 366;
	{8'd195,8'd171} : s = 365;
	{8'd195,8'd172} : s = 478;
	{8'd195,8'd173} : s = 86;
	{8'd195,8'd174} : s = 205;
	{8'd195,8'd175} : s = 203;
	{8'd195,8'd176} : s = 363;
	{8'd195,8'd177} : s = 199;
	{8'd195,8'd178} : s = 359;
	{8'd195,8'd179} : s = 350;
	{8'd195,8'd180} : s = 477;
	{8'd195,8'd181} : s = 188;
	{8'd195,8'd182} : s = 349;
	{8'd195,8'd183} : s = 347;
	{8'd195,8'd184} : s = 475;
	{8'd195,8'd185} : s = 343;
	{8'd195,8'd186} : s = 471;
	{8'd195,8'd187} : s = 463;
	{8'd195,8'd188} : s = 509;
	{8'd195,8'd189} : s = 3;
	{8'd195,8'd190} : s = 22;
	{8'd195,8'd191} : s = 21;
	{8'd195,8'd192} : s = 85;
	{8'd195,8'd193} : s = 19;
	{8'd195,8'd194} : s = 83;
	{8'd195,8'd195} : s = 78;
	{8'd195,8'd196} : s = 186;
	{8'd195,8'd197} : s = 14;
	{8'd195,8'd198} : s = 77;
	{8'd195,8'd199} : s = 75;
	{8'd195,8'd200} : s = 185;
	{8'd195,8'd201} : s = 71;
	{8'd195,8'd202} : s = 182;
	{8'd195,8'd203} : s = 181;
	{8'd195,8'd204} : s = 335;
	{8'd195,8'd205} : s = 13;
	{8'd195,8'd206} : s = 60;
	{8'd195,8'd207} : s = 58;
	{8'd195,8'd208} : s = 179;
	{8'd195,8'd209} : s = 57;
	{8'd195,8'd210} : s = 174;
	{8'd195,8'd211} : s = 173;
	{8'd195,8'd212} : s = 318;
	{8'd195,8'd213} : s = 54;
	{8'd195,8'd214} : s = 171;
	{8'd195,8'd215} : s = 167;
	{8'd195,8'd216} : s = 317;
	{8'd195,8'd217} : s = 158;
	{8'd195,8'd218} : s = 315;
	{8'd195,8'd219} : s = 311;
	{8'd195,8'd220} : s = 446;
	{8'd195,8'd221} : s = 11;
	{8'd195,8'd222} : s = 53;
	{8'd195,8'd223} : s = 51;
	{8'd195,8'd224} : s = 157;
	{8'd195,8'd225} : s = 46;
	{8'd195,8'd226} : s = 155;
	{8'd195,8'd227} : s = 151;
	{8'd195,8'd228} : s = 303;
	{8'd195,8'd229} : s = 45;
	{8'd195,8'd230} : s = 143;
	{8'd195,8'd231} : s = 124;
	{8'd195,8'd232} : s = 287;
	{8'd195,8'd233} : s = 122;
	{8'd195,8'd234} : s = 252;
	{8'd195,8'd235} : s = 250;
	{8'd195,8'd236} : s = 445;
	{8'd195,8'd237} : s = 43;
	{8'd195,8'd238} : s = 121;
	{8'd195,8'd239} : s = 118;
	{8'd195,8'd240} : s = 249;
	{8'd195,8'd241} : s = 117;
	{8'd195,8'd242} : s = 246;
	{8'd195,8'd243} : s = 245;
	{8'd195,8'd244} : s = 443;
	{8'd195,8'd245} : s = 115;
	{8'd195,8'd246} : s = 243;
	{8'd195,8'd247} : s = 238;
	{8'd195,8'd248} : s = 439;
	{8'd195,8'd249} : s = 237;
	{8'd195,8'd250} : s = 431;
	{8'd195,8'd251} : s = 415;
	{8'd195,8'd252} : s = 507;
	{8'd195,8'd253} : s = 7;
	{8'd195,8'd254} : s = 39;
	{8'd195,8'd255} : s = 30;
	{8'd196,8'd0} : s = 98;
	{8'd196,8'd1} : s = 240;
	{8'd196,8'd2} : s = 232;
	{8'd196,8'd3} : s = 372;
	{8'd196,8'd4} : s = 97;
	{8'd196,8'd5} : s = 228;
	{8'd196,8'd6} : s = 226;
	{8'd196,8'd7} : s = 370;
	{8'd196,8'd8} : s = 225;
	{8'd196,8'd9} : s = 369;
	{8'd196,8'd10} : s = 364;
	{8'd196,8'd11} : s = 470;
	{8'd196,8'd12} : s = 88;
	{8'd196,8'd13} : s = 216;
	{8'd196,8'd14} : s = 212;
	{8'd196,8'd15} : s = 362;
	{8'd196,8'd16} : s = 210;
	{8'd196,8'd17} : s = 361;
	{8'd196,8'd18} : s = 358;
	{8'd196,8'd19} : s = 469;
	{8'd196,8'd20} : s = 209;
	{8'd196,8'd21} : s = 357;
	{8'd196,8'd22} : s = 355;
	{8'd196,8'd23} : s = 467;
	{8'd196,8'd24} : s = 348;
	{8'd196,8'd25} : s = 462;
	{8'd196,8'd26} : s = 461;
	{8'd196,8'd27} : s = 505;
	{8'd196,8'd28} : s = 84;
	{8'd196,8'd29} : s = 204;
	{8'd196,8'd30} : s = 202;
	{8'd196,8'd31} : s = 346;
	{8'd196,8'd32} : s = 201;
	{8'd196,8'd33} : s = 345;
	{8'd196,8'd34} : s = 342;
	{8'd196,8'd35} : s = 459;
	{8'd196,8'd36} : s = 198;
	{8'd196,8'd37} : s = 341;
	{8'd196,8'd38} : s = 339;
	{8'd196,8'd39} : s = 455;
	{8'd196,8'd40} : s = 334;
	{8'd196,8'd41} : s = 444;
	{8'd196,8'd42} : s = 442;
	{8'd196,8'd43} : s = 502;
	{8'd196,8'd44} : s = 197;
	{8'd196,8'd45} : s = 333;
	{8'd196,8'd46} : s = 331;
	{8'd196,8'd47} : s = 441;
	{8'd196,8'd48} : s = 327;
	{8'd196,8'd49} : s = 438;
	{8'd196,8'd50} : s = 437;
	{8'd196,8'd51} : s = 501;
	{8'd196,8'd52} : s = 316;
	{8'd196,8'd53} : s = 435;
	{8'd196,8'd54} : s = 430;
	{8'd196,8'd55} : s = 499;
	{8'd196,8'd56} : s = 429;
	{8'd196,8'd57} : s = 494;
	{8'd196,8'd58} : s = 493;
	{8'd196,8'd59} : s = 510;
	{8'd196,8'd60} : s = 1;
	{8'd196,8'd61} : s = 18;
	{8'd196,8'd62} : s = 17;
	{8'd196,8'd63} : s = 82;
	{8'd196,8'd64} : s = 12;
	{8'd196,8'd65} : s = 81;
	{8'd196,8'd66} : s = 76;
	{8'd196,8'd67} : s = 195;
	{8'd196,8'd68} : s = 10;
	{8'd196,8'd69} : s = 74;
	{8'd196,8'd70} : s = 73;
	{8'd196,8'd71} : s = 184;
	{8'd196,8'd72} : s = 70;
	{8'd196,8'd73} : s = 180;
	{8'd196,8'd74} : s = 178;
	{8'd196,8'd75} : s = 314;
	{8'd196,8'd76} : s = 9;
	{8'd196,8'd77} : s = 69;
	{8'd196,8'd78} : s = 67;
	{8'd196,8'd79} : s = 177;
	{8'd196,8'd80} : s = 56;
	{8'd196,8'd81} : s = 172;
	{8'd196,8'd82} : s = 170;
	{8'd196,8'd83} : s = 313;
	{8'd196,8'd84} : s = 52;
	{8'd196,8'd85} : s = 169;
	{8'd196,8'd86} : s = 166;
	{8'd196,8'd87} : s = 310;
	{8'd196,8'd88} : s = 165;
	{8'd196,8'd89} : s = 309;
	{8'd196,8'd90} : s = 307;
	{8'd196,8'd91} : s = 427;
	{8'd196,8'd92} : s = 6;
	{8'd196,8'd93} : s = 50;
	{8'd196,8'd94} : s = 49;
	{8'd196,8'd95} : s = 163;
	{8'd196,8'd96} : s = 44;
	{8'd196,8'd97} : s = 156;
	{8'd196,8'd98} : s = 154;
	{8'd196,8'd99} : s = 302;
	{8'd196,8'd100} : s = 42;
	{8'd196,8'd101} : s = 153;
	{8'd196,8'd102} : s = 150;
	{8'd196,8'd103} : s = 301;
	{8'd196,8'd104} : s = 149;
	{8'd196,8'd105} : s = 299;
	{8'd196,8'd106} : s = 295;
	{8'd196,8'd107} : s = 423;
	{8'd196,8'd108} : s = 41;
	{8'd196,8'd109} : s = 147;
	{8'd196,8'd110} : s = 142;
	{8'd196,8'd111} : s = 286;
	{8'd196,8'd112} : s = 141;
	{8'd196,8'd113} : s = 285;
	{8'd196,8'd114} : s = 283;
	{8'd196,8'd115} : s = 414;
	{8'd196,8'd116} : s = 139;
	{8'd196,8'd117} : s = 279;
	{8'd196,8'd118} : s = 271;
	{8'd196,8'd119} : s = 413;
	{8'd196,8'd120} : s = 248;
	{8'd196,8'd121} : s = 411;
	{8'd196,8'd122} : s = 407;
	{8'd196,8'd123} : s = 491;
	{8'd196,8'd124} : s = 5;
	{8'd196,8'd125} : s = 38;
	{8'd196,8'd126} : s = 37;
	{8'd196,8'd127} : s = 135;
	{8'd196,8'd128} : s = 35;
	{8'd196,8'd129} : s = 120;
	{8'd196,8'd130} : s = 116;
	{8'd196,8'd131} : s = 244;
	{8'd196,8'd132} : s = 28;
	{8'd196,8'd133} : s = 114;
	{8'd196,8'd134} : s = 113;
	{8'd196,8'd135} : s = 242;
	{8'd196,8'd136} : s = 108;
	{8'd196,8'd137} : s = 241;
	{8'd196,8'd138} : s = 236;
	{8'd196,8'd139} : s = 399;
	{8'd196,8'd140} : s = 26;
	{8'd196,8'd141} : s = 106;
	{8'd196,8'd142} : s = 105;
	{8'd196,8'd143} : s = 234;
	{8'd196,8'd144} : s = 102;
	{8'd196,8'd145} : s = 233;
	{8'd196,8'd146} : s = 230;
	{8'd196,8'd147} : s = 380;
	{8'd196,8'd148} : s = 101;
	{8'd196,8'd149} : s = 229;
	{8'd196,8'd150} : s = 227;
	{8'd196,8'd151} : s = 378;
	{8'd196,8'd152} : s = 220;
	{8'd196,8'd153} : s = 377;
	{8'd196,8'd154} : s = 374;
	{8'd196,8'd155} : s = 487;
	{8'd196,8'd156} : s = 25;
	{8'd196,8'd157} : s = 99;
	{8'd196,8'd158} : s = 92;
	{8'd196,8'd159} : s = 218;
	{8'd196,8'd160} : s = 90;
	{8'd196,8'd161} : s = 217;
	{8'd196,8'd162} : s = 214;
	{8'd196,8'd163} : s = 373;
	{8'd196,8'd164} : s = 89;
	{8'd196,8'd165} : s = 213;
	{8'd196,8'd166} : s = 211;
	{8'd196,8'd167} : s = 371;
	{8'd196,8'd168} : s = 206;
	{8'd196,8'd169} : s = 366;
	{8'd196,8'd170} : s = 365;
	{8'd196,8'd171} : s = 478;
	{8'd196,8'd172} : s = 86;
	{8'd196,8'd173} : s = 205;
	{8'd196,8'd174} : s = 203;
	{8'd196,8'd175} : s = 363;
	{8'd196,8'd176} : s = 199;
	{8'd196,8'd177} : s = 359;
	{8'd196,8'd178} : s = 350;
	{8'd196,8'd179} : s = 477;
	{8'd196,8'd180} : s = 188;
	{8'd196,8'd181} : s = 349;
	{8'd196,8'd182} : s = 347;
	{8'd196,8'd183} : s = 475;
	{8'd196,8'd184} : s = 343;
	{8'd196,8'd185} : s = 471;
	{8'd196,8'd186} : s = 463;
	{8'd196,8'd187} : s = 509;
	{8'd196,8'd188} : s = 3;
	{8'd196,8'd189} : s = 22;
	{8'd196,8'd190} : s = 21;
	{8'd196,8'd191} : s = 85;
	{8'd196,8'd192} : s = 19;
	{8'd196,8'd193} : s = 83;
	{8'd196,8'd194} : s = 78;
	{8'd196,8'd195} : s = 186;
	{8'd196,8'd196} : s = 14;
	{8'd196,8'd197} : s = 77;
	{8'd196,8'd198} : s = 75;
	{8'd196,8'd199} : s = 185;
	{8'd196,8'd200} : s = 71;
	{8'd196,8'd201} : s = 182;
	{8'd196,8'd202} : s = 181;
	{8'd196,8'd203} : s = 335;
	{8'd196,8'd204} : s = 13;
	{8'd196,8'd205} : s = 60;
	{8'd196,8'd206} : s = 58;
	{8'd196,8'd207} : s = 179;
	{8'd196,8'd208} : s = 57;
	{8'd196,8'd209} : s = 174;
	{8'd196,8'd210} : s = 173;
	{8'd196,8'd211} : s = 318;
	{8'd196,8'd212} : s = 54;
	{8'd196,8'd213} : s = 171;
	{8'd196,8'd214} : s = 167;
	{8'd196,8'd215} : s = 317;
	{8'd196,8'd216} : s = 158;
	{8'd196,8'd217} : s = 315;
	{8'd196,8'd218} : s = 311;
	{8'd196,8'd219} : s = 446;
	{8'd196,8'd220} : s = 11;
	{8'd196,8'd221} : s = 53;
	{8'd196,8'd222} : s = 51;
	{8'd196,8'd223} : s = 157;
	{8'd196,8'd224} : s = 46;
	{8'd196,8'd225} : s = 155;
	{8'd196,8'd226} : s = 151;
	{8'd196,8'd227} : s = 303;
	{8'd196,8'd228} : s = 45;
	{8'd196,8'd229} : s = 143;
	{8'd196,8'd230} : s = 124;
	{8'd196,8'd231} : s = 287;
	{8'd196,8'd232} : s = 122;
	{8'd196,8'd233} : s = 252;
	{8'd196,8'd234} : s = 250;
	{8'd196,8'd235} : s = 445;
	{8'd196,8'd236} : s = 43;
	{8'd196,8'd237} : s = 121;
	{8'd196,8'd238} : s = 118;
	{8'd196,8'd239} : s = 249;
	{8'd196,8'd240} : s = 117;
	{8'd196,8'd241} : s = 246;
	{8'd196,8'd242} : s = 245;
	{8'd196,8'd243} : s = 443;
	{8'd196,8'd244} : s = 115;
	{8'd196,8'd245} : s = 243;
	{8'd196,8'd246} : s = 238;
	{8'd196,8'd247} : s = 439;
	{8'd196,8'd248} : s = 237;
	{8'd196,8'd249} : s = 431;
	{8'd196,8'd250} : s = 415;
	{8'd196,8'd251} : s = 507;
	{8'd196,8'd252} : s = 7;
	{8'd196,8'd253} : s = 39;
	{8'd196,8'd254} : s = 30;
	{8'd196,8'd255} : s = 110;
	{8'd197,8'd0} : s = 240;
	{8'd197,8'd1} : s = 232;
	{8'd197,8'd2} : s = 372;
	{8'd197,8'd3} : s = 97;
	{8'd197,8'd4} : s = 228;
	{8'd197,8'd5} : s = 226;
	{8'd197,8'd6} : s = 370;
	{8'd197,8'd7} : s = 225;
	{8'd197,8'd8} : s = 369;
	{8'd197,8'd9} : s = 364;
	{8'd197,8'd10} : s = 470;
	{8'd197,8'd11} : s = 88;
	{8'd197,8'd12} : s = 216;
	{8'd197,8'd13} : s = 212;
	{8'd197,8'd14} : s = 362;
	{8'd197,8'd15} : s = 210;
	{8'd197,8'd16} : s = 361;
	{8'd197,8'd17} : s = 358;
	{8'd197,8'd18} : s = 469;
	{8'd197,8'd19} : s = 209;
	{8'd197,8'd20} : s = 357;
	{8'd197,8'd21} : s = 355;
	{8'd197,8'd22} : s = 467;
	{8'd197,8'd23} : s = 348;
	{8'd197,8'd24} : s = 462;
	{8'd197,8'd25} : s = 461;
	{8'd197,8'd26} : s = 505;
	{8'd197,8'd27} : s = 84;
	{8'd197,8'd28} : s = 204;
	{8'd197,8'd29} : s = 202;
	{8'd197,8'd30} : s = 346;
	{8'd197,8'd31} : s = 201;
	{8'd197,8'd32} : s = 345;
	{8'd197,8'd33} : s = 342;
	{8'd197,8'd34} : s = 459;
	{8'd197,8'd35} : s = 198;
	{8'd197,8'd36} : s = 341;
	{8'd197,8'd37} : s = 339;
	{8'd197,8'd38} : s = 455;
	{8'd197,8'd39} : s = 334;
	{8'd197,8'd40} : s = 444;
	{8'd197,8'd41} : s = 442;
	{8'd197,8'd42} : s = 502;
	{8'd197,8'd43} : s = 197;
	{8'd197,8'd44} : s = 333;
	{8'd197,8'd45} : s = 331;
	{8'd197,8'd46} : s = 441;
	{8'd197,8'd47} : s = 327;
	{8'd197,8'd48} : s = 438;
	{8'd197,8'd49} : s = 437;
	{8'd197,8'd50} : s = 501;
	{8'd197,8'd51} : s = 316;
	{8'd197,8'd52} : s = 435;
	{8'd197,8'd53} : s = 430;
	{8'd197,8'd54} : s = 499;
	{8'd197,8'd55} : s = 429;
	{8'd197,8'd56} : s = 494;
	{8'd197,8'd57} : s = 493;
	{8'd197,8'd58} : s = 510;
	{8'd197,8'd59} : s = 1;
	{8'd197,8'd60} : s = 18;
	{8'd197,8'd61} : s = 17;
	{8'd197,8'd62} : s = 82;
	{8'd197,8'd63} : s = 12;
	{8'd197,8'd64} : s = 81;
	{8'd197,8'd65} : s = 76;
	{8'd197,8'd66} : s = 195;
	{8'd197,8'd67} : s = 10;
	{8'd197,8'd68} : s = 74;
	{8'd197,8'd69} : s = 73;
	{8'd197,8'd70} : s = 184;
	{8'd197,8'd71} : s = 70;
	{8'd197,8'd72} : s = 180;
	{8'd197,8'd73} : s = 178;
	{8'd197,8'd74} : s = 314;
	{8'd197,8'd75} : s = 9;
	{8'd197,8'd76} : s = 69;
	{8'd197,8'd77} : s = 67;
	{8'd197,8'd78} : s = 177;
	{8'd197,8'd79} : s = 56;
	{8'd197,8'd80} : s = 172;
	{8'd197,8'd81} : s = 170;
	{8'd197,8'd82} : s = 313;
	{8'd197,8'd83} : s = 52;
	{8'd197,8'd84} : s = 169;
	{8'd197,8'd85} : s = 166;
	{8'd197,8'd86} : s = 310;
	{8'd197,8'd87} : s = 165;
	{8'd197,8'd88} : s = 309;
	{8'd197,8'd89} : s = 307;
	{8'd197,8'd90} : s = 427;
	{8'd197,8'd91} : s = 6;
	{8'd197,8'd92} : s = 50;
	{8'd197,8'd93} : s = 49;
	{8'd197,8'd94} : s = 163;
	{8'd197,8'd95} : s = 44;
	{8'd197,8'd96} : s = 156;
	{8'd197,8'd97} : s = 154;
	{8'd197,8'd98} : s = 302;
	{8'd197,8'd99} : s = 42;
	{8'd197,8'd100} : s = 153;
	{8'd197,8'd101} : s = 150;
	{8'd197,8'd102} : s = 301;
	{8'd197,8'd103} : s = 149;
	{8'd197,8'd104} : s = 299;
	{8'd197,8'd105} : s = 295;
	{8'd197,8'd106} : s = 423;
	{8'd197,8'd107} : s = 41;
	{8'd197,8'd108} : s = 147;
	{8'd197,8'd109} : s = 142;
	{8'd197,8'd110} : s = 286;
	{8'd197,8'd111} : s = 141;
	{8'd197,8'd112} : s = 285;
	{8'd197,8'd113} : s = 283;
	{8'd197,8'd114} : s = 414;
	{8'd197,8'd115} : s = 139;
	{8'd197,8'd116} : s = 279;
	{8'd197,8'd117} : s = 271;
	{8'd197,8'd118} : s = 413;
	{8'd197,8'd119} : s = 248;
	{8'd197,8'd120} : s = 411;
	{8'd197,8'd121} : s = 407;
	{8'd197,8'd122} : s = 491;
	{8'd197,8'd123} : s = 5;
	{8'd197,8'd124} : s = 38;
	{8'd197,8'd125} : s = 37;
	{8'd197,8'd126} : s = 135;
	{8'd197,8'd127} : s = 35;
	{8'd197,8'd128} : s = 120;
	{8'd197,8'd129} : s = 116;
	{8'd197,8'd130} : s = 244;
	{8'd197,8'd131} : s = 28;
	{8'd197,8'd132} : s = 114;
	{8'd197,8'd133} : s = 113;
	{8'd197,8'd134} : s = 242;
	{8'd197,8'd135} : s = 108;
	{8'd197,8'd136} : s = 241;
	{8'd197,8'd137} : s = 236;
	{8'd197,8'd138} : s = 399;
	{8'd197,8'd139} : s = 26;
	{8'd197,8'd140} : s = 106;
	{8'd197,8'd141} : s = 105;
	{8'd197,8'd142} : s = 234;
	{8'd197,8'd143} : s = 102;
	{8'd197,8'd144} : s = 233;
	{8'd197,8'd145} : s = 230;
	{8'd197,8'd146} : s = 380;
	{8'd197,8'd147} : s = 101;
	{8'd197,8'd148} : s = 229;
	{8'd197,8'd149} : s = 227;
	{8'd197,8'd150} : s = 378;
	{8'd197,8'd151} : s = 220;
	{8'd197,8'd152} : s = 377;
	{8'd197,8'd153} : s = 374;
	{8'd197,8'd154} : s = 487;
	{8'd197,8'd155} : s = 25;
	{8'd197,8'd156} : s = 99;
	{8'd197,8'd157} : s = 92;
	{8'd197,8'd158} : s = 218;
	{8'd197,8'd159} : s = 90;
	{8'd197,8'd160} : s = 217;
	{8'd197,8'd161} : s = 214;
	{8'd197,8'd162} : s = 373;
	{8'd197,8'd163} : s = 89;
	{8'd197,8'd164} : s = 213;
	{8'd197,8'd165} : s = 211;
	{8'd197,8'd166} : s = 371;
	{8'd197,8'd167} : s = 206;
	{8'd197,8'd168} : s = 366;
	{8'd197,8'd169} : s = 365;
	{8'd197,8'd170} : s = 478;
	{8'd197,8'd171} : s = 86;
	{8'd197,8'd172} : s = 205;
	{8'd197,8'd173} : s = 203;
	{8'd197,8'd174} : s = 363;
	{8'd197,8'd175} : s = 199;
	{8'd197,8'd176} : s = 359;
	{8'd197,8'd177} : s = 350;
	{8'd197,8'd178} : s = 477;
	{8'd197,8'd179} : s = 188;
	{8'd197,8'd180} : s = 349;
	{8'd197,8'd181} : s = 347;
	{8'd197,8'd182} : s = 475;
	{8'd197,8'd183} : s = 343;
	{8'd197,8'd184} : s = 471;
	{8'd197,8'd185} : s = 463;
	{8'd197,8'd186} : s = 509;
	{8'd197,8'd187} : s = 3;
	{8'd197,8'd188} : s = 22;
	{8'd197,8'd189} : s = 21;
	{8'd197,8'd190} : s = 85;
	{8'd197,8'd191} : s = 19;
	{8'd197,8'd192} : s = 83;
	{8'd197,8'd193} : s = 78;
	{8'd197,8'd194} : s = 186;
	{8'd197,8'd195} : s = 14;
	{8'd197,8'd196} : s = 77;
	{8'd197,8'd197} : s = 75;
	{8'd197,8'd198} : s = 185;
	{8'd197,8'd199} : s = 71;
	{8'd197,8'd200} : s = 182;
	{8'd197,8'd201} : s = 181;
	{8'd197,8'd202} : s = 335;
	{8'd197,8'd203} : s = 13;
	{8'd197,8'd204} : s = 60;
	{8'd197,8'd205} : s = 58;
	{8'd197,8'd206} : s = 179;
	{8'd197,8'd207} : s = 57;
	{8'd197,8'd208} : s = 174;
	{8'd197,8'd209} : s = 173;
	{8'd197,8'd210} : s = 318;
	{8'd197,8'd211} : s = 54;
	{8'd197,8'd212} : s = 171;
	{8'd197,8'd213} : s = 167;
	{8'd197,8'd214} : s = 317;
	{8'd197,8'd215} : s = 158;
	{8'd197,8'd216} : s = 315;
	{8'd197,8'd217} : s = 311;
	{8'd197,8'd218} : s = 446;
	{8'd197,8'd219} : s = 11;
	{8'd197,8'd220} : s = 53;
	{8'd197,8'd221} : s = 51;
	{8'd197,8'd222} : s = 157;
	{8'd197,8'd223} : s = 46;
	{8'd197,8'd224} : s = 155;
	{8'd197,8'd225} : s = 151;
	{8'd197,8'd226} : s = 303;
	{8'd197,8'd227} : s = 45;
	{8'd197,8'd228} : s = 143;
	{8'd197,8'd229} : s = 124;
	{8'd197,8'd230} : s = 287;
	{8'd197,8'd231} : s = 122;
	{8'd197,8'd232} : s = 252;
	{8'd197,8'd233} : s = 250;
	{8'd197,8'd234} : s = 445;
	{8'd197,8'd235} : s = 43;
	{8'd197,8'd236} : s = 121;
	{8'd197,8'd237} : s = 118;
	{8'd197,8'd238} : s = 249;
	{8'd197,8'd239} : s = 117;
	{8'd197,8'd240} : s = 246;
	{8'd197,8'd241} : s = 245;
	{8'd197,8'd242} : s = 443;
	{8'd197,8'd243} : s = 115;
	{8'd197,8'd244} : s = 243;
	{8'd197,8'd245} : s = 238;
	{8'd197,8'd246} : s = 439;
	{8'd197,8'd247} : s = 237;
	{8'd197,8'd248} : s = 431;
	{8'd197,8'd249} : s = 415;
	{8'd197,8'd250} : s = 507;
	{8'd197,8'd251} : s = 7;
	{8'd197,8'd252} : s = 39;
	{8'd197,8'd253} : s = 30;
	{8'd197,8'd254} : s = 110;
	{8'd197,8'd255} : s = 29;
	{8'd198,8'd0} : s = 232;
	{8'd198,8'd1} : s = 372;
	{8'd198,8'd2} : s = 97;
	{8'd198,8'd3} : s = 228;
	{8'd198,8'd4} : s = 226;
	{8'd198,8'd5} : s = 370;
	{8'd198,8'd6} : s = 225;
	{8'd198,8'd7} : s = 369;
	{8'd198,8'd8} : s = 364;
	{8'd198,8'd9} : s = 470;
	{8'd198,8'd10} : s = 88;
	{8'd198,8'd11} : s = 216;
	{8'd198,8'd12} : s = 212;
	{8'd198,8'd13} : s = 362;
	{8'd198,8'd14} : s = 210;
	{8'd198,8'd15} : s = 361;
	{8'd198,8'd16} : s = 358;
	{8'd198,8'd17} : s = 469;
	{8'd198,8'd18} : s = 209;
	{8'd198,8'd19} : s = 357;
	{8'd198,8'd20} : s = 355;
	{8'd198,8'd21} : s = 467;
	{8'd198,8'd22} : s = 348;
	{8'd198,8'd23} : s = 462;
	{8'd198,8'd24} : s = 461;
	{8'd198,8'd25} : s = 505;
	{8'd198,8'd26} : s = 84;
	{8'd198,8'd27} : s = 204;
	{8'd198,8'd28} : s = 202;
	{8'd198,8'd29} : s = 346;
	{8'd198,8'd30} : s = 201;
	{8'd198,8'd31} : s = 345;
	{8'd198,8'd32} : s = 342;
	{8'd198,8'd33} : s = 459;
	{8'd198,8'd34} : s = 198;
	{8'd198,8'd35} : s = 341;
	{8'd198,8'd36} : s = 339;
	{8'd198,8'd37} : s = 455;
	{8'd198,8'd38} : s = 334;
	{8'd198,8'd39} : s = 444;
	{8'd198,8'd40} : s = 442;
	{8'd198,8'd41} : s = 502;
	{8'd198,8'd42} : s = 197;
	{8'd198,8'd43} : s = 333;
	{8'd198,8'd44} : s = 331;
	{8'd198,8'd45} : s = 441;
	{8'd198,8'd46} : s = 327;
	{8'd198,8'd47} : s = 438;
	{8'd198,8'd48} : s = 437;
	{8'd198,8'd49} : s = 501;
	{8'd198,8'd50} : s = 316;
	{8'd198,8'd51} : s = 435;
	{8'd198,8'd52} : s = 430;
	{8'd198,8'd53} : s = 499;
	{8'd198,8'd54} : s = 429;
	{8'd198,8'd55} : s = 494;
	{8'd198,8'd56} : s = 493;
	{8'd198,8'd57} : s = 510;
	{8'd198,8'd58} : s = 1;
	{8'd198,8'd59} : s = 18;
	{8'd198,8'd60} : s = 17;
	{8'd198,8'd61} : s = 82;
	{8'd198,8'd62} : s = 12;
	{8'd198,8'd63} : s = 81;
	{8'd198,8'd64} : s = 76;
	{8'd198,8'd65} : s = 195;
	{8'd198,8'd66} : s = 10;
	{8'd198,8'd67} : s = 74;
	{8'd198,8'd68} : s = 73;
	{8'd198,8'd69} : s = 184;
	{8'd198,8'd70} : s = 70;
	{8'd198,8'd71} : s = 180;
	{8'd198,8'd72} : s = 178;
	{8'd198,8'd73} : s = 314;
	{8'd198,8'd74} : s = 9;
	{8'd198,8'd75} : s = 69;
	{8'd198,8'd76} : s = 67;
	{8'd198,8'd77} : s = 177;
	{8'd198,8'd78} : s = 56;
	{8'd198,8'd79} : s = 172;
	{8'd198,8'd80} : s = 170;
	{8'd198,8'd81} : s = 313;
	{8'd198,8'd82} : s = 52;
	{8'd198,8'd83} : s = 169;
	{8'd198,8'd84} : s = 166;
	{8'd198,8'd85} : s = 310;
	{8'd198,8'd86} : s = 165;
	{8'd198,8'd87} : s = 309;
	{8'd198,8'd88} : s = 307;
	{8'd198,8'd89} : s = 427;
	{8'd198,8'd90} : s = 6;
	{8'd198,8'd91} : s = 50;
	{8'd198,8'd92} : s = 49;
	{8'd198,8'd93} : s = 163;
	{8'd198,8'd94} : s = 44;
	{8'd198,8'd95} : s = 156;
	{8'd198,8'd96} : s = 154;
	{8'd198,8'd97} : s = 302;
	{8'd198,8'd98} : s = 42;
	{8'd198,8'd99} : s = 153;
	{8'd198,8'd100} : s = 150;
	{8'd198,8'd101} : s = 301;
	{8'd198,8'd102} : s = 149;
	{8'd198,8'd103} : s = 299;
	{8'd198,8'd104} : s = 295;
	{8'd198,8'd105} : s = 423;
	{8'd198,8'd106} : s = 41;
	{8'd198,8'd107} : s = 147;
	{8'd198,8'd108} : s = 142;
	{8'd198,8'd109} : s = 286;
	{8'd198,8'd110} : s = 141;
	{8'd198,8'd111} : s = 285;
	{8'd198,8'd112} : s = 283;
	{8'd198,8'd113} : s = 414;
	{8'd198,8'd114} : s = 139;
	{8'd198,8'd115} : s = 279;
	{8'd198,8'd116} : s = 271;
	{8'd198,8'd117} : s = 413;
	{8'd198,8'd118} : s = 248;
	{8'd198,8'd119} : s = 411;
	{8'd198,8'd120} : s = 407;
	{8'd198,8'd121} : s = 491;
	{8'd198,8'd122} : s = 5;
	{8'd198,8'd123} : s = 38;
	{8'd198,8'd124} : s = 37;
	{8'd198,8'd125} : s = 135;
	{8'd198,8'd126} : s = 35;
	{8'd198,8'd127} : s = 120;
	{8'd198,8'd128} : s = 116;
	{8'd198,8'd129} : s = 244;
	{8'd198,8'd130} : s = 28;
	{8'd198,8'd131} : s = 114;
	{8'd198,8'd132} : s = 113;
	{8'd198,8'd133} : s = 242;
	{8'd198,8'd134} : s = 108;
	{8'd198,8'd135} : s = 241;
	{8'd198,8'd136} : s = 236;
	{8'd198,8'd137} : s = 399;
	{8'd198,8'd138} : s = 26;
	{8'd198,8'd139} : s = 106;
	{8'd198,8'd140} : s = 105;
	{8'd198,8'd141} : s = 234;
	{8'd198,8'd142} : s = 102;
	{8'd198,8'd143} : s = 233;
	{8'd198,8'd144} : s = 230;
	{8'd198,8'd145} : s = 380;
	{8'd198,8'd146} : s = 101;
	{8'd198,8'd147} : s = 229;
	{8'd198,8'd148} : s = 227;
	{8'd198,8'd149} : s = 378;
	{8'd198,8'd150} : s = 220;
	{8'd198,8'd151} : s = 377;
	{8'd198,8'd152} : s = 374;
	{8'd198,8'd153} : s = 487;
	{8'd198,8'd154} : s = 25;
	{8'd198,8'd155} : s = 99;
	{8'd198,8'd156} : s = 92;
	{8'd198,8'd157} : s = 218;
	{8'd198,8'd158} : s = 90;
	{8'd198,8'd159} : s = 217;
	{8'd198,8'd160} : s = 214;
	{8'd198,8'd161} : s = 373;
	{8'd198,8'd162} : s = 89;
	{8'd198,8'd163} : s = 213;
	{8'd198,8'd164} : s = 211;
	{8'd198,8'd165} : s = 371;
	{8'd198,8'd166} : s = 206;
	{8'd198,8'd167} : s = 366;
	{8'd198,8'd168} : s = 365;
	{8'd198,8'd169} : s = 478;
	{8'd198,8'd170} : s = 86;
	{8'd198,8'd171} : s = 205;
	{8'd198,8'd172} : s = 203;
	{8'd198,8'd173} : s = 363;
	{8'd198,8'd174} : s = 199;
	{8'd198,8'd175} : s = 359;
	{8'd198,8'd176} : s = 350;
	{8'd198,8'd177} : s = 477;
	{8'd198,8'd178} : s = 188;
	{8'd198,8'd179} : s = 349;
	{8'd198,8'd180} : s = 347;
	{8'd198,8'd181} : s = 475;
	{8'd198,8'd182} : s = 343;
	{8'd198,8'd183} : s = 471;
	{8'd198,8'd184} : s = 463;
	{8'd198,8'd185} : s = 509;
	{8'd198,8'd186} : s = 3;
	{8'd198,8'd187} : s = 22;
	{8'd198,8'd188} : s = 21;
	{8'd198,8'd189} : s = 85;
	{8'd198,8'd190} : s = 19;
	{8'd198,8'd191} : s = 83;
	{8'd198,8'd192} : s = 78;
	{8'd198,8'd193} : s = 186;
	{8'd198,8'd194} : s = 14;
	{8'd198,8'd195} : s = 77;
	{8'd198,8'd196} : s = 75;
	{8'd198,8'd197} : s = 185;
	{8'd198,8'd198} : s = 71;
	{8'd198,8'd199} : s = 182;
	{8'd198,8'd200} : s = 181;
	{8'd198,8'd201} : s = 335;
	{8'd198,8'd202} : s = 13;
	{8'd198,8'd203} : s = 60;
	{8'd198,8'd204} : s = 58;
	{8'd198,8'd205} : s = 179;
	{8'd198,8'd206} : s = 57;
	{8'd198,8'd207} : s = 174;
	{8'd198,8'd208} : s = 173;
	{8'd198,8'd209} : s = 318;
	{8'd198,8'd210} : s = 54;
	{8'd198,8'd211} : s = 171;
	{8'd198,8'd212} : s = 167;
	{8'd198,8'd213} : s = 317;
	{8'd198,8'd214} : s = 158;
	{8'd198,8'd215} : s = 315;
	{8'd198,8'd216} : s = 311;
	{8'd198,8'd217} : s = 446;
	{8'd198,8'd218} : s = 11;
	{8'd198,8'd219} : s = 53;
	{8'd198,8'd220} : s = 51;
	{8'd198,8'd221} : s = 157;
	{8'd198,8'd222} : s = 46;
	{8'd198,8'd223} : s = 155;
	{8'd198,8'd224} : s = 151;
	{8'd198,8'd225} : s = 303;
	{8'd198,8'd226} : s = 45;
	{8'd198,8'd227} : s = 143;
	{8'd198,8'd228} : s = 124;
	{8'd198,8'd229} : s = 287;
	{8'd198,8'd230} : s = 122;
	{8'd198,8'd231} : s = 252;
	{8'd198,8'd232} : s = 250;
	{8'd198,8'd233} : s = 445;
	{8'd198,8'd234} : s = 43;
	{8'd198,8'd235} : s = 121;
	{8'd198,8'd236} : s = 118;
	{8'd198,8'd237} : s = 249;
	{8'd198,8'd238} : s = 117;
	{8'd198,8'd239} : s = 246;
	{8'd198,8'd240} : s = 245;
	{8'd198,8'd241} : s = 443;
	{8'd198,8'd242} : s = 115;
	{8'd198,8'd243} : s = 243;
	{8'd198,8'd244} : s = 238;
	{8'd198,8'd245} : s = 439;
	{8'd198,8'd246} : s = 237;
	{8'd198,8'd247} : s = 431;
	{8'd198,8'd248} : s = 415;
	{8'd198,8'd249} : s = 507;
	{8'd198,8'd250} : s = 7;
	{8'd198,8'd251} : s = 39;
	{8'd198,8'd252} : s = 30;
	{8'd198,8'd253} : s = 110;
	{8'd198,8'd254} : s = 29;
	{8'd198,8'd255} : s = 109;
	{8'd199,8'd0} : s = 372;
	{8'd199,8'd1} : s = 97;
	{8'd199,8'd2} : s = 228;
	{8'd199,8'd3} : s = 226;
	{8'd199,8'd4} : s = 370;
	{8'd199,8'd5} : s = 225;
	{8'd199,8'd6} : s = 369;
	{8'd199,8'd7} : s = 364;
	{8'd199,8'd8} : s = 470;
	{8'd199,8'd9} : s = 88;
	{8'd199,8'd10} : s = 216;
	{8'd199,8'd11} : s = 212;
	{8'd199,8'd12} : s = 362;
	{8'd199,8'd13} : s = 210;
	{8'd199,8'd14} : s = 361;
	{8'd199,8'd15} : s = 358;
	{8'd199,8'd16} : s = 469;
	{8'd199,8'd17} : s = 209;
	{8'd199,8'd18} : s = 357;
	{8'd199,8'd19} : s = 355;
	{8'd199,8'd20} : s = 467;
	{8'd199,8'd21} : s = 348;
	{8'd199,8'd22} : s = 462;
	{8'd199,8'd23} : s = 461;
	{8'd199,8'd24} : s = 505;
	{8'd199,8'd25} : s = 84;
	{8'd199,8'd26} : s = 204;
	{8'd199,8'd27} : s = 202;
	{8'd199,8'd28} : s = 346;
	{8'd199,8'd29} : s = 201;
	{8'd199,8'd30} : s = 345;
	{8'd199,8'd31} : s = 342;
	{8'd199,8'd32} : s = 459;
	{8'd199,8'd33} : s = 198;
	{8'd199,8'd34} : s = 341;
	{8'd199,8'd35} : s = 339;
	{8'd199,8'd36} : s = 455;
	{8'd199,8'd37} : s = 334;
	{8'd199,8'd38} : s = 444;
	{8'd199,8'd39} : s = 442;
	{8'd199,8'd40} : s = 502;
	{8'd199,8'd41} : s = 197;
	{8'd199,8'd42} : s = 333;
	{8'd199,8'd43} : s = 331;
	{8'd199,8'd44} : s = 441;
	{8'd199,8'd45} : s = 327;
	{8'd199,8'd46} : s = 438;
	{8'd199,8'd47} : s = 437;
	{8'd199,8'd48} : s = 501;
	{8'd199,8'd49} : s = 316;
	{8'd199,8'd50} : s = 435;
	{8'd199,8'd51} : s = 430;
	{8'd199,8'd52} : s = 499;
	{8'd199,8'd53} : s = 429;
	{8'd199,8'd54} : s = 494;
	{8'd199,8'd55} : s = 493;
	{8'd199,8'd56} : s = 510;
	{8'd199,8'd57} : s = 1;
	{8'd199,8'd58} : s = 18;
	{8'd199,8'd59} : s = 17;
	{8'd199,8'd60} : s = 82;
	{8'd199,8'd61} : s = 12;
	{8'd199,8'd62} : s = 81;
	{8'd199,8'd63} : s = 76;
	{8'd199,8'd64} : s = 195;
	{8'd199,8'd65} : s = 10;
	{8'd199,8'd66} : s = 74;
	{8'd199,8'd67} : s = 73;
	{8'd199,8'd68} : s = 184;
	{8'd199,8'd69} : s = 70;
	{8'd199,8'd70} : s = 180;
	{8'd199,8'd71} : s = 178;
	{8'd199,8'd72} : s = 314;
	{8'd199,8'd73} : s = 9;
	{8'd199,8'd74} : s = 69;
	{8'd199,8'd75} : s = 67;
	{8'd199,8'd76} : s = 177;
	{8'd199,8'd77} : s = 56;
	{8'd199,8'd78} : s = 172;
	{8'd199,8'd79} : s = 170;
	{8'd199,8'd80} : s = 313;
	{8'd199,8'd81} : s = 52;
	{8'd199,8'd82} : s = 169;
	{8'd199,8'd83} : s = 166;
	{8'd199,8'd84} : s = 310;
	{8'd199,8'd85} : s = 165;
	{8'd199,8'd86} : s = 309;
	{8'd199,8'd87} : s = 307;
	{8'd199,8'd88} : s = 427;
	{8'd199,8'd89} : s = 6;
	{8'd199,8'd90} : s = 50;
	{8'd199,8'd91} : s = 49;
	{8'd199,8'd92} : s = 163;
	{8'd199,8'd93} : s = 44;
	{8'd199,8'd94} : s = 156;
	{8'd199,8'd95} : s = 154;
	{8'd199,8'd96} : s = 302;
	{8'd199,8'd97} : s = 42;
	{8'd199,8'd98} : s = 153;
	{8'd199,8'd99} : s = 150;
	{8'd199,8'd100} : s = 301;
	{8'd199,8'd101} : s = 149;
	{8'd199,8'd102} : s = 299;
	{8'd199,8'd103} : s = 295;
	{8'd199,8'd104} : s = 423;
	{8'd199,8'd105} : s = 41;
	{8'd199,8'd106} : s = 147;
	{8'd199,8'd107} : s = 142;
	{8'd199,8'd108} : s = 286;
	{8'd199,8'd109} : s = 141;
	{8'd199,8'd110} : s = 285;
	{8'd199,8'd111} : s = 283;
	{8'd199,8'd112} : s = 414;
	{8'd199,8'd113} : s = 139;
	{8'd199,8'd114} : s = 279;
	{8'd199,8'd115} : s = 271;
	{8'd199,8'd116} : s = 413;
	{8'd199,8'd117} : s = 248;
	{8'd199,8'd118} : s = 411;
	{8'd199,8'd119} : s = 407;
	{8'd199,8'd120} : s = 491;
	{8'd199,8'd121} : s = 5;
	{8'd199,8'd122} : s = 38;
	{8'd199,8'd123} : s = 37;
	{8'd199,8'd124} : s = 135;
	{8'd199,8'd125} : s = 35;
	{8'd199,8'd126} : s = 120;
	{8'd199,8'd127} : s = 116;
	{8'd199,8'd128} : s = 244;
	{8'd199,8'd129} : s = 28;
	{8'd199,8'd130} : s = 114;
	{8'd199,8'd131} : s = 113;
	{8'd199,8'd132} : s = 242;
	{8'd199,8'd133} : s = 108;
	{8'd199,8'd134} : s = 241;
	{8'd199,8'd135} : s = 236;
	{8'd199,8'd136} : s = 399;
	{8'd199,8'd137} : s = 26;
	{8'd199,8'd138} : s = 106;
	{8'd199,8'd139} : s = 105;
	{8'd199,8'd140} : s = 234;
	{8'd199,8'd141} : s = 102;
	{8'd199,8'd142} : s = 233;
	{8'd199,8'd143} : s = 230;
	{8'd199,8'd144} : s = 380;
	{8'd199,8'd145} : s = 101;
	{8'd199,8'd146} : s = 229;
	{8'd199,8'd147} : s = 227;
	{8'd199,8'd148} : s = 378;
	{8'd199,8'd149} : s = 220;
	{8'd199,8'd150} : s = 377;
	{8'd199,8'd151} : s = 374;
	{8'd199,8'd152} : s = 487;
	{8'd199,8'd153} : s = 25;
	{8'd199,8'd154} : s = 99;
	{8'd199,8'd155} : s = 92;
	{8'd199,8'd156} : s = 218;
	{8'd199,8'd157} : s = 90;
	{8'd199,8'd158} : s = 217;
	{8'd199,8'd159} : s = 214;
	{8'd199,8'd160} : s = 373;
	{8'd199,8'd161} : s = 89;
	{8'd199,8'd162} : s = 213;
	{8'd199,8'd163} : s = 211;
	{8'd199,8'd164} : s = 371;
	{8'd199,8'd165} : s = 206;
	{8'd199,8'd166} : s = 366;
	{8'd199,8'd167} : s = 365;
	{8'd199,8'd168} : s = 478;
	{8'd199,8'd169} : s = 86;
	{8'd199,8'd170} : s = 205;
	{8'd199,8'd171} : s = 203;
	{8'd199,8'd172} : s = 363;
	{8'd199,8'd173} : s = 199;
	{8'd199,8'd174} : s = 359;
	{8'd199,8'd175} : s = 350;
	{8'd199,8'd176} : s = 477;
	{8'd199,8'd177} : s = 188;
	{8'd199,8'd178} : s = 349;
	{8'd199,8'd179} : s = 347;
	{8'd199,8'd180} : s = 475;
	{8'd199,8'd181} : s = 343;
	{8'd199,8'd182} : s = 471;
	{8'd199,8'd183} : s = 463;
	{8'd199,8'd184} : s = 509;
	{8'd199,8'd185} : s = 3;
	{8'd199,8'd186} : s = 22;
	{8'd199,8'd187} : s = 21;
	{8'd199,8'd188} : s = 85;
	{8'd199,8'd189} : s = 19;
	{8'd199,8'd190} : s = 83;
	{8'd199,8'd191} : s = 78;
	{8'd199,8'd192} : s = 186;
	{8'd199,8'd193} : s = 14;
	{8'd199,8'd194} : s = 77;
	{8'd199,8'd195} : s = 75;
	{8'd199,8'd196} : s = 185;
	{8'd199,8'd197} : s = 71;
	{8'd199,8'd198} : s = 182;
	{8'd199,8'd199} : s = 181;
	{8'd199,8'd200} : s = 335;
	{8'd199,8'd201} : s = 13;
	{8'd199,8'd202} : s = 60;
	{8'd199,8'd203} : s = 58;
	{8'd199,8'd204} : s = 179;
	{8'd199,8'd205} : s = 57;
	{8'd199,8'd206} : s = 174;
	{8'd199,8'd207} : s = 173;
	{8'd199,8'd208} : s = 318;
	{8'd199,8'd209} : s = 54;
	{8'd199,8'd210} : s = 171;
	{8'd199,8'd211} : s = 167;
	{8'd199,8'd212} : s = 317;
	{8'd199,8'd213} : s = 158;
	{8'd199,8'd214} : s = 315;
	{8'd199,8'd215} : s = 311;
	{8'd199,8'd216} : s = 446;
	{8'd199,8'd217} : s = 11;
	{8'd199,8'd218} : s = 53;
	{8'd199,8'd219} : s = 51;
	{8'd199,8'd220} : s = 157;
	{8'd199,8'd221} : s = 46;
	{8'd199,8'd222} : s = 155;
	{8'd199,8'd223} : s = 151;
	{8'd199,8'd224} : s = 303;
	{8'd199,8'd225} : s = 45;
	{8'd199,8'd226} : s = 143;
	{8'd199,8'd227} : s = 124;
	{8'd199,8'd228} : s = 287;
	{8'd199,8'd229} : s = 122;
	{8'd199,8'd230} : s = 252;
	{8'd199,8'd231} : s = 250;
	{8'd199,8'd232} : s = 445;
	{8'd199,8'd233} : s = 43;
	{8'd199,8'd234} : s = 121;
	{8'd199,8'd235} : s = 118;
	{8'd199,8'd236} : s = 249;
	{8'd199,8'd237} : s = 117;
	{8'd199,8'd238} : s = 246;
	{8'd199,8'd239} : s = 245;
	{8'd199,8'd240} : s = 443;
	{8'd199,8'd241} : s = 115;
	{8'd199,8'd242} : s = 243;
	{8'd199,8'd243} : s = 238;
	{8'd199,8'd244} : s = 439;
	{8'd199,8'd245} : s = 237;
	{8'd199,8'd246} : s = 431;
	{8'd199,8'd247} : s = 415;
	{8'd199,8'd248} : s = 507;
	{8'd199,8'd249} : s = 7;
	{8'd199,8'd250} : s = 39;
	{8'd199,8'd251} : s = 30;
	{8'd199,8'd252} : s = 110;
	{8'd199,8'd253} : s = 29;
	{8'd199,8'd254} : s = 109;
	{8'd199,8'd255} : s = 107;
	{8'd200,8'd0} : s = 97;
	{8'd200,8'd1} : s = 228;
	{8'd200,8'd2} : s = 226;
	{8'd200,8'd3} : s = 370;
	{8'd200,8'd4} : s = 225;
	{8'd200,8'd5} : s = 369;
	{8'd200,8'd6} : s = 364;
	{8'd200,8'd7} : s = 470;
	{8'd200,8'd8} : s = 88;
	{8'd200,8'd9} : s = 216;
	{8'd200,8'd10} : s = 212;
	{8'd200,8'd11} : s = 362;
	{8'd200,8'd12} : s = 210;
	{8'd200,8'd13} : s = 361;
	{8'd200,8'd14} : s = 358;
	{8'd200,8'd15} : s = 469;
	{8'd200,8'd16} : s = 209;
	{8'd200,8'd17} : s = 357;
	{8'd200,8'd18} : s = 355;
	{8'd200,8'd19} : s = 467;
	{8'd200,8'd20} : s = 348;
	{8'd200,8'd21} : s = 462;
	{8'd200,8'd22} : s = 461;
	{8'd200,8'd23} : s = 505;
	{8'd200,8'd24} : s = 84;
	{8'd200,8'd25} : s = 204;
	{8'd200,8'd26} : s = 202;
	{8'd200,8'd27} : s = 346;
	{8'd200,8'd28} : s = 201;
	{8'd200,8'd29} : s = 345;
	{8'd200,8'd30} : s = 342;
	{8'd200,8'd31} : s = 459;
	{8'd200,8'd32} : s = 198;
	{8'd200,8'd33} : s = 341;
	{8'd200,8'd34} : s = 339;
	{8'd200,8'd35} : s = 455;
	{8'd200,8'd36} : s = 334;
	{8'd200,8'd37} : s = 444;
	{8'd200,8'd38} : s = 442;
	{8'd200,8'd39} : s = 502;
	{8'd200,8'd40} : s = 197;
	{8'd200,8'd41} : s = 333;
	{8'd200,8'd42} : s = 331;
	{8'd200,8'd43} : s = 441;
	{8'd200,8'd44} : s = 327;
	{8'd200,8'd45} : s = 438;
	{8'd200,8'd46} : s = 437;
	{8'd200,8'd47} : s = 501;
	{8'd200,8'd48} : s = 316;
	{8'd200,8'd49} : s = 435;
	{8'd200,8'd50} : s = 430;
	{8'd200,8'd51} : s = 499;
	{8'd200,8'd52} : s = 429;
	{8'd200,8'd53} : s = 494;
	{8'd200,8'd54} : s = 493;
	{8'd200,8'd55} : s = 510;
	{8'd200,8'd56} : s = 1;
	{8'd200,8'd57} : s = 18;
	{8'd200,8'd58} : s = 17;
	{8'd200,8'd59} : s = 82;
	{8'd200,8'd60} : s = 12;
	{8'd200,8'd61} : s = 81;
	{8'd200,8'd62} : s = 76;
	{8'd200,8'd63} : s = 195;
	{8'd200,8'd64} : s = 10;
	{8'd200,8'd65} : s = 74;
	{8'd200,8'd66} : s = 73;
	{8'd200,8'd67} : s = 184;
	{8'd200,8'd68} : s = 70;
	{8'd200,8'd69} : s = 180;
	{8'd200,8'd70} : s = 178;
	{8'd200,8'd71} : s = 314;
	{8'd200,8'd72} : s = 9;
	{8'd200,8'd73} : s = 69;
	{8'd200,8'd74} : s = 67;
	{8'd200,8'd75} : s = 177;
	{8'd200,8'd76} : s = 56;
	{8'd200,8'd77} : s = 172;
	{8'd200,8'd78} : s = 170;
	{8'd200,8'd79} : s = 313;
	{8'd200,8'd80} : s = 52;
	{8'd200,8'd81} : s = 169;
	{8'd200,8'd82} : s = 166;
	{8'd200,8'd83} : s = 310;
	{8'd200,8'd84} : s = 165;
	{8'd200,8'd85} : s = 309;
	{8'd200,8'd86} : s = 307;
	{8'd200,8'd87} : s = 427;
	{8'd200,8'd88} : s = 6;
	{8'd200,8'd89} : s = 50;
	{8'd200,8'd90} : s = 49;
	{8'd200,8'd91} : s = 163;
	{8'd200,8'd92} : s = 44;
	{8'd200,8'd93} : s = 156;
	{8'd200,8'd94} : s = 154;
	{8'd200,8'd95} : s = 302;
	{8'd200,8'd96} : s = 42;
	{8'd200,8'd97} : s = 153;
	{8'd200,8'd98} : s = 150;
	{8'd200,8'd99} : s = 301;
	{8'd200,8'd100} : s = 149;
	{8'd200,8'd101} : s = 299;
	{8'd200,8'd102} : s = 295;
	{8'd200,8'd103} : s = 423;
	{8'd200,8'd104} : s = 41;
	{8'd200,8'd105} : s = 147;
	{8'd200,8'd106} : s = 142;
	{8'd200,8'd107} : s = 286;
	{8'd200,8'd108} : s = 141;
	{8'd200,8'd109} : s = 285;
	{8'd200,8'd110} : s = 283;
	{8'd200,8'd111} : s = 414;
	{8'd200,8'd112} : s = 139;
	{8'd200,8'd113} : s = 279;
	{8'd200,8'd114} : s = 271;
	{8'd200,8'd115} : s = 413;
	{8'd200,8'd116} : s = 248;
	{8'd200,8'd117} : s = 411;
	{8'd200,8'd118} : s = 407;
	{8'd200,8'd119} : s = 491;
	{8'd200,8'd120} : s = 5;
	{8'd200,8'd121} : s = 38;
	{8'd200,8'd122} : s = 37;
	{8'd200,8'd123} : s = 135;
	{8'd200,8'd124} : s = 35;
	{8'd200,8'd125} : s = 120;
	{8'd200,8'd126} : s = 116;
	{8'd200,8'd127} : s = 244;
	{8'd200,8'd128} : s = 28;
	{8'd200,8'd129} : s = 114;
	{8'd200,8'd130} : s = 113;
	{8'd200,8'd131} : s = 242;
	{8'd200,8'd132} : s = 108;
	{8'd200,8'd133} : s = 241;
	{8'd200,8'd134} : s = 236;
	{8'd200,8'd135} : s = 399;
	{8'd200,8'd136} : s = 26;
	{8'd200,8'd137} : s = 106;
	{8'd200,8'd138} : s = 105;
	{8'd200,8'd139} : s = 234;
	{8'd200,8'd140} : s = 102;
	{8'd200,8'd141} : s = 233;
	{8'd200,8'd142} : s = 230;
	{8'd200,8'd143} : s = 380;
	{8'd200,8'd144} : s = 101;
	{8'd200,8'd145} : s = 229;
	{8'd200,8'd146} : s = 227;
	{8'd200,8'd147} : s = 378;
	{8'd200,8'd148} : s = 220;
	{8'd200,8'd149} : s = 377;
	{8'd200,8'd150} : s = 374;
	{8'd200,8'd151} : s = 487;
	{8'd200,8'd152} : s = 25;
	{8'd200,8'd153} : s = 99;
	{8'd200,8'd154} : s = 92;
	{8'd200,8'd155} : s = 218;
	{8'd200,8'd156} : s = 90;
	{8'd200,8'd157} : s = 217;
	{8'd200,8'd158} : s = 214;
	{8'd200,8'd159} : s = 373;
	{8'd200,8'd160} : s = 89;
	{8'd200,8'd161} : s = 213;
	{8'd200,8'd162} : s = 211;
	{8'd200,8'd163} : s = 371;
	{8'd200,8'd164} : s = 206;
	{8'd200,8'd165} : s = 366;
	{8'd200,8'd166} : s = 365;
	{8'd200,8'd167} : s = 478;
	{8'd200,8'd168} : s = 86;
	{8'd200,8'd169} : s = 205;
	{8'd200,8'd170} : s = 203;
	{8'd200,8'd171} : s = 363;
	{8'd200,8'd172} : s = 199;
	{8'd200,8'd173} : s = 359;
	{8'd200,8'd174} : s = 350;
	{8'd200,8'd175} : s = 477;
	{8'd200,8'd176} : s = 188;
	{8'd200,8'd177} : s = 349;
	{8'd200,8'd178} : s = 347;
	{8'd200,8'd179} : s = 475;
	{8'd200,8'd180} : s = 343;
	{8'd200,8'd181} : s = 471;
	{8'd200,8'd182} : s = 463;
	{8'd200,8'd183} : s = 509;
	{8'd200,8'd184} : s = 3;
	{8'd200,8'd185} : s = 22;
	{8'd200,8'd186} : s = 21;
	{8'd200,8'd187} : s = 85;
	{8'd200,8'd188} : s = 19;
	{8'd200,8'd189} : s = 83;
	{8'd200,8'd190} : s = 78;
	{8'd200,8'd191} : s = 186;
	{8'd200,8'd192} : s = 14;
	{8'd200,8'd193} : s = 77;
	{8'd200,8'd194} : s = 75;
	{8'd200,8'd195} : s = 185;
	{8'd200,8'd196} : s = 71;
	{8'd200,8'd197} : s = 182;
	{8'd200,8'd198} : s = 181;
	{8'd200,8'd199} : s = 335;
	{8'd200,8'd200} : s = 13;
	{8'd200,8'd201} : s = 60;
	{8'd200,8'd202} : s = 58;
	{8'd200,8'd203} : s = 179;
	{8'd200,8'd204} : s = 57;
	{8'd200,8'd205} : s = 174;
	{8'd200,8'd206} : s = 173;
	{8'd200,8'd207} : s = 318;
	{8'd200,8'd208} : s = 54;
	{8'd200,8'd209} : s = 171;
	{8'd200,8'd210} : s = 167;
	{8'd200,8'd211} : s = 317;
	{8'd200,8'd212} : s = 158;
	{8'd200,8'd213} : s = 315;
	{8'd200,8'd214} : s = 311;
	{8'd200,8'd215} : s = 446;
	{8'd200,8'd216} : s = 11;
	{8'd200,8'd217} : s = 53;
	{8'd200,8'd218} : s = 51;
	{8'd200,8'd219} : s = 157;
	{8'd200,8'd220} : s = 46;
	{8'd200,8'd221} : s = 155;
	{8'd200,8'd222} : s = 151;
	{8'd200,8'd223} : s = 303;
	{8'd200,8'd224} : s = 45;
	{8'd200,8'd225} : s = 143;
	{8'd200,8'd226} : s = 124;
	{8'd200,8'd227} : s = 287;
	{8'd200,8'd228} : s = 122;
	{8'd200,8'd229} : s = 252;
	{8'd200,8'd230} : s = 250;
	{8'd200,8'd231} : s = 445;
	{8'd200,8'd232} : s = 43;
	{8'd200,8'd233} : s = 121;
	{8'd200,8'd234} : s = 118;
	{8'd200,8'd235} : s = 249;
	{8'd200,8'd236} : s = 117;
	{8'd200,8'd237} : s = 246;
	{8'd200,8'd238} : s = 245;
	{8'd200,8'd239} : s = 443;
	{8'd200,8'd240} : s = 115;
	{8'd200,8'd241} : s = 243;
	{8'd200,8'd242} : s = 238;
	{8'd200,8'd243} : s = 439;
	{8'd200,8'd244} : s = 237;
	{8'd200,8'd245} : s = 431;
	{8'd200,8'd246} : s = 415;
	{8'd200,8'd247} : s = 507;
	{8'd200,8'd248} : s = 7;
	{8'd200,8'd249} : s = 39;
	{8'd200,8'd250} : s = 30;
	{8'd200,8'd251} : s = 110;
	{8'd200,8'd252} : s = 29;
	{8'd200,8'd253} : s = 109;
	{8'd200,8'd254} : s = 107;
	{8'd200,8'd255} : s = 235;
	{8'd201,8'd0} : s = 228;
	{8'd201,8'd1} : s = 226;
	{8'd201,8'd2} : s = 370;
	{8'd201,8'd3} : s = 225;
	{8'd201,8'd4} : s = 369;
	{8'd201,8'd5} : s = 364;
	{8'd201,8'd6} : s = 470;
	{8'd201,8'd7} : s = 88;
	{8'd201,8'd8} : s = 216;
	{8'd201,8'd9} : s = 212;
	{8'd201,8'd10} : s = 362;
	{8'd201,8'd11} : s = 210;
	{8'd201,8'd12} : s = 361;
	{8'd201,8'd13} : s = 358;
	{8'd201,8'd14} : s = 469;
	{8'd201,8'd15} : s = 209;
	{8'd201,8'd16} : s = 357;
	{8'd201,8'd17} : s = 355;
	{8'd201,8'd18} : s = 467;
	{8'd201,8'd19} : s = 348;
	{8'd201,8'd20} : s = 462;
	{8'd201,8'd21} : s = 461;
	{8'd201,8'd22} : s = 505;
	{8'd201,8'd23} : s = 84;
	{8'd201,8'd24} : s = 204;
	{8'd201,8'd25} : s = 202;
	{8'd201,8'd26} : s = 346;
	{8'd201,8'd27} : s = 201;
	{8'd201,8'd28} : s = 345;
	{8'd201,8'd29} : s = 342;
	{8'd201,8'd30} : s = 459;
	{8'd201,8'd31} : s = 198;
	{8'd201,8'd32} : s = 341;
	{8'd201,8'd33} : s = 339;
	{8'd201,8'd34} : s = 455;
	{8'd201,8'd35} : s = 334;
	{8'd201,8'd36} : s = 444;
	{8'd201,8'd37} : s = 442;
	{8'd201,8'd38} : s = 502;
	{8'd201,8'd39} : s = 197;
	{8'd201,8'd40} : s = 333;
	{8'd201,8'd41} : s = 331;
	{8'd201,8'd42} : s = 441;
	{8'd201,8'd43} : s = 327;
	{8'd201,8'd44} : s = 438;
	{8'd201,8'd45} : s = 437;
	{8'd201,8'd46} : s = 501;
	{8'd201,8'd47} : s = 316;
	{8'd201,8'd48} : s = 435;
	{8'd201,8'd49} : s = 430;
	{8'd201,8'd50} : s = 499;
	{8'd201,8'd51} : s = 429;
	{8'd201,8'd52} : s = 494;
	{8'd201,8'd53} : s = 493;
	{8'd201,8'd54} : s = 510;
	{8'd201,8'd55} : s = 1;
	{8'd201,8'd56} : s = 18;
	{8'd201,8'd57} : s = 17;
	{8'd201,8'd58} : s = 82;
	{8'd201,8'd59} : s = 12;
	{8'd201,8'd60} : s = 81;
	{8'd201,8'd61} : s = 76;
	{8'd201,8'd62} : s = 195;
	{8'd201,8'd63} : s = 10;
	{8'd201,8'd64} : s = 74;
	{8'd201,8'd65} : s = 73;
	{8'd201,8'd66} : s = 184;
	{8'd201,8'd67} : s = 70;
	{8'd201,8'd68} : s = 180;
	{8'd201,8'd69} : s = 178;
	{8'd201,8'd70} : s = 314;
	{8'd201,8'd71} : s = 9;
	{8'd201,8'd72} : s = 69;
	{8'd201,8'd73} : s = 67;
	{8'd201,8'd74} : s = 177;
	{8'd201,8'd75} : s = 56;
	{8'd201,8'd76} : s = 172;
	{8'd201,8'd77} : s = 170;
	{8'd201,8'd78} : s = 313;
	{8'd201,8'd79} : s = 52;
	{8'd201,8'd80} : s = 169;
	{8'd201,8'd81} : s = 166;
	{8'd201,8'd82} : s = 310;
	{8'd201,8'd83} : s = 165;
	{8'd201,8'd84} : s = 309;
	{8'd201,8'd85} : s = 307;
	{8'd201,8'd86} : s = 427;
	{8'd201,8'd87} : s = 6;
	{8'd201,8'd88} : s = 50;
	{8'd201,8'd89} : s = 49;
	{8'd201,8'd90} : s = 163;
	{8'd201,8'd91} : s = 44;
	{8'd201,8'd92} : s = 156;
	{8'd201,8'd93} : s = 154;
	{8'd201,8'd94} : s = 302;
	{8'd201,8'd95} : s = 42;
	{8'd201,8'd96} : s = 153;
	{8'd201,8'd97} : s = 150;
	{8'd201,8'd98} : s = 301;
	{8'd201,8'd99} : s = 149;
	{8'd201,8'd100} : s = 299;
	{8'd201,8'd101} : s = 295;
	{8'd201,8'd102} : s = 423;
	{8'd201,8'd103} : s = 41;
	{8'd201,8'd104} : s = 147;
	{8'd201,8'd105} : s = 142;
	{8'd201,8'd106} : s = 286;
	{8'd201,8'd107} : s = 141;
	{8'd201,8'd108} : s = 285;
	{8'd201,8'd109} : s = 283;
	{8'd201,8'd110} : s = 414;
	{8'd201,8'd111} : s = 139;
	{8'd201,8'd112} : s = 279;
	{8'd201,8'd113} : s = 271;
	{8'd201,8'd114} : s = 413;
	{8'd201,8'd115} : s = 248;
	{8'd201,8'd116} : s = 411;
	{8'd201,8'd117} : s = 407;
	{8'd201,8'd118} : s = 491;
	{8'd201,8'd119} : s = 5;
	{8'd201,8'd120} : s = 38;
	{8'd201,8'd121} : s = 37;
	{8'd201,8'd122} : s = 135;
	{8'd201,8'd123} : s = 35;
	{8'd201,8'd124} : s = 120;
	{8'd201,8'd125} : s = 116;
	{8'd201,8'd126} : s = 244;
	{8'd201,8'd127} : s = 28;
	{8'd201,8'd128} : s = 114;
	{8'd201,8'd129} : s = 113;
	{8'd201,8'd130} : s = 242;
	{8'd201,8'd131} : s = 108;
	{8'd201,8'd132} : s = 241;
	{8'd201,8'd133} : s = 236;
	{8'd201,8'd134} : s = 399;
	{8'd201,8'd135} : s = 26;
	{8'd201,8'd136} : s = 106;
	{8'd201,8'd137} : s = 105;
	{8'd201,8'd138} : s = 234;
	{8'd201,8'd139} : s = 102;
	{8'd201,8'd140} : s = 233;
	{8'd201,8'd141} : s = 230;
	{8'd201,8'd142} : s = 380;
	{8'd201,8'd143} : s = 101;
	{8'd201,8'd144} : s = 229;
	{8'd201,8'd145} : s = 227;
	{8'd201,8'd146} : s = 378;
	{8'd201,8'd147} : s = 220;
	{8'd201,8'd148} : s = 377;
	{8'd201,8'd149} : s = 374;
	{8'd201,8'd150} : s = 487;
	{8'd201,8'd151} : s = 25;
	{8'd201,8'd152} : s = 99;
	{8'd201,8'd153} : s = 92;
	{8'd201,8'd154} : s = 218;
	{8'd201,8'd155} : s = 90;
	{8'd201,8'd156} : s = 217;
	{8'd201,8'd157} : s = 214;
	{8'd201,8'd158} : s = 373;
	{8'd201,8'd159} : s = 89;
	{8'd201,8'd160} : s = 213;
	{8'd201,8'd161} : s = 211;
	{8'd201,8'd162} : s = 371;
	{8'd201,8'd163} : s = 206;
	{8'd201,8'd164} : s = 366;
	{8'd201,8'd165} : s = 365;
	{8'd201,8'd166} : s = 478;
	{8'd201,8'd167} : s = 86;
	{8'd201,8'd168} : s = 205;
	{8'd201,8'd169} : s = 203;
	{8'd201,8'd170} : s = 363;
	{8'd201,8'd171} : s = 199;
	{8'd201,8'd172} : s = 359;
	{8'd201,8'd173} : s = 350;
	{8'd201,8'd174} : s = 477;
	{8'd201,8'd175} : s = 188;
	{8'd201,8'd176} : s = 349;
	{8'd201,8'd177} : s = 347;
	{8'd201,8'd178} : s = 475;
	{8'd201,8'd179} : s = 343;
	{8'd201,8'd180} : s = 471;
	{8'd201,8'd181} : s = 463;
	{8'd201,8'd182} : s = 509;
	{8'd201,8'd183} : s = 3;
	{8'd201,8'd184} : s = 22;
	{8'd201,8'd185} : s = 21;
	{8'd201,8'd186} : s = 85;
	{8'd201,8'd187} : s = 19;
	{8'd201,8'd188} : s = 83;
	{8'd201,8'd189} : s = 78;
	{8'd201,8'd190} : s = 186;
	{8'd201,8'd191} : s = 14;
	{8'd201,8'd192} : s = 77;
	{8'd201,8'd193} : s = 75;
	{8'd201,8'd194} : s = 185;
	{8'd201,8'd195} : s = 71;
	{8'd201,8'd196} : s = 182;
	{8'd201,8'd197} : s = 181;
	{8'd201,8'd198} : s = 335;
	{8'd201,8'd199} : s = 13;
	{8'd201,8'd200} : s = 60;
	{8'd201,8'd201} : s = 58;
	{8'd201,8'd202} : s = 179;
	{8'd201,8'd203} : s = 57;
	{8'd201,8'd204} : s = 174;
	{8'd201,8'd205} : s = 173;
	{8'd201,8'd206} : s = 318;
	{8'd201,8'd207} : s = 54;
	{8'd201,8'd208} : s = 171;
	{8'd201,8'd209} : s = 167;
	{8'd201,8'd210} : s = 317;
	{8'd201,8'd211} : s = 158;
	{8'd201,8'd212} : s = 315;
	{8'd201,8'd213} : s = 311;
	{8'd201,8'd214} : s = 446;
	{8'd201,8'd215} : s = 11;
	{8'd201,8'd216} : s = 53;
	{8'd201,8'd217} : s = 51;
	{8'd201,8'd218} : s = 157;
	{8'd201,8'd219} : s = 46;
	{8'd201,8'd220} : s = 155;
	{8'd201,8'd221} : s = 151;
	{8'd201,8'd222} : s = 303;
	{8'd201,8'd223} : s = 45;
	{8'd201,8'd224} : s = 143;
	{8'd201,8'd225} : s = 124;
	{8'd201,8'd226} : s = 287;
	{8'd201,8'd227} : s = 122;
	{8'd201,8'd228} : s = 252;
	{8'd201,8'd229} : s = 250;
	{8'd201,8'd230} : s = 445;
	{8'd201,8'd231} : s = 43;
	{8'd201,8'd232} : s = 121;
	{8'd201,8'd233} : s = 118;
	{8'd201,8'd234} : s = 249;
	{8'd201,8'd235} : s = 117;
	{8'd201,8'd236} : s = 246;
	{8'd201,8'd237} : s = 245;
	{8'd201,8'd238} : s = 443;
	{8'd201,8'd239} : s = 115;
	{8'd201,8'd240} : s = 243;
	{8'd201,8'd241} : s = 238;
	{8'd201,8'd242} : s = 439;
	{8'd201,8'd243} : s = 237;
	{8'd201,8'd244} : s = 431;
	{8'd201,8'd245} : s = 415;
	{8'd201,8'd246} : s = 507;
	{8'd201,8'd247} : s = 7;
	{8'd201,8'd248} : s = 39;
	{8'd201,8'd249} : s = 30;
	{8'd201,8'd250} : s = 110;
	{8'd201,8'd251} : s = 29;
	{8'd201,8'd252} : s = 109;
	{8'd201,8'd253} : s = 107;
	{8'd201,8'd254} : s = 235;
	{8'd201,8'd255} : s = 27;
	{8'd202,8'd0} : s = 226;
	{8'd202,8'd1} : s = 370;
	{8'd202,8'd2} : s = 225;
	{8'd202,8'd3} : s = 369;
	{8'd202,8'd4} : s = 364;
	{8'd202,8'd5} : s = 470;
	{8'd202,8'd6} : s = 88;
	{8'd202,8'd7} : s = 216;
	{8'd202,8'd8} : s = 212;
	{8'd202,8'd9} : s = 362;
	{8'd202,8'd10} : s = 210;
	{8'd202,8'd11} : s = 361;
	{8'd202,8'd12} : s = 358;
	{8'd202,8'd13} : s = 469;
	{8'd202,8'd14} : s = 209;
	{8'd202,8'd15} : s = 357;
	{8'd202,8'd16} : s = 355;
	{8'd202,8'd17} : s = 467;
	{8'd202,8'd18} : s = 348;
	{8'd202,8'd19} : s = 462;
	{8'd202,8'd20} : s = 461;
	{8'd202,8'd21} : s = 505;
	{8'd202,8'd22} : s = 84;
	{8'd202,8'd23} : s = 204;
	{8'd202,8'd24} : s = 202;
	{8'd202,8'd25} : s = 346;
	{8'd202,8'd26} : s = 201;
	{8'd202,8'd27} : s = 345;
	{8'd202,8'd28} : s = 342;
	{8'd202,8'd29} : s = 459;
	{8'd202,8'd30} : s = 198;
	{8'd202,8'd31} : s = 341;
	{8'd202,8'd32} : s = 339;
	{8'd202,8'd33} : s = 455;
	{8'd202,8'd34} : s = 334;
	{8'd202,8'd35} : s = 444;
	{8'd202,8'd36} : s = 442;
	{8'd202,8'd37} : s = 502;
	{8'd202,8'd38} : s = 197;
	{8'd202,8'd39} : s = 333;
	{8'd202,8'd40} : s = 331;
	{8'd202,8'd41} : s = 441;
	{8'd202,8'd42} : s = 327;
	{8'd202,8'd43} : s = 438;
	{8'd202,8'd44} : s = 437;
	{8'd202,8'd45} : s = 501;
	{8'd202,8'd46} : s = 316;
	{8'd202,8'd47} : s = 435;
	{8'd202,8'd48} : s = 430;
	{8'd202,8'd49} : s = 499;
	{8'd202,8'd50} : s = 429;
	{8'd202,8'd51} : s = 494;
	{8'd202,8'd52} : s = 493;
	{8'd202,8'd53} : s = 510;
	{8'd202,8'd54} : s = 1;
	{8'd202,8'd55} : s = 18;
	{8'd202,8'd56} : s = 17;
	{8'd202,8'd57} : s = 82;
	{8'd202,8'd58} : s = 12;
	{8'd202,8'd59} : s = 81;
	{8'd202,8'd60} : s = 76;
	{8'd202,8'd61} : s = 195;
	{8'd202,8'd62} : s = 10;
	{8'd202,8'd63} : s = 74;
	{8'd202,8'd64} : s = 73;
	{8'd202,8'd65} : s = 184;
	{8'd202,8'd66} : s = 70;
	{8'd202,8'd67} : s = 180;
	{8'd202,8'd68} : s = 178;
	{8'd202,8'd69} : s = 314;
	{8'd202,8'd70} : s = 9;
	{8'd202,8'd71} : s = 69;
	{8'd202,8'd72} : s = 67;
	{8'd202,8'd73} : s = 177;
	{8'd202,8'd74} : s = 56;
	{8'd202,8'd75} : s = 172;
	{8'd202,8'd76} : s = 170;
	{8'd202,8'd77} : s = 313;
	{8'd202,8'd78} : s = 52;
	{8'd202,8'd79} : s = 169;
	{8'd202,8'd80} : s = 166;
	{8'd202,8'd81} : s = 310;
	{8'd202,8'd82} : s = 165;
	{8'd202,8'd83} : s = 309;
	{8'd202,8'd84} : s = 307;
	{8'd202,8'd85} : s = 427;
	{8'd202,8'd86} : s = 6;
	{8'd202,8'd87} : s = 50;
	{8'd202,8'd88} : s = 49;
	{8'd202,8'd89} : s = 163;
	{8'd202,8'd90} : s = 44;
	{8'd202,8'd91} : s = 156;
	{8'd202,8'd92} : s = 154;
	{8'd202,8'd93} : s = 302;
	{8'd202,8'd94} : s = 42;
	{8'd202,8'd95} : s = 153;
	{8'd202,8'd96} : s = 150;
	{8'd202,8'd97} : s = 301;
	{8'd202,8'd98} : s = 149;
	{8'd202,8'd99} : s = 299;
	{8'd202,8'd100} : s = 295;
	{8'd202,8'd101} : s = 423;
	{8'd202,8'd102} : s = 41;
	{8'd202,8'd103} : s = 147;
	{8'd202,8'd104} : s = 142;
	{8'd202,8'd105} : s = 286;
	{8'd202,8'd106} : s = 141;
	{8'd202,8'd107} : s = 285;
	{8'd202,8'd108} : s = 283;
	{8'd202,8'd109} : s = 414;
	{8'd202,8'd110} : s = 139;
	{8'd202,8'd111} : s = 279;
	{8'd202,8'd112} : s = 271;
	{8'd202,8'd113} : s = 413;
	{8'd202,8'd114} : s = 248;
	{8'd202,8'd115} : s = 411;
	{8'd202,8'd116} : s = 407;
	{8'd202,8'd117} : s = 491;
	{8'd202,8'd118} : s = 5;
	{8'd202,8'd119} : s = 38;
	{8'd202,8'd120} : s = 37;
	{8'd202,8'd121} : s = 135;
	{8'd202,8'd122} : s = 35;
	{8'd202,8'd123} : s = 120;
	{8'd202,8'd124} : s = 116;
	{8'd202,8'd125} : s = 244;
	{8'd202,8'd126} : s = 28;
	{8'd202,8'd127} : s = 114;
	{8'd202,8'd128} : s = 113;
	{8'd202,8'd129} : s = 242;
	{8'd202,8'd130} : s = 108;
	{8'd202,8'd131} : s = 241;
	{8'd202,8'd132} : s = 236;
	{8'd202,8'd133} : s = 399;
	{8'd202,8'd134} : s = 26;
	{8'd202,8'd135} : s = 106;
	{8'd202,8'd136} : s = 105;
	{8'd202,8'd137} : s = 234;
	{8'd202,8'd138} : s = 102;
	{8'd202,8'd139} : s = 233;
	{8'd202,8'd140} : s = 230;
	{8'd202,8'd141} : s = 380;
	{8'd202,8'd142} : s = 101;
	{8'd202,8'd143} : s = 229;
	{8'd202,8'd144} : s = 227;
	{8'd202,8'd145} : s = 378;
	{8'd202,8'd146} : s = 220;
	{8'd202,8'd147} : s = 377;
	{8'd202,8'd148} : s = 374;
	{8'd202,8'd149} : s = 487;
	{8'd202,8'd150} : s = 25;
	{8'd202,8'd151} : s = 99;
	{8'd202,8'd152} : s = 92;
	{8'd202,8'd153} : s = 218;
	{8'd202,8'd154} : s = 90;
	{8'd202,8'd155} : s = 217;
	{8'd202,8'd156} : s = 214;
	{8'd202,8'd157} : s = 373;
	{8'd202,8'd158} : s = 89;
	{8'd202,8'd159} : s = 213;
	{8'd202,8'd160} : s = 211;
	{8'd202,8'd161} : s = 371;
	{8'd202,8'd162} : s = 206;
	{8'd202,8'd163} : s = 366;
	{8'd202,8'd164} : s = 365;
	{8'd202,8'd165} : s = 478;
	{8'd202,8'd166} : s = 86;
	{8'd202,8'd167} : s = 205;
	{8'd202,8'd168} : s = 203;
	{8'd202,8'd169} : s = 363;
	{8'd202,8'd170} : s = 199;
	{8'd202,8'd171} : s = 359;
	{8'd202,8'd172} : s = 350;
	{8'd202,8'd173} : s = 477;
	{8'd202,8'd174} : s = 188;
	{8'd202,8'd175} : s = 349;
	{8'd202,8'd176} : s = 347;
	{8'd202,8'd177} : s = 475;
	{8'd202,8'd178} : s = 343;
	{8'd202,8'd179} : s = 471;
	{8'd202,8'd180} : s = 463;
	{8'd202,8'd181} : s = 509;
	{8'd202,8'd182} : s = 3;
	{8'd202,8'd183} : s = 22;
	{8'd202,8'd184} : s = 21;
	{8'd202,8'd185} : s = 85;
	{8'd202,8'd186} : s = 19;
	{8'd202,8'd187} : s = 83;
	{8'd202,8'd188} : s = 78;
	{8'd202,8'd189} : s = 186;
	{8'd202,8'd190} : s = 14;
	{8'd202,8'd191} : s = 77;
	{8'd202,8'd192} : s = 75;
	{8'd202,8'd193} : s = 185;
	{8'd202,8'd194} : s = 71;
	{8'd202,8'd195} : s = 182;
	{8'd202,8'd196} : s = 181;
	{8'd202,8'd197} : s = 335;
	{8'd202,8'd198} : s = 13;
	{8'd202,8'd199} : s = 60;
	{8'd202,8'd200} : s = 58;
	{8'd202,8'd201} : s = 179;
	{8'd202,8'd202} : s = 57;
	{8'd202,8'd203} : s = 174;
	{8'd202,8'd204} : s = 173;
	{8'd202,8'd205} : s = 318;
	{8'd202,8'd206} : s = 54;
	{8'd202,8'd207} : s = 171;
	{8'd202,8'd208} : s = 167;
	{8'd202,8'd209} : s = 317;
	{8'd202,8'd210} : s = 158;
	{8'd202,8'd211} : s = 315;
	{8'd202,8'd212} : s = 311;
	{8'd202,8'd213} : s = 446;
	{8'd202,8'd214} : s = 11;
	{8'd202,8'd215} : s = 53;
	{8'd202,8'd216} : s = 51;
	{8'd202,8'd217} : s = 157;
	{8'd202,8'd218} : s = 46;
	{8'd202,8'd219} : s = 155;
	{8'd202,8'd220} : s = 151;
	{8'd202,8'd221} : s = 303;
	{8'd202,8'd222} : s = 45;
	{8'd202,8'd223} : s = 143;
	{8'd202,8'd224} : s = 124;
	{8'd202,8'd225} : s = 287;
	{8'd202,8'd226} : s = 122;
	{8'd202,8'd227} : s = 252;
	{8'd202,8'd228} : s = 250;
	{8'd202,8'd229} : s = 445;
	{8'd202,8'd230} : s = 43;
	{8'd202,8'd231} : s = 121;
	{8'd202,8'd232} : s = 118;
	{8'd202,8'd233} : s = 249;
	{8'd202,8'd234} : s = 117;
	{8'd202,8'd235} : s = 246;
	{8'd202,8'd236} : s = 245;
	{8'd202,8'd237} : s = 443;
	{8'd202,8'd238} : s = 115;
	{8'd202,8'd239} : s = 243;
	{8'd202,8'd240} : s = 238;
	{8'd202,8'd241} : s = 439;
	{8'd202,8'd242} : s = 237;
	{8'd202,8'd243} : s = 431;
	{8'd202,8'd244} : s = 415;
	{8'd202,8'd245} : s = 507;
	{8'd202,8'd246} : s = 7;
	{8'd202,8'd247} : s = 39;
	{8'd202,8'd248} : s = 30;
	{8'd202,8'd249} : s = 110;
	{8'd202,8'd250} : s = 29;
	{8'd202,8'd251} : s = 109;
	{8'd202,8'd252} : s = 107;
	{8'd202,8'd253} : s = 235;
	{8'd202,8'd254} : s = 27;
	{8'd202,8'd255} : s = 103;
	{8'd203,8'd0} : s = 370;
	{8'd203,8'd1} : s = 225;
	{8'd203,8'd2} : s = 369;
	{8'd203,8'd3} : s = 364;
	{8'd203,8'd4} : s = 470;
	{8'd203,8'd5} : s = 88;
	{8'd203,8'd6} : s = 216;
	{8'd203,8'd7} : s = 212;
	{8'd203,8'd8} : s = 362;
	{8'd203,8'd9} : s = 210;
	{8'd203,8'd10} : s = 361;
	{8'd203,8'd11} : s = 358;
	{8'd203,8'd12} : s = 469;
	{8'd203,8'd13} : s = 209;
	{8'd203,8'd14} : s = 357;
	{8'd203,8'd15} : s = 355;
	{8'd203,8'd16} : s = 467;
	{8'd203,8'd17} : s = 348;
	{8'd203,8'd18} : s = 462;
	{8'd203,8'd19} : s = 461;
	{8'd203,8'd20} : s = 505;
	{8'd203,8'd21} : s = 84;
	{8'd203,8'd22} : s = 204;
	{8'd203,8'd23} : s = 202;
	{8'd203,8'd24} : s = 346;
	{8'd203,8'd25} : s = 201;
	{8'd203,8'd26} : s = 345;
	{8'd203,8'd27} : s = 342;
	{8'd203,8'd28} : s = 459;
	{8'd203,8'd29} : s = 198;
	{8'd203,8'd30} : s = 341;
	{8'd203,8'd31} : s = 339;
	{8'd203,8'd32} : s = 455;
	{8'd203,8'd33} : s = 334;
	{8'd203,8'd34} : s = 444;
	{8'd203,8'd35} : s = 442;
	{8'd203,8'd36} : s = 502;
	{8'd203,8'd37} : s = 197;
	{8'd203,8'd38} : s = 333;
	{8'd203,8'd39} : s = 331;
	{8'd203,8'd40} : s = 441;
	{8'd203,8'd41} : s = 327;
	{8'd203,8'd42} : s = 438;
	{8'd203,8'd43} : s = 437;
	{8'd203,8'd44} : s = 501;
	{8'd203,8'd45} : s = 316;
	{8'd203,8'd46} : s = 435;
	{8'd203,8'd47} : s = 430;
	{8'd203,8'd48} : s = 499;
	{8'd203,8'd49} : s = 429;
	{8'd203,8'd50} : s = 494;
	{8'd203,8'd51} : s = 493;
	{8'd203,8'd52} : s = 510;
	{8'd203,8'd53} : s = 1;
	{8'd203,8'd54} : s = 18;
	{8'd203,8'd55} : s = 17;
	{8'd203,8'd56} : s = 82;
	{8'd203,8'd57} : s = 12;
	{8'd203,8'd58} : s = 81;
	{8'd203,8'd59} : s = 76;
	{8'd203,8'd60} : s = 195;
	{8'd203,8'd61} : s = 10;
	{8'd203,8'd62} : s = 74;
	{8'd203,8'd63} : s = 73;
	{8'd203,8'd64} : s = 184;
	{8'd203,8'd65} : s = 70;
	{8'd203,8'd66} : s = 180;
	{8'd203,8'd67} : s = 178;
	{8'd203,8'd68} : s = 314;
	{8'd203,8'd69} : s = 9;
	{8'd203,8'd70} : s = 69;
	{8'd203,8'd71} : s = 67;
	{8'd203,8'd72} : s = 177;
	{8'd203,8'd73} : s = 56;
	{8'd203,8'd74} : s = 172;
	{8'd203,8'd75} : s = 170;
	{8'd203,8'd76} : s = 313;
	{8'd203,8'd77} : s = 52;
	{8'd203,8'd78} : s = 169;
	{8'd203,8'd79} : s = 166;
	{8'd203,8'd80} : s = 310;
	{8'd203,8'd81} : s = 165;
	{8'd203,8'd82} : s = 309;
	{8'd203,8'd83} : s = 307;
	{8'd203,8'd84} : s = 427;
	{8'd203,8'd85} : s = 6;
	{8'd203,8'd86} : s = 50;
	{8'd203,8'd87} : s = 49;
	{8'd203,8'd88} : s = 163;
	{8'd203,8'd89} : s = 44;
	{8'd203,8'd90} : s = 156;
	{8'd203,8'd91} : s = 154;
	{8'd203,8'd92} : s = 302;
	{8'd203,8'd93} : s = 42;
	{8'd203,8'd94} : s = 153;
	{8'd203,8'd95} : s = 150;
	{8'd203,8'd96} : s = 301;
	{8'd203,8'd97} : s = 149;
	{8'd203,8'd98} : s = 299;
	{8'd203,8'd99} : s = 295;
	{8'd203,8'd100} : s = 423;
	{8'd203,8'd101} : s = 41;
	{8'd203,8'd102} : s = 147;
	{8'd203,8'd103} : s = 142;
	{8'd203,8'd104} : s = 286;
	{8'd203,8'd105} : s = 141;
	{8'd203,8'd106} : s = 285;
	{8'd203,8'd107} : s = 283;
	{8'd203,8'd108} : s = 414;
	{8'd203,8'd109} : s = 139;
	{8'd203,8'd110} : s = 279;
	{8'd203,8'd111} : s = 271;
	{8'd203,8'd112} : s = 413;
	{8'd203,8'd113} : s = 248;
	{8'd203,8'd114} : s = 411;
	{8'd203,8'd115} : s = 407;
	{8'd203,8'd116} : s = 491;
	{8'd203,8'd117} : s = 5;
	{8'd203,8'd118} : s = 38;
	{8'd203,8'd119} : s = 37;
	{8'd203,8'd120} : s = 135;
	{8'd203,8'd121} : s = 35;
	{8'd203,8'd122} : s = 120;
	{8'd203,8'd123} : s = 116;
	{8'd203,8'd124} : s = 244;
	{8'd203,8'd125} : s = 28;
	{8'd203,8'd126} : s = 114;
	{8'd203,8'd127} : s = 113;
	{8'd203,8'd128} : s = 242;
	{8'd203,8'd129} : s = 108;
	{8'd203,8'd130} : s = 241;
	{8'd203,8'd131} : s = 236;
	{8'd203,8'd132} : s = 399;
	{8'd203,8'd133} : s = 26;
	{8'd203,8'd134} : s = 106;
	{8'd203,8'd135} : s = 105;
	{8'd203,8'd136} : s = 234;
	{8'd203,8'd137} : s = 102;
	{8'd203,8'd138} : s = 233;
	{8'd203,8'd139} : s = 230;
	{8'd203,8'd140} : s = 380;
	{8'd203,8'd141} : s = 101;
	{8'd203,8'd142} : s = 229;
	{8'd203,8'd143} : s = 227;
	{8'd203,8'd144} : s = 378;
	{8'd203,8'd145} : s = 220;
	{8'd203,8'd146} : s = 377;
	{8'd203,8'd147} : s = 374;
	{8'd203,8'd148} : s = 487;
	{8'd203,8'd149} : s = 25;
	{8'd203,8'd150} : s = 99;
	{8'd203,8'd151} : s = 92;
	{8'd203,8'd152} : s = 218;
	{8'd203,8'd153} : s = 90;
	{8'd203,8'd154} : s = 217;
	{8'd203,8'd155} : s = 214;
	{8'd203,8'd156} : s = 373;
	{8'd203,8'd157} : s = 89;
	{8'd203,8'd158} : s = 213;
	{8'd203,8'd159} : s = 211;
	{8'd203,8'd160} : s = 371;
	{8'd203,8'd161} : s = 206;
	{8'd203,8'd162} : s = 366;
	{8'd203,8'd163} : s = 365;
	{8'd203,8'd164} : s = 478;
	{8'd203,8'd165} : s = 86;
	{8'd203,8'd166} : s = 205;
	{8'd203,8'd167} : s = 203;
	{8'd203,8'd168} : s = 363;
	{8'd203,8'd169} : s = 199;
	{8'd203,8'd170} : s = 359;
	{8'd203,8'd171} : s = 350;
	{8'd203,8'd172} : s = 477;
	{8'd203,8'd173} : s = 188;
	{8'd203,8'd174} : s = 349;
	{8'd203,8'd175} : s = 347;
	{8'd203,8'd176} : s = 475;
	{8'd203,8'd177} : s = 343;
	{8'd203,8'd178} : s = 471;
	{8'd203,8'd179} : s = 463;
	{8'd203,8'd180} : s = 509;
	{8'd203,8'd181} : s = 3;
	{8'd203,8'd182} : s = 22;
	{8'd203,8'd183} : s = 21;
	{8'd203,8'd184} : s = 85;
	{8'd203,8'd185} : s = 19;
	{8'd203,8'd186} : s = 83;
	{8'd203,8'd187} : s = 78;
	{8'd203,8'd188} : s = 186;
	{8'd203,8'd189} : s = 14;
	{8'd203,8'd190} : s = 77;
	{8'd203,8'd191} : s = 75;
	{8'd203,8'd192} : s = 185;
	{8'd203,8'd193} : s = 71;
	{8'd203,8'd194} : s = 182;
	{8'd203,8'd195} : s = 181;
	{8'd203,8'd196} : s = 335;
	{8'd203,8'd197} : s = 13;
	{8'd203,8'd198} : s = 60;
	{8'd203,8'd199} : s = 58;
	{8'd203,8'd200} : s = 179;
	{8'd203,8'd201} : s = 57;
	{8'd203,8'd202} : s = 174;
	{8'd203,8'd203} : s = 173;
	{8'd203,8'd204} : s = 318;
	{8'd203,8'd205} : s = 54;
	{8'd203,8'd206} : s = 171;
	{8'd203,8'd207} : s = 167;
	{8'd203,8'd208} : s = 317;
	{8'd203,8'd209} : s = 158;
	{8'd203,8'd210} : s = 315;
	{8'd203,8'd211} : s = 311;
	{8'd203,8'd212} : s = 446;
	{8'd203,8'd213} : s = 11;
	{8'd203,8'd214} : s = 53;
	{8'd203,8'd215} : s = 51;
	{8'd203,8'd216} : s = 157;
	{8'd203,8'd217} : s = 46;
	{8'd203,8'd218} : s = 155;
	{8'd203,8'd219} : s = 151;
	{8'd203,8'd220} : s = 303;
	{8'd203,8'd221} : s = 45;
	{8'd203,8'd222} : s = 143;
	{8'd203,8'd223} : s = 124;
	{8'd203,8'd224} : s = 287;
	{8'd203,8'd225} : s = 122;
	{8'd203,8'd226} : s = 252;
	{8'd203,8'd227} : s = 250;
	{8'd203,8'd228} : s = 445;
	{8'd203,8'd229} : s = 43;
	{8'd203,8'd230} : s = 121;
	{8'd203,8'd231} : s = 118;
	{8'd203,8'd232} : s = 249;
	{8'd203,8'd233} : s = 117;
	{8'd203,8'd234} : s = 246;
	{8'd203,8'd235} : s = 245;
	{8'd203,8'd236} : s = 443;
	{8'd203,8'd237} : s = 115;
	{8'd203,8'd238} : s = 243;
	{8'd203,8'd239} : s = 238;
	{8'd203,8'd240} : s = 439;
	{8'd203,8'd241} : s = 237;
	{8'd203,8'd242} : s = 431;
	{8'd203,8'd243} : s = 415;
	{8'd203,8'd244} : s = 507;
	{8'd203,8'd245} : s = 7;
	{8'd203,8'd246} : s = 39;
	{8'd203,8'd247} : s = 30;
	{8'd203,8'd248} : s = 110;
	{8'd203,8'd249} : s = 29;
	{8'd203,8'd250} : s = 109;
	{8'd203,8'd251} : s = 107;
	{8'd203,8'd252} : s = 235;
	{8'd203,8'd253} : s = 27;
	{8'd203,8'd254} : s = 103;
	{8'd203,8'd255} : s = 94;
	{8'd204,8'd0} : s = 225;
	{8'd204,8'd1} : s = 369;
	{8'd204,8'd2} : s = 364;
	{8'd204,8'd3} : s = 470;
	{8'd204,8'd4} : s = 88;
	{8'd204,8'd5} : s = 216;
	{8'd204,8'd6} : s = 212;
	{8'd204,8'd7} : s = 362;
	{8'd204,8'd8} : s = 210;
	{8'd204,8'd9} : s = 361;
	{8'd204,8'd10} : s = 358;
	{8'd204,8'd11} : s = 469;
	{8'd204,8'd12} : s = 209;
	{8'd204,8'd13} : s = 357;
	{8'd204,8'd14} : s = 355;
	{8'd204,8'd15} : s = 467;
	{8'd204,8'd16} : s = 348;
	{8'd204,8'd17} : s = 462;
	{8'd204,8'd18} : s = 461;
	{8'd204,8'd19} : s = 505;
	{8'd204,8'd20} : s = 84;
	{8'd204,8'd21} : s = 204;
	{8'd204,8'd22} : s = 202;
	{8'd204,8'd23} : s = 346;
	{8'd204,8'd24} : s = 201;
	{8'd204,8'd25} : s = 345;
	{8'd204,8'd26} : s = 342;
	{8'd204,8'd27} : s = 459;
	{8'd204,8'd28} : s = 198;
	{8'd204,8'd29} : s = 341;
	{8'd204,8'd30} : s = 339;
	{8'd204,8'd31} : s = 455;
	{8'd204,8'd32} : s = 334;
	{8'd204,8'd33} : s = 444;
	{8'd204,8'd34} : s = 442;
	{8'd204,8'd35} : s = 502;
	{8'd204,8'd36} : s = 197;
	{8'd204,8'd37} : s = 333;
	{8'd204,8'd38} : s = 331;
	{8'd204,8'd39} : s = 441;
	{8'd204,8'd40} : s = 327;
	{8'd204,8'd41} : s = 438;
	{8'd204,8'd42} : s = 437;
	{8'd204,8'd43} : s = 501;
	{8'd204,8'd44} : s = 316;
	{8'd204,8'd45} : s = 435;
	{8'd204,8'd46} : s = 430;
	{8'd204,8'd47} : s = 499;
	{8'd204,8'd48} : s = 429;
	{8'd204,8'd49} : s = 494;
	{8'd204,8'd50} : s = 493;
	{8'd204,8'd51} : s = 510;
	{8'd204,8'd52} : s = 1;
	{8'd204,8'd53} : s = 18;
	{8'd204,8'd54} : s = 17;
	{8'd204,8'd55} : s = 82;
	{8'd204,8'd56} : s = 12;
	{8'd204,8'd57} : s = 81;
	{8'd204,8'd58} : s = 76;
	{8'd204,8'd59} : s = 195;
	{8'd204,8'd60} : s = 10;
	{8'd204,8'd61} : s = 74;
	{8'd204,8'd62} : s = 73;
	{8'd204,8'd63} : s = 184;
	{8'd204,8'd64} : s = 70;
	{8'd204,8'd65} : s = 180;
	{8'd204,8'd66} : s = 178;
	{8'd204,8'd67} : s = 314;
	{8'd204,8'd68} : s = 9;
	{8'd204,8'd69} : s = 69;
	{8'd204,8'd70} : s = 67;
	{8'd204,8'd71} : s = 177;
	{8'd204,8'd72} : s = 56;
	{8'd204,8'd73} : s = 172;
	{8'd204,8'd74} : s = 170;
	{8'd204,8'd75} : s = 313;
	{8'd204,8'd76} : s = 52;
	{8'd204,8'd77} : s = 169;
	{8'd204,8'd78} : s = 166;
	{8'd204,8'd79} : s = 310;
	{8'd204,8'd80} : s = 165;
	{8'd204,8'd81} : s = 309;
	{8'd204,8'd82} : s = 307;
	{8'd204,8'd83} : s = 427;
	{8'd204,8'd84} : s = 6;
	{8'd204,8'd85} : s = 50;
	{8'd204,8'd86} : s = 49;
	{8'd204,8'd87} : s = 163;
	{8'd204,8'd88} : s = 44;
	{8'd204,8'd89} : s = 156;
	{8'd204,8'd90} : s = 154;
	{8'd204,8'd91} : s = 302;
	{8'd204,8'd92} : s = 42;
	{8'd204,8'd93} : s = 153;
	{8'd204,8'd94} : s = 150;
	{8'd204,8'd95} : s = 301;
	{8'd204,8'd96} : s = 149;
	{8'd204,8'd97} : s = 299;
	{8'd204,8'd98} : s = 295;
	{8'd204,8'd99} : s = 423;
	{8'd204,8'd100} : s = 41;
	{8'd204,8'd101} : s = 147;
	{8'd204,8'd102} : s = 142;
	{8'd204,8'd103} : s = 286;
	{8'd204,8'd104} : s = 141;
	{8'd204,8'd105} : s = 285;
	{8'd204,8'd106} : s = 283;
	{8'd204,8'd107} : s = 414;
	{8'd204,8'd108} : s = 139;
	{8'd204,8'd109} : s = 279;
	{8'd204,8'd110} : s = 271;
	{8'd204,8'd111} : s = 413;
	{8'd204,8'd112} : s = 248;
	{8'd204,8'd113} : s = 411;
	{8'd204,8'd114} : s = 407;
	{8'd204,8'd115} : s = 491;
	{8'd204,8'd116} : s = 5;
	{8'd204,8'd117} : s = 38;
	{8'd204,8'd118} : s = 37;
	{8'd204,8'd119} : s = 135;
	{8'd204,8'd120} : s = 35;
	{8'd204,8'd121} : s = 120;
	{8'd204,8'd122} : s = 116;
	{8'd204,8'd123} : s = 244;
	{8'd204,8'd124} : s = 28;
	{8'd204,8'd125} : s = 114;
	{8'd204,8'd126} : s = 113;
	{8'd204,8'd127} : s = 242;
	{8'd204,8'd128} : s = 108;
	{8'd204,8'd129} : s = 241;
	{8'd204,8'd130} : s = 236;
	{8'd204,8'd131} : s = 399;
	{8'd204,8'd132} : s = 26;
	{8'd204,8'd133} : s = 106;
	{8'd204,8'd134} : s = 105;
	{8'd204,8'd135} : s = 234;
	{8'd204,8'd136} : s = 102;
	{8'd204,8'd137} : s = 233;
	{8'd204,8'd138} : s = 230;
	{8'd204,8'd139} : s = 380;
	{8'd204,8'd140} : s = 101;
	{8'd204,8'd141} : s = 229;
	{8'd204,8'd142} : s = 227;
	{8'd204,8'd143} : s = 378;
	{8'd204,8'd144} : s = 220;
	{8'd204,8'd145} : s = 377;
	{8'd204,8'd146} : s = 374;
	{8'd204,8'd147} : s = 487;
	{8'd204,8'd148} : s = 25;
	{8'd204,8'd149} : s = 99;
	{8'd204,8'd150} : s = 92;
	{8'd204,8'd151} : s = 218;
	{8'd204,8'd152} : s = 90;
	{8'd204,8'd153} : s = 217;
	{8'd204,8'd154} : s = 214;
	{8'd204,8'd155} : s = 373;
	{8'd204,8'd156} : s = 89;
	{8'd204,8'd157} : s = 213;
	{8'd204,8'd158} : s = 211;
	{8'd204,8'd159} : s = 371;
	{8'd204,8'd160} : s = 206;
	{8'd204,8'd161} : s = 366;
	{8'd204,8'd162} : s = 365;
	{8'd204,8'd163} : s = 478;
	{8'd204,8'd164} : s = 86;
	{8'd204,8'd165} : s = 205;
	{8'd204,8'd166} : s = 203;
	{8'd204,8'd167} : s = 363;
	{8'd204,8'd168} : s = 199;
	{8'd204,8'd169} : s = 359;
	{8'd204,8'd170} : s = 350;
	{8'd204,8'd171} : s = 477;
	{8'd204,8'd172} : s = 188;
	{8'd204,8'd173} : s = 349;
	{8'd204,8'd174} : s = 347;
	{8'd204,8'd175} : s = 475;
	{8'd204,8'd176} : s = 343;
	{8'd204,8'd177} : s = 471;
	{8'd204,8'd178} : s = 463;
	{8'd204,8'd179} : s = 509;
	{8'd204,8'd180} : s = 3;
	{8'd204,8'd181} : s = 22;
	{8'd204,8'd182} : s = 21;
	{8'd204,8'd183} : s = 85;
	{8'd204,8'd184} : s = 19;
	{8'd204,8'd185} : s = 83;
	{8'd204,8'd186} : s = 78;
	{8'd204,8'd187} : s = 186;
	{8'd204,8'd188} : s = 14;
	{8'd204,8'd189} : s = 77;
	{8'd204,8'd190} : s = 75;
	{8'd204,8'd191} : s = 185;
	{8'd204,8'd192} : s = 71;
	{8'd204,8'd193} : s = 182;
	{8'd204,8'd194} : s = 181;
	{8'd204,8'd195} : s = 335;
	{8'd204,8'd196} : s = 13;
	{8'd204,8'd197} : s = 60;
	{8'd204,8'd198} : s = 58;
	{8'd204,8'd199} : s = 179;
	{8'd204,8'd200} : s = 57;
	{8'd204,8'd201} : s = 174;
	{8'd204,8'd202} : s = 173;
	{8'd204,8'd203} : s = 318;
	{8'd204,8'd204} : s = 54;
	{8'd204,8'd205} : s = 171;
	{8'd204,8'd206} : s = 167;
	{8'd204,8'd207} : s = 317;
	{8'd204,8'd208} : s = 158;
	{8'd204,8'd209} : s = 315;
	{8'd204,8'd210} : s = 311;
	{8'd204,8'd211} : s = 446;
	{8'd204,8'd212} : s = 11;
	{8'd204,8'd213} : s = 53;
	{8'd204,8'd214} : s = 51;
	{8'd204,8'd215} : s = 157;
	{8'd204,8'd216} : s = 46;
	{8'd204,8'd217} : s = 155;
	{8'd204,8'd218} : s = 151;
	{8'd204,8'd219} : s = 303;
	{8'd204,8'd220} : s = 45;
	{8'd204,8'd221} : s = 143;
	{8'd204,8'd222} : s = 124;
	{8'd204,8'd223} : s = 287;
	{8'd204,8'd224} : s = 122;
	{8'd204,8'd225} : s = 252;
	{8'd204,8'd226} : s = 250;
	{8'd204,8'd227} : s = 445;
	{8'd204,8'd228} : s = 43;
	{8'd204,8'd229} : s = 121;
	{8'd204,8'd230} : s = 118;
	{8'd204,8'd231} : s = 249;
	{8'd204,8'd232} : s = 117;
	{8'd204,8'd233} : s = 246;
	{8'd204,8'd234} : s = 245;
	{8'd204,8'd235} : s = 443;
	{8'd204,8'd236} : s = 115;
	{8'd204,8'd237} : s = 243;
	{8'd204,8'd238} : s = 238;
	{8'd204,8'd239} : s = 439;
	{8'd204,8'd240} : s = 237;
	{8'd204,8'd241} : s = 431;
	{8'd204,8'd242} : s = 415;
	{8'd204,8'd243} : s = 507;
	{8'd204,8'd244} : s = 7;
	{8'd204,8'd245} : s = 39;
	{8'd204,8'd246} : s = 30;
	{8'd204,8'd247} : s = 110;
	{8'd204,8'd248} : s = 29;
	{8'd204,8'd249} : s = 109;
	{8'd204,8'd250} : s = 107;
	{8'd204,8'd251} : s = 235;
	{8'd204,8'd252} : s = 27;
	{8'd204,8'd253} : s = 103;
	{8'd204,8'd254} : s = 94;
	{8'd204,8'd255} : s = 231;
	{8'd205,8'd0} : s = 369;
	{8'd205,8'd1} : s = 364;
	{8'd205,8'd2} : s = 470;
	{8'd205,8'd3} : s = 88;
	{8'd205,8'd4} : s = 216;
	{8'd205,8'd5} : s = 212;
	{8'd205,8'd6} : s = 362;
	{8'd205,8'd7} : s = 210;
	{8'd205,8'd8} : s = 361;
	{8'd205,8'd9} : s = 358;
	{8'd205,8'd10} : s = 469;
	{8'd205,8'd11} : s = 209;
	{8'd205,8'd12} : s = 357;
	{8'd205,8'd13} : s = 355;
	{8'd205,8'd14} : s = 467;
	{8'd205,8'd15} : s = 348;
	{8'd205,8'd16} : s = 462;
	{8'd205,8'd17} : s = 461;
	{8'd205,8'd18} : s = 505;
	{8'd205,8'd19} : s = 84;
	{8'd205,8'd20} : s = 204;
	{8'd205,8'd21} : s = 202;
	{8'd205,8'd22} : s = 346;
	{8'd205,8'd23} : s = 201;
	{8'd205,8'd24} : s = 345;
	{8'd205,8'd25} : s = 342;
	{8'd205,8'd26} : s = 459;
	{8'd205,8'd27} : s = 198;
	{8'd205,8'd28} : s = 341;
	{8'd205,8'd29} : s = 339;
	{8'd205,8'd30} : s = 455;
	{8'd205,8'd31} : s = 334;
	{8'd205,8'd32} : s = 444;
	{8'd205,8'd33} : s = 442;
	{8'd205,8'd34} : s = 502;
	{8'd205,8'd35} : s = 197;
	{8'd205,8'd36} : s = 333;
	{8'd205,8'd37} : s = 331;
	{8'd205,8'd38} : s = 441;
	{8'd205,8'd39} : s = 327;
	{8'd205,8'd40} : s = 438;
	{8'd205,8'd41} : s = 437;
	{8'd205,8'd42} : s = 501;
	{8'd205,8'd43} : s = 316;
	{8'd205,8'd44} : s = 435;
	{8'd205,8'd45} : s = 430;
	{8'd205,8'd46} : s = 499;
	{8'd205,8'd47} : s = 429;
	{8'd205,8'd48} : s = 494;
	{8'd205,8'd49} : s = 493;
	{8'd205,8'd50} : s = 510;
	{8'd205,8'd51} : s = 1;
	{8'd205,8'd52} : s = 18;
	{8'd205,8'd53} : s = 17;
	{8'd205,8'd54} : s = 82;
	{8'd205,8'd55} : s = 12;
	{8'd205,8'd56} : s = 81;
	{8'd205,8'd57} : s = 76;
	{8'd205,8'd58} : s = 195;
	{8'd205,8'd59} : s = 10;
	{8'd205,8'd60} : s = 74;
	{8'd205,8'd61} : s = 73;
	{8'd205,8'd62} : s = 184;
	{8'd205,8'd63} : s = 70;
	{8'd205,8'd64} : s = 180;
	{8'd205,8'd65} : s = 178;
	{8'd205,8'd66} : s = 314;
	{8'd205,8'd67} : s = 9;
	{8'd205,8'd68} : s = 69;
	{8'd205,8'd69} : s = 67;
	{8'd205,8'd70} : s = 177;
	{8'd205,8'd71} : s = 56;
	{8'd205,8'd72} : s = 172;
	{8'd205,8'd73} : s = 170;
	{8'd205,8'd74} : s = 313;
	{8'd205,8'd75} : s = 52;
	{8'd205,8'd76} : s = 169;
	{8'd205,8'd77} : s = 166;
	{8'd205,8'd78} : s = 310;
	{8'd205,8'd79} : s = 165;
	{8'd205,8'd80} : s = 309;
	{8'd205,8'd81} : s = 307;
	{8'd205,8'd82} : s = 427;
	{8'd205,8'd83} : s = 6;
	{8'd205,8'd84} : s = 50;
	{8'd205,8'd85} : s = 49;
	{8'd205,8'd86} : s = 163;
	{8'd205,8'd87} : s = 44;
	{8'd205,8'd88} : s = 156;
	{8'd205,8'd89} : s = 154;
	{8'd205,8'd90} : s = 302;
	{8'd205,8'd91} : s = 42;
	{8'd205,8'd92} : s = 153;
	{8'd205,8'd93} : s = 150;
	{8'd205,8'd94} : s = 301;
	{8'd205,8'd95} : s = 149;
	{8'd205,8'd96} : s = 299;
	{8'd205,8'd97} : s = 295;
	{8'd205,8'd98} : s = 423;
	{8'd205,8'd99} : s = 41;
	{8'd205,8'd100} : s = 147;
	{8'd205,8'd101} : s = 142;
	{8'd205,8'd102} : s = 286;
	{8'd205,8'd103} : s = 141;
	{8'd205,8'd104} : s = 285;
	{8'd205,8'd105} : s = 283;
	{8'd205,8'd106} : s = 414;
	{8'd205,8'd107} : s = 139;
	{8'd205,8'd108} : s = 279;
	{8'd205,8'd109} : s = 271;
	{8'd205,8'd110} : s = 413;
	{8'd205,8'd111} : s = 248;
	{8'd205,8'd112} : s = 411;
	{8'd205,8'd113} : s = 407;
	{8'd205,8'd114} : s = 491;
	{8'd205,8'd115} : s = 5;
	{8'd205,8'd116} : s = 38;
	{8'd205,8'd117} : s = 37;
	{8'd205,8'd118} : s = 135;
	{8'd205,8'd119} : s = 35;
	{8'd205,8'd120} : s = 120;
	{8'd205,8'd121} : s = 116;
	{8'd205,8'd122} : s = 244;
	{8'd205,8'd123} : s = 28;
	{8'd205,8'd124} : s = 114;
	{8'd205,8'd125} : s = 113;
	{8'd205,8'd126} : s = 242;
	{8'd205,8'd127} : s = 108;
	{8'd205,8'd128} : s = 241;
	{8'd205,8'd129} : s = 236;
	{8'd205,8'd130} : s = 399;
	{8'd205,8'd131} : s = 26;
	{8'd205,8'd132} : s = 106;
	{8'd205,8'd133} : s = 105;
	{8'd205,8'd134} : s = 234;
	{8'd205,8'd135} : s = 102;
	{8'd205,8'd136} : s = 233;
	{8'd205,8'd137} : s = 230;
	{8'd205,8'd138} : s = 380;
	{8'd205,8'd139} : s = 101;
	{8'd205,8'd140} : s = 229;
	{8'd205,8'd141} : s = 227;
	{8'd205,8'd142} : s = 378;
	{8'd205,8'd143} : s = 220;
	{8'd205,8'd144} : s = 377;
	{8'd205,8'd145} : s = 374;
	{8'd205,8'd146} : s = 487;
	{8'd205,8'd147} : s = 25;
	{8'd205,8'd148} : s = 99;
	{8'd205,8'd149} : s = 92;
	{8'd205,8'd150} : s = 218;
	{8'd205,8'd151} : s = 90;
	{8'd205,8'd152} : s = 217;
	{8'd205,8'd153} : s = 214;
	{8'd205,8'd154} : s = 373;
	{8'd205,8'd155} : s = 89;
	{8'd205,8'd156} : s = 213;
	{8'd205,8'd157} : s = 211;
	{8'd205,8'd158} : s = 371;
	{8'd205,8'd159} : s = 206;
	{8'd205,8'd160} : s = 366;
	{8'd205,8'd161} : s = 365;
	{8'd205,8'd162} : s = 478;
	{8'd205,8'd163} : s = 86;
	{8'd205,8'd164} : s = 205;
	{8'd205,8'd165} : s = 203;
	{8'd205,8'd166} : s = 363;
	{8'd205,8'd167} : s = 199;
	{8'd205,8'd168} : s = 359;
	{8'd205,8'd169} : s = 350;
	{8'd205,8'd170} : s = 477;
	{8'd205,8'd171} : s = 188;
	{8'd205,8'd172} : s = 349;
	{8'd205,8'd173} : s = 347;
	{8'd205,8'd174} : s = 475;
	{8'd205,8'd175} : s = 343;
	{8'd205,8'd176} : s = 471;
	{8'd205,8'd177} : s = 463;
	{8'd205,8'd178} : s = 509;
	{8'd205,8'd179} : s = 3;
	{8'd205,8'd180} : s = 22;
	{8'd205,8'd181} : s = 21;
	{8'd205,8'd182} : s = 85;
	{8'd205,8'd183} : s = 19;
	{8'd205,8'd184} : s = 83;
	{8'd205,8'd185} : s = 78;
	{8'd205,8'd186} : s = 186;
	{8'd205,8'd187} : s = 14;
	{8'd205,8'd188} : s = 77;
	{8'd205,8'd189} : s = 75;
	{8'd205,8'd190} : s = 185;
	{8'd205,8'd191} : s = 71;
	{8'd205,8'd192} : s = 182;
	{8'd205,8'd193} : s = 181;
	{8'd205,8'd194} : s = 335;
	{8'd205,8'd195} : s = 13;
	{8'd205,8'd196} : s = 60;
	{8'd205,8'd197} : s = 58;
	{8'd205,8'd198} : s = 179;
	{8'd205,8'd199} : s = 57;
	{8'd205,8'd200} : s = 174;
	{8'd205,8'd201} : s = 173;
	{8'd205,8'd202} : s = 318;
	{8'd205,8'd203} : s = 54;
	{8'd205,8'd204} : s = 171;
	{8'd205,8'd205} : s = 167;
	{8'd205,8'd206} : s = 317;
	{8'd205,8'd207} : s = 158;
	{8'd205,8'd208} : s = 315;
	{8'd205,8'd209} : s = 311;
	{8'd205,8'd210} : s = 446;
	{8'd205,8'd211} : s = 11;
	{8'd205,8'd212} : s = 53;
	{8'd205,8'd213} : s = 51;
	{8'd205,8'd214} : s = 157;
	{8'd205,8'd215} : s = 46;
	{8'd205,8'd216} : s = 155;
	{8'd205,8'd217} : s = 151;
	{8'd205,8'd218} : s = 303;
	{8'd205,8'd219} : s = 45;
	{8'd205,8'd220} : s = 143;
	{8'd205,8'd221} : s = 124;
	{8'd205,8'd222} : s = 287;
	{8'd205,8'd223} : s = 122;
	{8'd205,8'd224} : s = 252;
	{8'd205,8'd225} : s = 250;
	{8'd205,8'd226} : s = 445;
	{8'd205,8'd227} : s = 43;
	{8'd205,8'd228} : s = 121;
	{8'd205,8'd229} : s = 118;
	{8'd205,8'd230} : s = 249;
	{8'd205,8'd231} : s = 117;
	{8'd205,8'd232} : s = 246;
	{8'd205,8'd233} : s = 245;
	{8'd205,8'd234} : s = 443;
	{8'd205,8'd235} : s = 115;
	{8'd205,8'd236} : s = 243;
	{8'd205,8'd237} : s = 238;
	{8'd205,8'd238} : s = 439;
	{8'd205,8'd239} : s = 237;
	{8'd205,8'd240} : s = 431;
	{8'd205,8'd241} : s = 415;
	{8'd205,8'd242} : s = 507;
	{8'd205,8'd243} : s = 7;
	{8'd205,8'd244} : s = 39;
	{8'd205,8'd245} : s = 30;
	{8'd205,8'd246} : s = 110;
	{8'd205,8'd247} : s = 29;
	{8'd205,8'd248} : s = 109;
	{8'd205,8'd249} : s = 107;
	{8'd205,8'd250} : s = 235;
	{8'd205,8'd251} : s = 27;
	{8'd205,8'd252} : s = 103;
	{8'd205,8'd253} : s = 94;
	{8'd205,8'd254} : s = 231;
	{8'd205,8'd255} : s = 93;
	{8'd206,8'd0} : s = 364;
	{8'd206,8'd1} : s = 470;
	{8'd206,8'd2} : s = 88;
	{8'd206,8'd3} : s = 216;
	{8'd206,8'd4} : s = 212;
	{8'd206,8'd5} : s = 362;
	{8'd206,8'd6} : s = 210;
	{8'd206,8'd7} : s = 361;
	{8'd206,8'd8} : s = 358;
	{8'd206,8'd9} : s = 469;
	{8'd206,8'd10} : s = 209;
	{8'd206,8'd11} : s = 357;
	{8'd206,8'd12} : s = 355;
	{8'd206,8'd13} : s = 467;
	{8'd206,8'd14} : s = 348;
	{8'd206,8'd15} : s = 462;
	{8'd206,8'd16} : s = 461;
	{8'd206,8'd17} : s = 505;
	{8'd206,8'd18} : s = 84;
	{8'd206,8'd19} : s = 204;
	{8'd206,8'd20} : s = 202;
	{8'd206,8'd21} : s = 346;
	{8'd206,8'd22} : s = 201;
	{8'd206,8'd23} : s = 345;
	{8'd206,8'd24} : s = 342;
	{8'd206,8'd25} : s = 459;
	{8'd206,8'd26} : s = 198;
	{8'd206,8'd27} : s = 341;
	{8'd206,8'd28} : s = 339;
	{8'd206,8'd29} : s = 455;
	{8'd206,8'd30} : s = 334;
	{8'd206,8'd31} : s = 444;
	{8'd206,8'd32} : s = 442;
	{8'd206,8'd33} : s = 502;
	{8'd206,8'd34} : s = 197;
	{8'd206,8'd35} : s = 333;
	{8'd206,8'd36} : s = 331;
	{8'd206,8'd37} : s = 441;
	{8'd206,8'd38} : s = 327;
	{8'd206,8'd39} : s = 438;
	{8'd206,8'd40} : s = 437;
	{8'd206,8'd41} : s = 501;
	{8'd206,8'd42} : s = 316;
	{8'd206,8'd43} : s = 435;
	{8'd206,8'd44} : s = 430;
	{8'd206,8'd45} : s = 499;
	{8'd206,8'd46} : s = 429;
	{8'd206,8'd47} : s = 494;
	{8'd206,8'd48} : s = 493;
	{8'd206,8'd49} : s = 510;
	{8'd206,8'd50} : s = 1;
	{8'd206,8'd51} : s = 18;
	{8'd206,8'd52} : s = 17;
	{8'd206,8'd53} : s = 82;
	{8'd206,8'd54} : s = 12;
	{8'd206,8'd55} : s = 81;
	{8'd206,8'd56} : s = 76;
	{8'd206,8'd57} : s = 195;
	{8'd206,8'd58} : s = 10;
	{8'd206,8'd59} : s = 74;
	{8'd206,8'd60} : s = 73;
	{8'd206,8'd61} : s = 184;
	{8'd206,8'd62} : s = 70;
	{8'd206,8'd63} : s = 180;
	{8'd206,8'd64} : s = 178;
	{8'd206,8'd65} : s = 314;
	{8'd206,8'd66} : s = 9;
	{8'd206,8'd67} : s = 69;
	{8'd206,8'd68} : s = 67;
	{8'd206,8'd69} : s = 177;
	{8'd206,8'd70} : s = 56;
	{8'd206,8'd71} : s = 172;
	{8'd206,8'd72} : s = 170;
	{8'd206,8'd73} : s = 313;
	{8'd206,8'd74} : s = 52;
	{8'd206,8'd75} : s = 169;
	{8'd206,8'd76} : s = 166;
	{8'd206,8'd77} : s = 310;
	{8'd206,8'd78} : s = 165;
	{8'd206,8'd79} : s = 309;
	{8'd206,8'd80} : s = 307;
	{8'd206,8'd81} : s = 427;
	{8'd206,8'd82} : s = 6;
	{8'd206,8'd83} : s = 50;
	{8'd206,8'd84} : s = 49;
	{8'd206,8'd85} : s = 163;
	{8'd206,8'd86} : s = 44;
	{8'd206,8'd87} : s = 156;
	{8'd206,8'd88} : s = 154;
	{8'd206,8'd89} : s = 302;
	{8'd206,8'd90} : s = 42;
	{8'd206,8'd91} : s = 153;
	{8'd206,8'd92} : s = 150;
	{8'd206,8'd93} : s = 301;
	{8'd206,8'd94} : s = 149;
	{8'd206,8'd95} : s = 299;
	{8'd206,8'd96} : s = 295;
	{8'd206,8'd97} : s = 423;
	{8'd206,8'd98} : s = 41;
	{8'd206,8'd99} : s = 147;
	{8'd206,8'd100} : s = 142;
	{8'd206,8'd101} : s = 286;
	{8'd206,8'd102} : s = 141;
	{8'd206,8'd103} : s = 285;
	{8'd206,8'd104} : s = 283;
	{8'd206,8'd105} : s = 414;
	{8'd206,8'd106} : s = 139;
	{8'd206,8'd107} : s = 279;
	{8'd206,8'd108} : s = 271;
	{8'd206,8'd109} : s = 413;
	{8'd206,8'd110} : s = 248;
	{8'd206,8'd111} : s = 411;
	{8'd206,8'd112} : s = 407;
	{8'd206,8'd113} : s = 491;
	{8'd206,8'd114} : s = 5;
	{8'd206,8'd115} : s = 38;
	{8'd206,8'd116} : s = 37;
	{8'd206,8'd117} : s = 135;
	{8'd206,8'd118} : s = 35;
	{8'd206,8'd119} : s = 120;
	{8'd206,8'd120} : s = 116;
	{8'd206,8'd121} : s = 244;
	{8'd206,8'd122} : s = 28;
	{8'd206,8'd123} : s = 114;
	{8'd206,8'd124} : s = 113;
	{8'd206,8'd125} : s = 242;
	{8'd206,8'd126} : s = 108;
	{8'd206,8'd127} : s = 241;
	{8'd206,8'd128} : s = 236;
	{8'd206,8'd129} : s = 399;
	{8'd206,8'd130} : s = 26;
	{8'd206,8'd131} : s = 106;
	{8'd206,8'd132} : s = 105;
	{8'd206,8'd133} : s = 234;
	{8'd206,8'd134} : s = 102;
	{8'd206,8'd135} : s = 233;
	{8'd206,8'd136} : s = 230;
	{8'd206,8'd137} : s = 380;
	{8'd206,8'd138} : s = 101;
	{8'd206,8'd139} : s = 229;
	{8'd206,8'd140} : s = 227;
	{8'd206,8'd141} : s = 378;
	{8'd206,8'd142} : s = 220;
	{8'd206,8'd143} : s = 377;
	{8'd206,8'd144} : s = 374;
	{8'd206,8'd145} : s = 487;
	{8'd206,8'd146} : s = 25;
	{8'd206,8'd147} : s = 99;
	{8'd206,8'd148} : s = 92;
	{8'd206,8'd149} : s = 218;
	{8'd206,8'd150} : s = 90;
	{8'd206,8'd151} : s = 217;
	{8'd206,8'd152} : s = 214;
	{8'd206,8'd153} : s = 373;
	{8'd206,8'd154} : s = 89;
	{8'd206,8'd155} : s = 213;
	{8'd206,8'd156} : s = 211;
	{8'd206,8'd157} : s = 371;
	{8'd206,8'd158} : s = 206;
	{8'd206,8'd159} : s = 366;
	{8'd206,8'd160} : s = 365;
	{8'd206,8'd161} : s = 478;
	{8'd206,8'd162} : s = 86;
	{8'd206,8'd163} : s = 205;
	{8'd206,8'd164} : s = 203;
	{8'd206,8'd165} : s = 363;
	{8'd206,8'd166} : s = 199;
	{8'd206,8'd167} : s = 359;
	{8'd206,8'd168} : s = 350;
	{8'd206,8'd169} : s = 477;
	{8'd206,8'd170} : s = 188;
	{8'd206,8'd171} : s = 349;
	{8'd206,8'd172} : s = 347;
	{8'd206,8'd173} : s = 475;
	{8'd206,8'd174} : s = 343;
	{8'd206,8'd175} : s = 471;
	{8'd206,8'd176} : s = 463;
	{8'd206,8'd177} : s = 509;
	{8'd206,8'd178} : s = 3;
	{8'd206,8'd179} : s = 22;
	{8'd206,8'd180} : s = 21;
	{8'd206,8'd181} : s = 85;
	{8'd206,8'd182} : s = 19;
	{8'd206,8'd183} : s = 83;
	{8'd206,8'd184} : s = 78;
	{8'd206,8'd185} : s = 186;
	{8'd206,8'd186} : s = 14;
	{8'd206,8'd187} : s = 77;
	{8'd206,8'd188} : s = 75;
	{8'd206,8'd189} : s = 185;
	{8'd206,8'd190} : s = 71;
	{8'd206,8'd191} : s = 182;
	{8'd206,8'd192} : s = 181;
	{8'd206,8'd193} : s = 335;
	{8'd206,8'd194} : s = 13;
	{8'd206,8'd195} : s = 60;
	{8'd206,8'd196} : s = 58;
	{8'd206,8'd197} : s = 179;
	{8'd206,8'd198} : s = 57;
	{8'd206,8'd199} : s = 174;
	{8'd206,8'd200} : s = 173;
	{8'd206,8'd201} : s = 318;
	{8'd206,8'd202} : s = 54;
	{8'd206,8'd203} : s = 171;
	{8'd206,8'd204} : s = 167;
	{8'd206,8'd205} : s = 317;
	{8'd206,8'd206} : s = 158;
	{8'd206,8'd207} : s = 315;
	{8'd206,8'd208} : s = 311;
	{8'd206,8'd209} : s = 446;
	{8'd206,8'd210} : s = 11;
	{8'd206,8'd211} : s = 53;
	{8'd206,8'd212} : s = 51;
	{8'd206,8'd213} : s = 157;
	{8'd206,8'd214} : s = 46;
	{8'd206,8'd215} : s = 155;
	{8'd206,8'd216} : s = 151;
	{8'd206,8'd217} : s = 303;
	{8'd206,8'd218} : s = 45;
	{8'd206,8'd219} : s = 143;
	{8'd206,8'd220} : s = 124;
	{8'd206,8'd221} : s = 287;
	{8'd206,8'd222} : s = 122;
	{8'd206,8'd223} : s = 252;
	{8'd206,8'd224} : s = 250;
	{8'd206,8'd225} : s = 445;
	{8'd206,8'd226} : s = 43;
	{8'd206,8'd227} : s = 121;
	{8'd206,8'd228} : s = 118;
	{8'd206,8'd229} : s = 249;
	{8'd206,8'd230} : s = 117;
	{8'd206,8'd231} : s = 246;
	{8'd206,8'd232} : s = 245;
	{8'd206,8'd233} : s = 443;
	{8'd206,8'd234} : s = 115;
	{8'd206,8'd235} : s = 243;
	{8'd206,8'd236} : s = 238;
	{8'd206,8'd237} : s = 439;
	{8'd206,8'd238} : s = 237;
	{8'd206,8'd239} : s = 431;
	{8'd206,8'd240} : s = 415;
	{8'd206,8'd241} : s = 507;
	{8'd206,8'd242} : s = 7;
	{8'd206,8'd243} : s = 39;
	{8'd206,8'd244} : s = 30;
	{8'd206,8'd245} : s = 110;
	{8'd206,8'd246} : s = 29;
	{8'd206,8'd247} : s = 109;
	{8'd206,8'd248} : s = 107;
	{8'd206,8'd249} : s = 235;
	{8'd206,8'd250} : s = 27;
	{8'd206,8'd251} : s = 103;
	{8'd206,8'd252} : s = 94;
	{8'd206,8'd253} : s = 231;
	{8'd206,8'd254} : s = 93;
	{8'd206,8'd255} : s = 222;
	{8'd207,8'd0} : s = 470;
	{8'd207,8'd1} : s = 88;
	{8'd207,8'd2} : s = 216;
	{8'd207,8'd3} : s = 212;
	{8'd207,8'd4} : s = 362;
	{8'd207,8'd5} : s = 210;
	{8'd207,8'd6} : s = 361;
	{8'd207,8'd7} : s = 358;
	{8'd207,8'd8} : s = 469;
	{8'd207,8'd9} : s = 209;
	{8'd207,8'd10} : s = 357;
	{8'd207,8'd11} : s = 355;
	{8'd207,8'd12} : s = 467;
	{8'd207,8'd13} : s = 348;
	{8'd207,8'd14} : s = 462;
	{8'd207,8'd15} : s = 461;
	{8'd207,8'd16} : s = 505;
	{8'd207,8'd17} : s = 84;
	{8'd207,8'd18} : s = 204;
	{8'd207,8'd19} : s = 202;
	{8'd207,8'd20} : s = 346;
	{8'd207,8'd21} : s = 201;
	{8'd207,8'd22} : s = 345;
	{8'd207,8'd23} : s = 342;
	{8'd207,8'd24} : s = 459;
	{8'd207,8'd25} : s = 198;
	{8'd207,8'd26} : s = 341;
	{8'd207,8'd27} : s = 339;
	{8'd207,8'd28} : s = 455;
	{8'd207,8'd29} : s = 334;
	{8'd207,8'd30} : s = 444;
	{8'd207,8'd31} : s = 442;
	{8'd207,8'd32} : s = 502;
	{8'd207,8'd33} : s = 197;
	{8'd207,8'd34} : s = 333;
	{8'd207,8'd35} : s = 331;
	{8'd207,8'd36} : s = 441;
	{8'd207,8'd37} : s = 327;
	{8'd207,8'd38} : s = 438;
	{8'd207,8'd39} : s = 437;
	{8'd207,8'd40} : s = 501;
	{8'd207,8'd41} : s = 316;
	{8'd207,8'd42} : s = 435;
	{8'd207,8'd43} : s = 430;
	{8'd207,8'd44} : s = 499;
	{8'd207,8'd45} : s = 429;
	{8'd207,8'd46} : s = 494;
	{8'd207,8'd47} : s = 493;
	{8'd207,8'd48} : s = 510;
	{8'd207,8'd49} : s = 1;
	{8'd207,8'd50} : s = 18;
	{8'd207,8'd51} : s = 17;
	{8'd207,8'd52} : s = 82;
	{8'd207,8'd53} : s = 12;
	{8'd207,8'd54} : s = 81;
	{8'd207,8'd55} : s = 76;
	{8'd207,8'd56} : s = 195;
	{8'd207,8'd57} : s = 10;
	{8'd207,8'd58} : s = 74;
	{8'd207,8'd59} : s = 73;
	{8'd207,8'd60} : s = 184;
	{8'd207,8'd61} : s = 70;
	{8'd207,8'd62} : s = 180;
	{8'd207,8'd63} : s = 178;
	{8'd207,8'd64} : s = 314;
	{8'd207,8'd65} : s = 9;
	{8'd207,8'd66} : s = 69;
	{8'd207,8'd67} : s = 67;
	{8'd207,8'd68} : s = 177;
	{8'd207,8'd69} : s = 56;
	{8'd207,8'd70} : s = 172;
	{8'd207,8'd71} : s = 170;
	{8'd207,8'd72} : s = 313;
	{8'd207,8'd73} : s = 52;
	{8'd207,8'd74} : s = 169;
	{8'd207,8'd75} : s = 166;
	{8'd207,8'd76} : s = 310;
	{8'd207,8'd77} : s = 165;
	{8'd207,8'd78} : s = 309;
	{8'd207,8'd79} : s = 307;
	{8'd207,8'd80} : s = 427;
	{8'd207,8'd81} : s = 6;
	{8'd207,8'd82} : s = 50;
	{8'd207,8'd83} : s = 49;
	{8'd207,8'd84} : s = 163;
	{8'd207,8'd85} : s = 44;
	{8'd207,8'd86} : s = 156;
	{8'd207,8'd87} : s = 154;
	{8'd207,8'd88} : s = 302;
	{8'd207,8'd89} : s = 42;
	{8'd207,8'd90} : s = 153;
	{8'd207,8'd91} : s = 150;
	{8'd207,8'd92} : s = 301;
	{8'd207,8'd93} : s = 149;
	{8'd207,8'd94} : s = 299;
	{8'd207,8'd95} : s = 295;
	{8'd207,8'd96} : s = 423;
	{8'd207,8'd97} : s = 41;
	{8'd207,8'd98} : s = 147;
	{8'd207,8'd99} : s = 142;
	{8'd207,8'd100} : s = 286;
	{8'd207,8'd101} : s = 141;
	{8'd207,8'd102} : s = 285;
	{8'd207,8'd103} : s = 283;
	{8'd207,8'd104} : s = 414;
	{8'd207,8'd105} : s = 139;
	{8'd207,8'd106} : s = 279;
	{8'd207,8'd107} : s = 271;
	{8'd207,8'd108} : s = 413;
	{8'd207,8'd109} : s = 248;
	{8'd207,8'd110} : s = 411;
	{8'd207,8'd111} : s = 407;
	{8'd207,8'd112} : s = 491;
	{8'd207,8'd113} : s = 5;
	{8'd207,8'd114} : s = 38;
	{8'd207,8'd115} : s = 37;
	{8'd207,8'd116} : s = 135;
	{8'd207,8'd117} : s = 35;
	{8'd207,8'd118} : s = 120;
	{8'd207,8'd119} : s = 116;
	{8'd207,8'd120} : s = 244;
	{8'd207,8'd121} : s = 28;
	{8'd207,8'd122} : s = 114;
	{8'd207,8'd123} : s = 113;
	{8'd207,8'd124} : s = 242;
	{8'd207,8'd125} : s = 108;
	{8'd207,8'd126} : s = 241;
	{8'd207,8'd127} : s = 236;
	{8'd207,8'd128} : s = 399;
	{8'd207,8'd129} : s = 26;
	{8'd207,8'd130} : s = 106;
	{8'd207,8'd131} : s = 105;
	{8'd207,8'd132} : s = 234;
	{8'd207,8'd133} : s = 102;
	{8'd207,8'd134} : s = 233;
	{8'd207,8'd135} : s = 230;
	{8'd207,8'd136} : s = 380;
	{8'd207,8'd137} : s = 101;
	{8'd207,8'd138} : s = 229;
	{8'd207,8'd139} : s = 227;
	{8'd207,8'd140} : s = 378;
	{8'd207,8'd141} : s = 220;
	{8'd207,8'd142} : s = 377;
	{8'd207,8'd143} : s = 374;
	{8'd207,8'd144} : s = 487;
	{8'd207,8'd145} : s = 25;
	{8'd207,8'd146} : s = 99;
	{8'd207,8'd147} : s = 92;
	{8'd207,8'd148} : s = 218;
	{8'd207,8'd149} : s = 90;
	{8'd207,8'd150} : s = 217;
	{8'd207,8'd151} : s = 214;
	{8'd207,8'd152} : s = 373;
	{8'd207,8'd153} : s = 89;
	{8'd207,8'd154} : s = 213;
	{8'd207,8'd155} : s = 211;
	{8'd207,8'd156} : s = 371;
	{8'd207,8'd157} : s = 206;
	{8'd207,8'd158} : s = 366;
	{8'd207,8'd159} : s = 365;
	{8'd207,8'd160} : s = 478;
	{8'd207,8'd161} : s = 86;
	{8'd207,8'd162} : s = 205;
	{8'd207,8'd163} : s = 203;
	{8'd207,8'd164} : s = 363;
	{8'd207,8'd165} : s = 199;
	{8'd207,8'd166} : s = 359;
	{8'd207,8'd167} : s = 350;
	{8'd207,8'd168} : s = 477;
	{8'd207,8'd169} : s = 188;
	{8'd207,8'd170} : s = 349;
	{8'd207,8'd171} : s = 347;
	{8'd207,8'd172} : s = 475;
	{8'd207,8'd173} : s = 343;
	{8'd207,8'd174} : s = 471;
	{8'd207,8'd175} : s = 463;
	{8'd207,8'd176} : s = 509;
	{8'd207,8'd177} : s = 3;
	{8'd207,8'd178} : s = 22;
	{8'd207,8'd179} : s = 21;
	{8'd207,8'd180} : s = 85;
	{8'd207,8'd181} : s = 19;
	{8'd207,8'd182} : s = 83;
	{8'd207,8'd183} : s = 78;
	{8'd207,8'd184} : s = 186;
	{8'd207,8'd185} : s = 14;
	{8'd207,8'd186} : s = 77;
	{8'd207,8'd187} : s = 75;
	{8'd207,8'd188} : s = 185;
	{8'd207,8'd189} : s = 71;
	{8'd207,8'd190} : s = 182;
	{8'd207,8'd191} : s = 181;
	{8'd207,8'd192} : s = 335;
	{8'd207,8'd193} : s = 13;
	{8'd207,8'd194} : s = 60;
	{8'd207,8'd195} : s = 58;
	{8'd207,8'd196} : s = 179;
	{8'd207,8'd197} : s = 57;
	{8'd207,8'd198} : s = 174;
	{8'd207,8'd199} : s = 173;
	{8'd207,8'd200} : s = 318;
	{8'd207,8'd201} : s = 54;
	{8'd207,8'd202} : s = 171;
	{8'd207,8'd203} : s = 167;
	{8'd207,8'd204} : s = 317;
	{8'd207,8'd205} : s = 158;
	{8'd207,8'd206} : s = 315;
	{8'd207,8'd207} : s = 311;
	{8'd207,8'd208} : s = 446;
	{8'd207,8'd209} : s = 11;
	{8'd207,8'd210} : s = 53;
	{8'd207,8'd211} : s = 51;
	{8'd207,8'd212} : s = 157;
	{8'd207,8'd213} : s = 46;
	{8'd207,8'd214} : s = 155;
	{8'd207,8'd215} : s = 151;
	{8'd207,8'd216} : s = 303;
	{8'd207,8'd217} : s = 45;
	{8'd207,8'd218} : s = 143;
	{8'd207,8'd219} : s = 124;
	{8'd207,8'd220} : s = 287;
	{8'd207,8'd221} : s = 122;
	{8'd207,8'd222} : s = 252;
	{8'd207,8'd223} : s = 250;
	{8'd207,8'd224} : s = 445;
	{8'd207,8'd225} : s = 43;
	{8'd207,8'd226} : s = 121;
	{8'd207,8'd227} : s = 118;
	{8'd207,8'd228} : s = 249;
	{8'd207,8'd229} : s = 117;
	{8'd207,8'd230} : s = 246;
	{8'd207,8'd231} : s = 245;
	{8'd207,8'd232} : s = 443;
	{8'd207,8'd233} : s = 115;
	{8'd207,8'd234} : s = 243;
	{8'd207,8'd235} : s = 238;
	{8'd207,8'd236} : s = 439;
	{8'd207,8'd237} : s = 237;
	{8'd207,8'd238} : s = 431;
	{8'd207,8'd239} : s = 415;
	{8'd207,8'd240} : s = 507;
	{8'd207,8'd241} : s = 7;
	{8'd207,8'd242} : s = 39;
	{8'd207,8'd243} : s = 30;
	{8'd207,8'd244} : s = 110;
	{8'd207,8'd245} : s = 29;
	{8'd207,8'd246} : s = 109;
	{8'd207,8'd247} : s = 107;
	{8'd207,8'd248} : s = 235;
	{8'd207,8'd249} : s = 27;
	{8'd207,8'd250} : s = 103;
	{8'd207,8'd251} : s = 94;
	{8'd207,8'd252} : s = 231;
	{8'd207,8'd253} : s = 93;
	{8'd207,8'd254} : s = 222;
	{8'd207,8'd255} : s = 221;
	{8'd208,8'd0} : s = 88;
	{8'd208,8'd1} : s = 216;
	{8'd208,8'd2} : s = 212;
	{8'd208,8'd3} : s = 362;
	{8'd208,8'd4} : s = 210;
	{8'd208,8'd5} : s = 361;
	{8'd208,8'd6} : s = 358;
	{8'd208,8'd7} : s = 469;
	{8'd208,8'd8} : s = 209;
	{8'd208,8'd9} : s = 357;
	{8'd208,8'd10} : s = 355;
	{8'd208,8'd11} : s = 467;
	{8'd208,8'd12} : s = 348;
	{8'd208,8'd13} : s = 462;
	{8'd208,8'd14} : s = 461;
	{8'd208,8'd15} : s = 505;
	{8'd208,8'd16} : s = 84;
	{8'd208,8'd17} : s = 204;
	{8'd208,8'd18} : s = 202;
	{8'd208,8'd19} : s = 346;
	{8'd208,8'd20} : s = 201;
	{8'd208,8'd21} : s = 345;
	{8'd208,8'd22} : s = 342;
	{8'd208,8'd23} : s = 459;
	{8'd208,8'd24} : s = 198;
	{8'd208,8'd25} : s = 341;
	{8'd208,8'd26} : s = 339;
	{8'd208,8'd27} : s = 455;
	{8'd208,8'd28} : s = 334;
	{8'd208,8'd29} : s = 444;
	{8'd208,8'd30} : s = 442;
	{8'd208,8'd31} : s = 502;
	{8'd208,8'd32} : s = 197;
	{8'd208,8'd33} : s = 333;
	{8'd208,8'd34} : s = 331;
	{8'd208,8'd35} : s = 441;
	{8'd208,8'd36} : s = 327;
	{8'd208,8'd37} : s = 438;
	{8'd208,8'd38} : s = 437;
	{8'd208,8'd39} : s = 501;
	{8'd208,8'd40} : s = 316;
	{8'd208,8'd41} : s = 435;
	{8'd208,8'd42} : s = 430;
	{8'd208,8'd43} : s = 499;
	{8'd208,8'd44} : s = 429;
	{8'd208,8'd45} : s = 494;
	{8'd208,8'd46} : s = 493;
	{8'd208,8'd47} : s = 510;
	{8'd208,8'd48} : s = 1;
	{8'd208,8'd49} : s = 18;
	{8'd208,8'd50} : s = 17;
	{8'd208,8'd51} : s = 82;
	{8'd208,8'd52} : s = 12;
	{8'd208,8'd53} : s = 81;
	{8'd208,8'd54} : s = 76;
	{8'd208,8'd55} : s = 195;
	{8'd208,8'd56} : s = 10;
	{8'd208,8'd57} : s = 74;
	{8'd208,8'd58} : s = 73;
	{8'd208,8'd59} : s = 184;
	{8'd208,8'd60} : s = 70;
	{8'd208,8'd61} : s = 180;
	{8'd208,8'd62} : s = 178;
	{8'd208,8'd63} : s = 314;
	{8'd208,8'd64} : s = 9;
	{8'd208,8'd65} : s = 69;
	{8'd208,8'd66} : s = 67;
	{8'd208,8'd67} : s = 177;
	{8'd208,8'd68} : s = 56;
	{8'd208,8'd69} : s = 172;
	{8'd208,8'd70} : s = 170;
	{8'd208,8'd71} : s = 313;
	{8'd208,8'd72} : s = 52;
	{8'd208,8'd73} : s = 169;
	{8'd208,8'd74} : s = 166;
	{8'd208,8'd75} : s = 310;
	{8'd208,8'd76} : s = 165;
	{8'd208,8'd77} : s = 309;
	{8'd208,8'd78} : s = 307;
	{8'd208,8'd79} : s = 427;
	{8'd208,8'd80} : s = 6;
	{8'd208,8'd81} : s = 50;
	{8'd208,8'd82} : s = 49;
	{8'd208,8'd83} : s = 163;
	{8'd208,8'd84} : s = 44;
	{8'd208,8'd85} : s = 156;
	{8'd208,8'd86} : s = 154;
	{8'd208,8'd87} : s = 302;
	{8'd208,8'd88} : s = 42;
	{8'd208,8'd89} : s = 153;
	{8'd208,8'd90} : s = 150;
	{8'd208,8'd91} : s = 301;
	{8'd208,8'd92} : s = 149;
	{8'd208,8'd93} : s = 299;
	{8'd208,8'd94} : s = 295;
	{8'd208,8'd95} : s = 423;
	{8'd208,8'd96} : s = 41;
	{8'd208,8'd97} : s = 147;
	{8'd208,8'd98} : s = 142;
	{8'd208,8'd99} : s = 286;
	{8'd208,8'd100} : s = 141;
	{8'd208,8'd101} : s = 285;
	{8'd208,8'd102} : s = 283;
	{8'd208,8'd103} : s = 414;
	{8'd208,8'd104} : s = 139;
	{8'd208,8'd105} : s = 279;
	{8'd208,8'd106} : s = 271;
	{8'd208,8'd107} : s = 413;
	{8'd208,8'd108} : s = 248;
	{8'd208,8'd109} : s = 411;
	{8'd208,8'd110} : s = 407;
	{8'd208,8'd111} : s = 491;
	{8'd208,8'd112} : s = 5;
	{8'd208,8'd113} : s = 38;
	{8'd208,8'd114} : s = 37;
	{8'd208,8'd115} : s = 135;
	{8'd208,8'd116} : s = 35;
	{8'd208,8'd117} : s = 120;
	{8'd208,8'd118} : s = 116;
	{8'd208,8'd119} : s = 244;
	{8'd208,8'd120} : s = 28;
	{8'd208,8'd121} : s = 114;
	{8'd208,8'd122} : s = 113;
	{8'd208,8'd123} : s = 242;
	{8'd208,8'd124} : s = 108;
	{8'd208,8'd125} : s = 241;
	{8'd208,8'd126} : s = 236;
	{8'd208,8'd127} : s = 399;
	{8'd208,8'd128} : s = 26;
	{8'd208,8'd129} : s = 106;
	{8'd208,8'd130} : s = 105;
	{8'd208,8'd131} : s = 234;
	{8'd208,8'd132} : s = 102;
	{8'd208,8'd133} : s = 233;
	{8'd208,8'd134} : s = 230;
	{8'd208,8'd135} : s = 380;
	{8'd208,8'd136} : s = 101;
	{8'd208,8'd137} : s = 229;
	{8'd208,8'd138} : s = 227;
	{8'd208,8'd139} : s = 378;
	{8'd208,8'd140} : s = 220;
	{8'd208,8'd141} : s = 377;
	{8'd208,8'd142} : s = 374;
	{8'd208,8'd143} : s = 487;
	{8'd208,8'd144} : s = 25;
	{8'd208,8'd145} : s = 99;
	{8'd208,8'd146} : s = 92;
	{8'd208,8'd147} : s = 218;
	{8'd208,8'd148} : s = 90;
	{8'd208,8'd149} : s = 217;
	{8'd208,8'd150} : s = 214;
	{8'd208,8'd151} : s = 373;
	{8'd208,8'd152} : s = 89;
	{8'd208,8'd153} : s = 213;
	{8'd208,8'd154} : s = 211;
	{8'd208,8'd155} : s = 371;
	{8'd208,8'd156} : s = 206;
	{8'd208,8'd157} : s = 366;
	{8'd208,8'd158} : s = 365;
	{8'd208,8'd159} : s = 478;
	{8'd208,8'd160} : s = 86;
	{8'd208,8'd161} : s = 205;
	{8'd208,8'd162} : s = 203;
	{8'd208,8'd163} : s = 363;
	{8'd208,8'd164} : s = 199;
	{8'd208,8'd165} : s = 359;
	{8'd208,8'd166} : s = 350;
	{8'd208,8'd167} : s = 477;
	{8'd208,8'd168} : s = 188;
	{8'd208,8'd169} : s = 349;
	{8'd208,8'd170} : s = 347;
	{8'd208,8'd171} : s = 475;
	{8'd208,8'd172} : s = 343;
	{8'd208,8'd173} : s = 471;
	{8'd208,8'd174} : s = 463;
	{8'd208,8'd175} : s = 509;
	{8'd208,8'd176} : s = 3;
	{8'd208,8'd177} : s = 22;
	{8'd208,8'd178} : s = 21;
	{8'd208,8'd179} : s = 85;
	{8'd208,8'd180} : s = 19;
	{8'd208,8'd181} : s = 83;
	{8'd208,8'd182} : s = 78;
	{8'd208,8'd183} : s = 186;
	{8'd208,8'd184} : s = 14;
	{8'd208,8'd185} : s = 77;
	{8'd208,8'd186} : s = 75;
	{8'd208,8'd187} : s = 185;
	{8'd208,8'd188} : s = 71;
	{8'd208,8'd189} : s = 182;
	{8'd208,8'd190} : s = 181;
	{8'd208,8'd191} : s = 335;
	{8'd208,8'd192} : s = 13;
	{8'd208,8'd193} : s = 60;
	{8'd208,8'd194} : s = 58;
	{8'd208,8'd195} : s = 179;
	{8'd208,8'd196} : s = 57;
	{8'd208,8'd197} : s = 174;
	{8'd208,8'd198} : s = 173;
	{8'd208,8'd199} : s = 318;
	{8'd208,8'd200} : s = 54;
	{8'd208,8'd201} : s = 171;
	{8'd208,8'd202} : s = 167;
	{8'd208,8'd203} : s = 317;
	{8'd208,8'd204} : s = 158;
	{8'd208,8'd205} : s = 315;
	{8'd208,8'd206} : s = 311;
	{8'd208,8'd207} : s = 446;
	{8'd208,8'd208} : s = 11;
	{8'd208,8'd209} : s = 53;
	{8'd208,8'd210} : s = 51;
	{8'd208,8'd211} : s = 157;
	{8'd208,8'd212} : s = 46;
	{8'd208,8'd213} : s = 155;
	{8'd208,8'd214} : s = 151;
	{8'd208,8'd215} : s = 303;
	{8'd208,8'd216} : s = 45;
	{8'd208,8'd217} : s = 143;
	{8'd208,8'd218} : s = 124;
	{8'd208,8'd219} : s = 287;
	{8'd208,8'd220} : s = 122;
	{8'd208,8'd221} : s = 252;
	{8'd208,8'd222} : s = 250;
	{8'd208,8'd223} : s = 445;
	{8'd208,8'd224} : s = 43;
	{8'd208,8'd225} : s = 121;
	{8'd208,8'd226} : s = 118;
	{8'd208,8'd227} : s = 249;
	{8'd208,8'd228} : s = 117;
	{8'd208,8'd229} : s = 246;
	{8'd208,8'd230} : s = 245;
	{8'd208,8'd231} : s = 443;
	{8'd208,8'd232} : s = 115;
	{8'd208,8'd233} : s = 243;
	{8'd208,8'd234} : s = 238;
	{8'd208,8'd235} : s = 439;
	{8'd208,8'd236} : s = 237;
	{8'd208,8'd237} : s = 431;
	{8'd208,8'd238} : s = 415;
	{8'd208,8'd239} : s = 507;
	{8'd208,8'd240} : s = 7;
	{8'd208,8'd241} : s = 39;
	{8'd208,8'd242} : s = 30;
	{8'd208,8'd243} : s = 110;
	{8'd208,8'd244} : s = 29;
	{8'd208,8'd245} : s = 109;
	{8'd208,8'd246} : s = 107;
	{8'd208,8'd247} : s = 235;
	{8'd208,8'd248} : s = 27;
	{8'd208,8'd249} : s = 103;
	{8'd208,8'd250} : s = 94;
	{8'd208,8'd251} : s = 231;
	{8'd208,8'd252} : s = 93;
	{8'd208,8'd253} : s = 222;
	{8'd208,8'd254} : s = 221;
	{8'd208,8'd255} : s = 382;
	{8'd209,8'd0} : s = 216;
	{8'd209,8'd1} : s = 212;
	{8'd209,8'd2} : s = 362;
	{8'd209,8'd3} : s = 210;
	{8'd209,8'd4} : s = 361;
	{8'd209,8'd5} : s = 358;
	{8'd209,8'd6} : s = 469;
	{8'd209,8'd7} : s = 209;
	{8'd209,8'd8} : s = 357;
	{8'd209,8'd9} : s = 355;
	{8'd209,8'd10} : s = 467;
	{8'd209,8'd11} : s = 348;
	{8'd209,8'd12} : s = 462;
	{8'd209,8'd13} : s = 461;
	{8'd209,8'd14} : s = 505;
	{8'd209,8'd15} : s = 84;
	{8'd209,8'd16} : s = 204;
	{8'd209,8'd17} : s = 202;
	{8'd209,8'd18} : s = 346;
	{8'd209,8'd19} : s = 201;
	{8'd209,8'd20} : s = 345;
	{8'd209,8'd21} : s = 342;
	{8'd209,8'd22} : s = 459;
	{8'd209,8'd23} : s = 198;
	{8'd209,8'd24} : s = 341;
	{8'd209,8'd25} : s = 339;
	{8'd209,8'd26} : s = 455;
	{8'd209,8'd27} : s = 334;
	{8'd209,8'd28} : s = 444;
	{8'd209,8'd29} : s = 442;
	{8'd209,8'd30} : s = 502;
	{8'd209,8'd31} : s = 197;
	{8'd209,8'd32} : s = 333;
	{8'd209,8'd33} : s = 331;
	{8'd209,8'd34} : s = 441;
	{8'd209,8'd35} : s = 327;
	{8'd209,8'd36} : s = 438;
	{8'd209,8'd37} : s = 437;
	{8'd209,8'd38} : s = 501;
	{8'd209,8'd39} : s = 316;
	{8'd209,8'd40} : s = 435;
	{8'd209,8'd41} : s = 430;
	{8'd209,8'd42} : s = 499;
	{8'd209,8'd43} : s = 429;
	{8'd209,8'd44} : s = 494;
	{8'd209,8'd45} : s = 493;
	{8'd209,8'd46} : s = 510;
	{8'd209,8'd47} : s = 1;
	{8'd209,8'd48} : s = 18;
	{8'd209,8'd49} : s = 17;
	{8'd209,8'd50} : s = 82;
	{8'd209,8'd51} : s = 12;
	{8'd209,8'd52} : s = 81;
	{8'd209,8'd53} : s = 76;
	{8'd209,8'd54} : s = 195;
	{8'd209,8'd55} : s = 10;
	{8'd209,8'd56} : s = 74;
	{8'd209,8'd57} : s = 73;
	{8'd209,8'd58} : s = 184;
	{8'd209,8'd59} : s = 70;
	{8'd209,8'd60} : s = 180;
	{8'd209,8'd61} : s = 178;
	{8'd209,8'd62} : s = 314;
	{8'd209,8'd63} : s = 9;
	{8'd209,8'd64} : s = 69;
	{8'd209,8'd65} : s = 67;
	{8'd209,8'd66} : s = 177;
	{8'd209,8'd67} : s = 56;
	{8'd209,8'd68} : s = 172;
	{8'd209,8'd69} : s = 170;
	{8'd209,8'd70} : s = 313;
	{8'd209,8'd71} : s = 52;
	{8'd209,8'd72} : s = 169;
	{8'd209,8'd73} : s = 166;
	{8'd209,8'd74} : s = 310;
	{8'd209,8'd75} : s = 165;
	{8'd209,8'd76} : s = 309;
	{8'd209,8'd77} : s = 307;
	{8'd209,8'd78} : s = 427;
	{8'd209,8'd79} : s = 6;
	{8'd209,8'd80} : s = 50;
	{8'd209,8'd81} : s = 49;
	{8'd209,8'd82} : s = 163;
	{8'd209,8'd83} : s = 44;
	{8'd209,8'd84} : s = 156;
	{8'd209,8'd85} : s = 154;
	{8'd209,8'd86} : s = 302;
	{8'd209,8'd87} : s = 42;
	{8'd209,8'd88} : s = 153;
	{8'd209,8'd89} : s = 150;
	{8'd209,8'd90} : s = 301;
	{8'd209,8'd91} : s = 149;
	{8'd209,8'd92} : s = 299;
	{8'd209,8'd93} : s = 295;
	{8'd209,8'd94} : s = 423;
	{8'd209,8'd95} : s = 41;
	{8'd209,8'd96} : s = 147;
	{8'd209,8'd97} : s = 142;
	{8'd209,8'd98} : s = 286;
	{8'd209,8'd99} : s = 141;
	{8'd209,8'd100} : s = 285;
	{8'd209,8'd101} : s = 283;
	{8'd209,8'd102} : s = 414;
	{8'd209,8'd103} : s = 139;
	{8'd209,8'd104} : s = 279;
	{8'd209,8'd105} : s = 271;
	{8'd209,8'd106} : s = 413;
	{8'd209,8'd107} : s = 248;
	{8'd209,8'd108} : s = 411;
	{8'd209,8'd109} : s = 407;
	{8'd209,8'd110} : s = 491;
	{8'd209,8'd111} : s = 5;
	{8'd209,8'd112} : s = 38;
	{8'd209,8'd113} : s = 37;
	{8'd209,8'd114} : s = 135;
	{8'd209,8'd115} : s = 35;
	{8'd209,8'd116} : s = 120;
	{8'd209,8'd117} : s = 116;
	{8'd209,8'd118} : s = 244;
	{8'd209,8'd119} : s = 28;
	{8'd209,8'd120} : s = 114;
	{8'd209,8'd121} : s = 113;
	{8'd209,8'd122} : s = 242;
	{8'd209,8'd123} : s = 108;
	{8'd209,8'd124} : s = 241;
	{8'd209,8'd125} : s = 236;
	{8'd209,8'd126} : s = 399;
	{8'd209,8'd127} : s = 26;
	{8'd209,8'd128} : s = 106;
	{8'd209,8'd129} : s = 105;
	{8'd209,8'd130} : s = 234;
	{8'd209,8'd131} : s = 102;
	{8'd209,8'd132} : s = 233;
	{8'd209,8'd133} : s = 230;
	{8'd209,8'd134} : s = 380;
	{8'd209,8'd135} : s = 101;
	{8'd209,8'd136} : s = 229;
	{8'd209,8'd137} : s = 227;
	{8'd209,8'd138} : s = 378;
	{8'd209,8'd139} : s = 220;
	{8'd209,8'd140} : s = 377;
	{8'd209,8'd141} : s = 374;
	{8'd209,8'd142} : s = 487;
	{8'd209,8'd143} : s = 25;
	{8'd209,8'd144} : s = 99;
	{8'd209,8'd145} : s = 92;
	{8'd209,8'd146} : s = 218;
	{8'd209,8'd147} : s = 90;
	{8'd209,8'd148} : s = 217;
	{8'd209,8'd149} : s = 214;
	{8'd209,8'd150} : s = 373;
	{8'd209,8'd151} : s = 89;
	{8'd209,8'd152} : s = 213;
	{8'd209,8'd153} : s = 211;
	{8'd209,8'd154} : s = 371;
	{8'd209,8'd155} : s = 206;
	{8'd209,8'd156} : s = 366;
	{8'd209,8'd157} : s = 365;
	{8'd209,8'd158} : s = 478;
	{8'd209,8'd159} : s = 86;
	{8'd209,8'd160} : s = 205;
	{8'd209,8'd161} : s = 203;
	{8'd209,8'd162} : s = 363;
	{8'd209,8'd163} : s = 199;
	{8'd209,8'd164} : s = 359;
	{8'd209,8'd165} : s = 350;
	{8'd209,8'd166} : s = 477;
	{8'd209,8'd167} : s = 188;
	{8'd209,8'd168} : s = 349;
	{8'd209,8'd169} : s = 347;
	{8'd209,8'd170} : s = 475;
	{8'd209,8'd171} : s = 343;
	{8'd209,8'd172} : s = 471;
	{8'd209,8'd173} : s = 463;
	{8'd209,8'd174} : s = 509;
	{8'd209,8'd175} : s = 3;
	{8'd209,8'd176} : s = 22;
	{8'd209,8'd177} : s = 21;
	{8'd209,8'd178} : s = 85;
	{8'd209,8'd179} : s = 19;
	{8'd209,8'd180} : s = 83;
	{8'd209,8'd181} : s = 78;
	{8'd209,8'd182} : s = 186;
	{8'd209,8'd183} : s = 14;
	{8'd209,8'd184} : s = 77;
	{8'd209,8'd185} : s = 75;
	{8'd209,8'd186} : s = 185;
	{8'd209,8'd187} : s = 71;
	{8'd209,8'd188} : s = 182;
	{8'd209,8'd189} : s = 181;
	{8'd209,8'd190} : s = 335;
	{8'd209,8'd191} : s = 13;
	{8'd209,8'd192} : s = 60;
	{8'd209,8'd193} : s = 58;
	{8'd209,8'd194} : s = 179;
	{8'd209,8'd195} : s = 57;
	{8'd209,8'd196} : s = 174;
	{8'd209,8'd197} : s = 173;
	{8'd209,8'd198} : s = 318;
	{8'd209,8'd199} : s = 54;
	{8'd209,8'd200} : s = 171;
	{8'd209,8'd201} : s = 167;
	{8'd209,8'd202} : s = 317;
	{8'd209,8'd203} : s = 158;
	{8'd209,8'd204} : s = 315;
	{8'd209,8'd205} : s = 311;
	{8'd209,8'd206} : s = 446;
	{8'd209,8'd207} : s = 11;
	{8'd209,8'd208} : s = 53;
	{8'd209,8'd209} : s = 51;
	{8'd209,8'd210} : s = 157;
	{8'd209,8'd211} : s = 46;
	{8'd209,8'd212} : s = 155;
	{8'd209,8'd213} : s = 151;
	{8'd209,8'd214} : s = 303;
	{8'd209,8'd215} : s = 45;
	{8'd209,8'd216} : s = 143;
	{8'd209,8'd217} : s = 124;
	{8'd209,8'd218} : s = 287;
	{8'd209,8'd219} : s = 122;
	{8'd209,8'd220} : s = 252;
	{8'd209,8'd221} : s = 250;
	{8'd209,8'd222} : s = 445;
	{8'd209,8'd223} : s = 43;
	{8'd209,8'd224} : s = 121;
	{8'd209,8'd225} : s = 118;
	{8'd209,8'd226} : s = 249;
	{8'd209,8'd227} : s = 117;
	{8'd209,8'd228} : s = 246;
	{8'd209,8'd229} : s = 245;
	{8'd209,8'd230} : s = 443;
	{8'd209,8'd231} : s = 115;
	{8'd209,8'd232} : s = 243;
	{8'd209,8'd233} : s = 238;
	{8'd209,8'd234} : s = 439;
	{8'd209,8'd235} : s = 237;
	{8'd209,8'd236} : s = 431;
	{8'd209,8'd237} : s = 415;
	{8'd209,8'd238} : s = 507;
	{8'd209,8'd239} : s = 7;
	{8'd209,8'd240} : s = 39;
	{8'd209,8'd241} : s = 30;
	{8'd209,8'd242} : s = 110;
	{8'd209,8'd243} : s = 29;
	{8'd209,8'd244} : s = 109;
	{8'd209,8'd245} : s = 107;
	{8'd209,8'd246} : s = 235;
	{8'd209,8'd247} : s = 27;
	{8'd209,8'd248} : s = 103;
	{8'd209,8'd249} : s = 94;
	{8'd209,8'd250} : s = 231;
	{8'd209,8'd251} : s = 93;
	{8'd209,8'd252} : s = 222;
	{8'd209,8'd253} : s = 221;
	{8'd209,8'd254} : s = 382;
	{8'd209,8'd255} : s = 23;
	{8'd210,8'd0} : s = 212;
	{8'd210,8'd1} : s = 362;
	{8'd210,8'd2} : s = 210;
	{8'd210,8'd3} : s = 361;
	{8'd210,8'd4} : s = 358;
	{8'd210,8'd5} : s = 469;
	{8'd210,8'd6} : s = 209;
	{8'd210,8'd7} : s = 357;
	{8'd210,8'd8} : s = 355;
	{8'd210,8'd9} : s = 467;
	{8'd210,8'd10} : s = 348;
	{8'd210,8'd11} : s = 462;
	{8'd210,8'd12} : s = 461;
	{8'd210,8'd13} : s = 505;
	{8'd210,8'd14} : s = 84;
	{8'd210,8'd15} : s = 204;
	{8'd210,8'd16} : s = 202;
	{8'd210,8'd17} : s = 346;
	{8'd210,8'd18} : s = 201;
	{8'd210,8'd19} : s = 345;
	{8'd210,8'd20} : s = 342;
	{8'd210,8'd21} : s = 459;
	{8'd210,8'd22} : s = 198;
	{8'd210,8'd23} : s = 341;
	{8'd210,8'd24} : s = 339;
	{8'd210,8'd25} : s = 455;
	{8'd210,8'd26} : s = 334;
	{8'd210,8'd27} : s = 444;
	{8'd210,8'd28} : s = 442;
	{8'd210,8'd29} : s = 502;
	{8'd210,8'd30} : s = 197;
	{8'd210,8'd31} : s = 333;
	{8'd210,8'd32} : s = 331;
	{8'd210,8'd33} : s = 441;
	{8'd210,8'd34} : s = 327;
	{8'd210,8'd35} : s = 438;
	{8'd210,8'd36} : s = 437;
	{8'd210,8'd37} : s = 501;
	{8'd210,8'd38} : s = 316;
	{8'd210,8'd39} : s = 435;
	{8'd210,8'd40} : s = 430;
	{8'd210,8'd41} : s = 499;
	{8'd210,8'd42} : s = 429;
	{8'd210,8'd43} : s = 494;
	{8'd210,8'd44} : s = 493;
	{8'd210,8'd45} : s = 510;
	{8'd210,8'd46} : s = 1;
	{8'd210,8'd47} : s = 18;
	{8'd210,8'd48} : s = 17;
	{8'd210,8'd49} : s = 82;
	{8'd210,8'd50} : s = 12;
	{8'd210,8'd51} : s = 81;
	{8'd210,8'd52} : s = 76;
	{8'd210,8'd53} : s = 195;
	{8'd210,8'd54} : s = 10;
	{8'd210,8'd55} : s = 74;
	{8'd210,8'd56} : s = 73;
	{8'd210,8'd57} : s = 184;
	{8'd210,8'd58} : s = 70;
	{8'd210,8'd59} : s = 180;
	{8'd210,8'd60} : s = 178;
	{8'd210,8'd61} : s = 314;
	{8'd210,8'd62} : s = 9;
	{8'd210,8'd63} : s = 69;
	{8'd210,8'd64} : s = 67;
	{8'd210,8'd65} : s = 177;
	{8'd210,8'd66} : s = 56;
	{8'd210,8'd67} : s = 172;
	{8'd210,8'd68} : s = 170;
	{8'd210,8'd69} : s = 313;
	{8'd210,8'd70} : s = 52;
	{8'd210,8'd71} : s = 169;
	{8'd210,8'd72} : s = 166;
	{8'd210,8'd73} : s = 310;
	{8'd210,8'd74} : s = 165;
	{8'd210,8'd75} : s = 309;
	{8'd210,8'd76} : s = 307;
	{8'd210,8'd77} : s = 427;
	{8'd210,8'd78} : s = 6;
	{8'd210,8'd79} : s = 50;
	{8'd210,8'd80} : s = 49;
	{8'd210,8'd81} : s = 163;
	{8'd210,8'd82} : s = 44;
	{8'd210,8'd83} : s = 156;
	{8'd210,8'd84} : s = 154;
	{8'd210,8'd85} : s = 302;
	{8'd210,8'd86} : s = 42;
	{8'd210,8'd87} : s = 153;
	{8'd210,8'd88} : s = 150;
	{8'd210,8'd89} : s = 301;
	{8'd210,8'd90} : s = 149;
	{8'd210,8'd91} : s = 299;
	{8'd210,8'd92} : s = 295;
	{8'd210,8'd93} : s = 423;
	{8'd210,8'd94} : s = 41;
	{8'd210,8'd95} : s = 147;
	{8'd210,8'd96} : s = 142;
	{8'd210,8'd97} : s = 286;
	{8'd210,8'd98} : s = 141;
	{8'd210,8'd99} : s = 285;
	{8'd210,8'd100} : s = 283;
	{8'd210,8'd101} : s = 414;
	{8'd210,8'd102} : s = 139;
	{8'd210,8'd103} : s = 279;
	{8'd210,8'd104} : s = 271;
	{8'd210,8'd105} : s = 413;
	{8'd210,8'd106} : s = 248;
	{8'd210,8'd107} : s = 411;
	{8'd210,8'd108} : s = 407;
	{8'd210,8'd109} : s = 491;
	{8'd210,8'd110} : s = 5;
	{8'd210,8'd111} : s = 38;
	{8'd210,8'd112} : s = 37;
	{8'd210,8'd113} : s = 135;
	{8'd210,8'd114} : s = 35;
	{8'd210,8'd115} : s = 120;
	{8'd210,8'd116} : s = 116;
	{8'd210,8'd117} : s = 244;
	{8'd210,8'd118} : s = 28;
	{8'd210,8'd119} : s = 114;
	{8'd210,8'd120} : s = 113;
	{8'd210,8'd121} : s = 242;
	{8'd210,8'd122} : s = 108;
	{8'd210,8'd123} : s = 241;
	{8'd210,8'd124} : s = 236;
	{8'd210,8'd125} : s = 399;
	{8'd210,8'd126} : s = 26;
	{8'd210,8'd127} : s = 106;
	{8'd210,8'd128} : s = 105;
	{8'd210,8'd129} : s = 234;
	{8'd210,8'd130} : s = 102;
	{8'd210,8'd131} : s = 233;
	{8'd210,8'd132} : s = 230;
	{8'd210,8'd133} : s = 380;
	{8'd210,8'd134} : s = 101;
	{8'd210,8'd135} : s = 229;
	{8'd210,8'd136} : s = 227;
	{8'd210,8'd137} : s = 378;
	{8'd210,8'd138} : s = 220;
	{8'd210,8'd139} : s = 377;
	{8'd210,8'd140} : s = 374;
	{8'd210,8'd141} : s = 487;
	{8'd210,8'd142} : s = 25;
	{8'd210,8'd143} : s = 99;
	{8'd210,8'd144} : s = 92;
	{8'd210,8'd145} : s = 218;
	{8'd210,8'd146} : s = 90;
	{8'd210,8'd147} : s = 217;
	{8'd210,8'd148} : s = 214;
	{8'd210,8'd149} : s = 373;
	{8'd210,8'd150} : s = 89;
	{8'd210,8'd151} : s = 213;
	{8'd210,8'd152} : s = 211;
	{8'd210,8'd153} : s = 371;
	{8'd210,8'd154} : s = 206;
	{8'd210,8'd155} : s = 366;
	{8'd210,8'd156} : s = 365;
	{8'd210,8'd157} : s = 478;
	{8'd210,8'd158} : s = 86;
	{8'd210,8'd159} : s = 205;
	{8'd210,8'd160} : s = 203;
	{8'd210,8'd161} : s = 363;
	{8'd210,8'd162} : s = 199;
	{8'd210,8'd163} : s = 359;
	{8'd210,8'd164} : s = 350;
	{8'd210,8'd165} : s = 477;
	{8'd210,8'd166} : s = 188;
	{8'd210,8'd167} : s = 349;
	{8'd210,8'd168} : s = 347;
	{8'd210,8'd169} : s = 475;
	{8'd210,8'd170} : s = 343;
	{8'd210,8'd171} : s = 471;
	{8'd210,8'd172} : s = 463;
	{8'd210,8'd173} : s = 509;
	{8'd210,8'd174} : s = 3;
	{8'd210,8'd175} : s = 22;
	{8'd210,8'd176} : s = 21;
	{8'd210,8'd177} : s = 85;
	{8'd210,8'd178} : s = 19;
	{8'd210,8'd179} : s = 83;
	{8'd210,8'd180} : s = 78;
	{8'd210,8'd181} : s = 186;
	{8'd210,8'd182} : s = 14;
	{8'd210,8'd183} : s = 77;
	{8'd210,8'd184} : s = 75;
	{8'd210,8'd185} : s = 185;
	{8'd210,8'd186} : s = 71;
	{8'd210,8'd187} : s = 182;
	{8'd210,8'd188} : s = 181;
	{8'd210,8'd189} : s = 335;
	{8'd210,8'd190} : s = 13;
	{8'd210,8'd191} : s = 60;
	{8'd210,8'd192} : s = 58;
	{8'd210,8'd193} : s = 179;
	{8'd210,8'd194} : s = 57;
	{8'd210,8'd195} : s = 174;
	{8'd210,8'd196} : s = 173;
	{8'd210,8'd197} : s = 318;
	{8'd210,8'd198} : s = 54;
	{8'd210,8'd199} : s = 171;
	{8'd210,8'd200} : s = 167;
	{8'd210,8'd201} : s = 317;
	{8'd210,8'd202} : s = 158;
	{8'd210,8'd203} : s = 315;
	{8'd210,8'd204} : s = 311;
	{8'd210,8'd205} : s = 446;
	{8'd210,8'd206} : s = 11;
	{8'd210,8'd207} : s = 53;
	{8'd210,8'd208} : s = 51;
	{8'd210,8'd209} : s = 157;
	{8'd210,8'd210} : s = 46;
	{8'd210,8'd211} : s = 155;
	{8'd210,8'd212} : s = 151;
	{8'd210,8'd213} : s = 303;
	{8'd210,8'd214} : s = 45;
	{8'd210,8'd215} : s = 143;
	{8'd210,8'd216} : s = 124;
	{8'd210,8'd217} : s = 287;
	{8'd210,8'd218} : s = 122;
	{8'd210,8'd219} : s = 252;
	{8'd210,8'd220} : s = 250;
	{8'd210,8'd221} : s = 445;
	{8'd210,8'd222} : s = 43;
	{8'd210,8'd223} : s = 121;
	{8'd210,8'd224} : s = 118;
	{8'd210,8'd225} : s = 249;
	{8'd210,8'd226} : s = 117;
	{8'd210,8'd227} : s = 246;
	{8'd210,8'd228} : s = 245;
	{8'd210,8'd229} : s = 443;
	{8'd210,8'd230} : s = 115;
	{8'd210,8'd231} : s = 243;
	{8'd210,8'd232} : s = 238;
	{8'd210,8'd233} : s = 439;
	{8'd210,8'd234} : s = 237;
	{8'd210,8'd235} : s = 431;
	{8'd210,8'd236} : s = 415;
	{8'd210,8'd237} : s = 507;
	{8'd210,8'd238} : s = 7;
	{8'd210,8'd239} : s = 39;
	{8'd210,8'd240} : s = 30;
	{8'd210,8'd241} : s = 110;
	{8'd210,8'd242} : s = 29;
	{8'd210,8'd243} : s = 109;
	{8'd210,8'd244} : s = 107;
	{8'd210,8'd245} : s = 235;
	{8'd210,8'd246} : s = 27;
	{8'd210,8'd247} : s = 103;
	{8'd210,8'd248} : s = 94;
	{8'd210,8'd249} : s = 231;
	{8'd210,8'd250} : s = 93;
	{8'd210,8'd251} : s = 222;
	{8'd210,8'd252} : s = 221;
	{8'd210,8'd253} : s = 382;
	{8'd210,8'd254} : s = 23;
	{8'd210,8'd255} : s = 91;
	{8'd211,8'd0} : s = 362;
	{8'd211,8'd1} : s = 210;
	{8'd211,8'd2} : s = 361;
	{8'd211,8'd3} : s = 358;
	{8'd211,8'd4} : s = 469;
	{8'd211,8'd5} : s = 209;
	{8'd211,8'd6} : s = 357;
	{8'd211,8'd7} : s = 355;
	{8'd211,8'd8} : s = 467;
	{8'd211,8'd9} : s = 348;
	{8'd211,8'd10} : s = 462;
	{8'd211,8'd11} : s = 461;
	{8'd211,8'd12} : s = 505;
	{8'd211,8'd13} : s = 84;
	{8'd211,8'd14} : s = 204;
	{8'd211,8'd15} : s = 202;
	{8'd211,8'd16} : s = 346;
	{8'd211,8'd17} : s = 201;
	{8'd211,8'd18} : s = 345;
	{8'd211,8'd19} : s = 342;
	{8'd211,8'd20} : s = 459;
	{8'd211,8'd21} : s = 198;
	{8'd211,8'd22} : s = 341;
	{8'd211,8'd23} : s = 339;
	{8'd211,8'd24} : s = 455;
	{8'd211,8'd25} : s = 334;
	{8'd211,8'd26} : s = 444;
	{8'd211,8'd27} : s = 442;
	{8'd211,8'd28} : s = 502;
	{8'd211,8'd29} : s = 197;
	{8'd211,8'd30} : s = 333;
	{8'd211,8'd31} : s = 331;
	{8'd211,8'd32} : s = 441;
	{8'd211,8'd33} : s = 327;
	{8'd211,8'd34} : s = 438;
	{8'd211,8'd35} : s = 437;
	{8'd211,8'd36} : s = 501;
	{8'd211,8'd37} : s = 316;
	{8'd211,8'd38} : s = 435;
	{8'd211,8'd39} : s = 430;
	{8'd211,8'd40} : s = 499;
	{8'd211,8'd41} : s = 429;
	{8'd211,8'd42} : s = 494;
	{8'd211,8'd43} : s = 493;
	{8'd211,8'd44} : s = 510;
	{8'd211,8'd45} : s = 1;
	{8'd211,8'd46} : s = 18;
	{8'd211,8'd47} : s = 17;
	{8'd211,8'd48} : s = 82;
	{8'd211,8'd49} : s = 12;
	{8'd211,8'd50} : s = 81;
	{8'd211,8'd51} : s = 76;
	{8'd211,8'd52} : s = 195;
	{8'd211,8'd53} : s = 10;
	{8'd211,8'd54} : s = 74;
	{8'd211,8'd55} : s = 73;
	{8'd211,8'd56} : s = 184;
	{8'd211,8'd57} : s = 70;
	{8'd211,8'd58} : s = 180;
	{8'd211,8'd59} : s = 178;
	{8'd211,8'd60} : s = 314;
	{8'd211,8'd61} : s = 9;
	{8'd211,8'd62} : s = 69;
	{8'd211,8'd63} : s = 67;
	{8'd211,8'd64} : s = 177;
	{8'd211,8'd65} : s = 56;
	{8'd211,8'd66} : s = 172;
	{8'd211,8'd67} : s = 170;
	{8'd211,8'd68} : s = 313;
	{8'd211,8'd69} : s = 52;
	{8'd211,8'd70} : s = 169;
	{8'd211,8'd71} : s = 166;
	{8'd211,8'd72} : s = 310;
	{8'd211,8'd73} : s = 165;
	{8'd211,8'd74} : s = 309;
	{8'd211,8'd75} : s = 307;
	{8'd211,8'd76} : s = 427;
	{8'd211,8'd77} : s = 6;
	{8'd211,8'd78} : s = 50;
	{8'd211,8'd79} : s = 49;
	{8'd211,8'd80} : s = 163;
	{8'd211,8'd81} : s = 44;
	{8'd211,8'd82} : s = 156;
	{8'd211,8'd83} : s = 154;
	{8'd211,8'd84} : s = 302;
	{8'd211,8'd85} : s = 42;
	{8'd211,8'd86} : s = 153;
	{8'd211,8'd87} : s = 150;
	{8'd211,8'd88} : s = 301;
	{8'd211,8'd89} : s = 149;
	{8'd211,8'd90} : s = 299;
	{8'd211,8'd91} : s = 295;
	{8'd211,8'd92} : s = 423;
	{8'd211,8'd93} : s = 41;
	{8'd211,8'd94} : s = 147;
	{8'd211,8'd95} : s = 142;
	{8'd211,8'd96} : s = 286;
	{8'd211,8'd97} : s = 141;
	{8'd211,8'd98} : s = 285;
	{8'd211,8'd99} : s = 283;
	{8'd211,8'd100} : s = 414;
	{8'd211,8'd101} : s = 139;
	{8'd211,8'd102} : s = 279;
	{8'd211,8'd103} : s = 271;
	{8'd211,8'd104} : s = 413;
	{8'd211,8'd105} : s = 248;
	{8'd211,8'd106} : s = 411;
	{8'd211,8'd107} : s = 407;
	{8'd211,8'd108} : s = 491;
	{8'd211,8'd109} : s = 5;
	{8'd211,8'd110} : s = 38;
	{8'd211,8'd111} : s = 37;
	{8'd211,8'd112} : s = 135;
	{8'd211,8'd113} : s = 35;
	{8'd211,8'd114} : s = 120;
	{8'd211,8'd115} : s = 116;
	{8'd211,8'd116} : s = 244;
	{8'd211,8'd117} : s = 28;
	{8'd211,8'd118} : s = 114;
	{8'd211,8'd119} : s = 113;
	{8'd211,8'd120} : s = 242;
	{8'd211,8'd121} : s = 108;
	{8'd211,8'd122} : s = 241;
	{8'd211,8'd123} : s = 236;
	{8'd211,8'd124} : s = 399;
	{8'd211,8'd125} : s = 26;
	{8'd211,8'd126} : s = 106;
	{8'd211,8'd127} : s = 105;
	{8'd211,8'd128} : s = 234;
	{8'd211,8'd129} : s = 102;
	{8'd211,8'd130} : s = 233;
	{8'd211,8'd131} : s = 230;
	{8'd211,8'd132} : s = 380;
	{8'd211,8'd133} : s = 101;
	{8'd211,8'd134} : s = 229;
	{8'd211,8'd135} : s = 227;
	{8'd211,8'd136} : s = 378;
	{8'd211,8'd137} : s = 220;
	{8'd211,8'd138} : s = 377;
	{8'd211,8'd139} : s = 374;
	{8'd211,8'd140} : s = 487;
	{8'd211,8'd141} : s = 25;
	{8'd211,8'd142} : s = 99;
	{8'd211,8'd143} : s = 92;
	{8'd211,8'd144} : s = 218;
	{8'd211,8'd145} : s = 90;
	{8'd211,8'd146} : s = 217;
	{8'd211,8'd147} : s = 214;
	{8'd211,8'd148} : s = 373;
	{8'd211,8'd149} : s = 89;
	{8'd211,8'd150} : s = 213;
	{8'd211,8'd151} : s = 211;
	{8'd211,8'd152} : s = 371;
	{8'd211,8'd153} : s = 206;
	{8'd211,8'd154} : s = 366;
	{8'd211,8'd155} : s = 365;
	{8'd211,8'd156} : s = 478;
	{8'd211,8'd157} : s = 86;
	{8'd211,8'd158} : s = 205;
	{8'd211,8'd159} : s = 203;
	{8'd211,8'd160} : s = 363;
	{8'd211,8'd161} : s = 199;
	{8'd211,8'd162} : s = 359;
	{8'd211,8'd163} : s = 350;
	{8'd211,8'd164} : s = 477;
	{8'd211,8'd165} : s = 188;
	{8'd211,8'd166} : s = 349;
	{8'd211,8'd167} : s = 347;
	{8'd211,8'd168} : s = 475;
	{8'd211,8'd169} : s = 343;
	{8'd211,8'd170} : s = 471;
	{8'd211,8'd171} : s = 463;
	{8'd211,8'd172} : s = 509;
	{8'd211,8'd173} : s = 3;
	{8'd211,8'd174} : s = 22;
	{8'd211,8'd175} : s = 21;
	{8'd211,8'd176} : s = 85;
	{8'd211,8'd177} : s = 19;
	{8'd211,8'd178} : s = 83;
	{8'd211,8'd179} : s = 78;
	{8'd211,8'd180} : s = 186;
	{8'd211,8'd181} : s = 14;
	{8'd211,8'd182} : s = 77;
	{8'd211,8'd183} : s = 75;
	{8'd211,8'd184} : s = 185;
	{8'd211,8'd185} : s = 71;
	{8'd211,8'd186} : s = 182;
	{8'd211,8'd187} : s = 181;
	{8'd211,8'd188} : s = 335;
	{8'd211,8'd189} : s = 13;
	{8'd211,8'd190} : s = 60;
	{8'd211,8'd191} : s = 58;
	{8'd211,8'd192} : s = 179;
	{8'd211,8'd193} : s = 57;
	{8'd211,8'd194} : s = 174;
	{8'd211,8'd195} : s = 173;
	{8'd211,8'd196} : s = 318;
	{8'd211,8'd197} : s = 54;
	{8'd211,8'd198} : s = 171;
	{8'd211,8'd199} : s = 167;
	{8'd211,8'd200} : s = 317;
	{8'd211,8'd201} : s = 158;
	{8'd211,8'd202} : s = 315;
	{8'd211,8'd203} : s = 311;
	{8'd211,8'd204} : s = 446;
	{8'd211,8'd205} : s = 11;
	{8'd211,8'd206} : s = 53;
	{8'd211,8'd207} : s = 51;
	{8'd211,8'd208} : s = 157;
	{8'd211,8'd209} : s = 46;
	{8'd211,8'd210} : s = 155;
	{8'd211,8'd211} : s = 151;
	{8'd211,8'd212} : s = 303;
	{8'd211,8'd213} : s = 45;
	{8'd211,8'd214} : s = 143;
	{8'd211,8'd215} : s = 124;
	{8'd211,8'd216} : s = 287;
	{8'd211,8'd217} : s = 122;
	{8'd211,8'd218} : s = 252;
	{8'd211,8'd219} : s = 250;
	{8'd211,8'd220} : s = 445;
	{8'd211,8'd221} : s = 43;
	{8'd211,8'd222} : s = 121;
	{8'd211,8'd223} : s = 118;
	{8'd211,8'd224} : s = 249;
	{8'd211,8'd225} : s = 117;
	{8'd211,8'd226} : s = 246;
	{8'd211,8'd227} : s = 245;
	{8'd211,8'd228} : s = 443;
	{8'd211,8'd229} : s = 115;
	{8'd211,8'd230} : s = 243;
	{8'd211,8'd231} : s = 238;
	{8'd211,8'd232} : s = 439;
	{8'd211,8'd233} : s = 237;
	{8'd211,8'd234} : s = 431;
	{8'd211,8'd235} : s = 415;
	{8'd211,8'd236} : s = 507;
	{8'd211,8'd237} : s = 7;
	{8'd211,8'd238} : s = 39;
	{8'd211,8'd239} : s = 30;
	{8'd211,8'd240} : s = 110;
	{8'd211,8'd241} : s = 29;
	{8'd211,8'd242} : s = 109;
	{8'd211,8'd243} : s = 107;
	{8'd211,8'd244} : s = 235;
	{8'd211,8'd245} : s = 27;
	{8'd211,8'd246} : s = 103;
	{8'd211,8'd247} : s = 94;
	{8'd211,8'd248} : s = 231;
	{8'd211,8'd249} : s = 93;
	{8'd211,8'd250} : s = 222;
	{8'd211,8'd251} : s = 221;
	{8'd211,8'd252} : s = 382;
	{8'd211,8'd253} : s = 23;
	{8'd211,8'd254} : s = 91;
	{8'd211,8'd255} : s = 87;
	{8'd212,8'd0} : s = 210;
	{8'd212,8'd1} : s = 361;
	{8'd212,8'd2} : s = 358;
	{8'd212,8'd3} : s = 469;
	{8'd212,8'd4} : s = 209;
	{8'd212,8'd5} : s = 357;
	{8'd212,8'd6} : s = 355;
	{8'd212,8'd7} : s = 467;
	{8'd212,8'd8} : s = 348;
	{8'd212,8'd9} : s = 462;
	{8'd212,8'd10} : s = 461;
	{8'd212,8'd11} : s = 505;
	{8'd212,8'd12} : s = 84;
	{8'd212,8'd13} : s = 204;
	{8'd212,8'd14} : s = 202;
	{8'd212,8'd15} : s = 346;
	{8'd212,8'd16} : s = 201;
	{8'd212,8'd17} : s = 345;
	{8'd212,8'd18} : s = 342;
	{8'd212,8'd19} : s = 459;
	{8'd212,8'd20} : s = 198;
	{8'd212,8'd21} : s = 341;
	{8'd212,8'd22} : s = 339;
	{8'd212,8'd23} : s = 455;
	{8'd212,8'd24} : s = 334;
	{8'd212,8'd25} : s = 444;
	{8'd212,8'd26} : s = 442;
	{8'd212,8'd27} : s = 502;
	{8'd212,8'd28} : s = 197;
	{8'd212,8'd29} : s = 333;
	{8'd212,8'd30} : s = 331;
	{8'd212,8'd31} : s = 441;
	{8'd212,8'd32} : s = 327;
	{8'd212,8'd33} : s = 438;
	{8'd212,8'd34} : s = 437;
	{8'd212,8'd35} : s = 501;
	{8'd212,8'd36} : s = 316;
	{8'd212,8'd37} : s = 435;
	{8'd212,8'd38} : s = 430;
	{8'd212,8'd39} : s = 499;
	{8'd212,8'd40} : s = 429;
	{8'd212,8'd41} : s = 494;
	{8'd212,8'd42} : s = 493;
	{8'd212,8'd43} : s = 510;
	{8'd212,8'd44} : s = 1;
	{8'd212,8'd45} : s = 18;
	{8'd212,8'd46} : s = 17;
	{8'd212,8'd47} : s = 82;
	{8'd212,8'd48} : s = 12;
	{8'd212,8'd49} : s = 81;
	{8'd212,8'd50} : s = 76;
	{8'd212,8'd51} : s = 195;
	{8'd212,8'd52} : s = 10;
	{8'd212,8'd53} : s = 74;
	{8'd212,8'd54} : s = 73;
	{8'd212,8'd55} : s = 184;
	{8'd212,8'd56} : s = 70;
	{8'd212,8'd57} : s = 180;
	{8'd212,8'd58} : s = 178;
	{8'd212,8'd59} : s = 314;
	{8'd212,8'd60} : s = 9;
	{8'd212,8'd61} : s = 69;
	{8'd212,8'd62} : s = 67;
	{8'd212,8'd63} : s = 177;
	{8'd212,8'd64} : s = 56;
	{8'd212,8'd65} : s = 172;
	{8'd212,8'd66} : s = 170;
	{8'd212,8'd67} : s = 313;
	{8'd212,8'd68} : s = 52;
	{8'd212,8'd69} : s = 169;
	{8'd212,8'd70} : s = 166;
	{8'd212,8'd71} : s = 310;
	{8'd212,8'd72} : s = 165;
	{8'd212,8'd73} : s = 309;
	{8'd212,8'd74} : s = 307;
	{8'd212,8'd75} : s = 427;
	{8'd212,8'd76} : s = 6;
	{8'd212,8'd77} : s = 50;
	{8'd212,8'd78} : s = 49;
	{8'd212,8'd79} : s = 163;
	{8'd212,8'd80} : s = 44;
	{8'd212,8'd81} : s = 156;
	{8'd212,8'd82} : s = 154;
	{8'd212,8'd83} : s = 302;
	{8'd212,8'd84} : s = 42;
	{8'd212,8'd85} : s = 153;
	{8'd212,8'd86} : s = 150;
	{8'd212,8'd87} : s = 301;
	{8'd212,8'd88} : s = 149;
	{8'd212,8'd89} : s = 299;
	{8'd212,8'd90} : s = 295;
	{8'd212,8'd91} : s = 423;
	{8'd212,8'd92} : s = 41;
	{8'd212,8'd93} : s = 147;
	{8'd212,8'd94} : s = 142;
	{8'd212,8'd95} : s = 286;
	{8'd212,8'd96} : s = 141;
	{8'd212,8'd97} : s = 285;
	{8'd212,8'd98} : s = 283;
	{8'd212,8'd99} : s = 414;
	{8'd212,8'd100} : s = 139;
	{8'd212,8'd101} : s = 279;
	{8'd212,8'd102} : s = 271;
	{8'd212,8'd103} : s = 413;
	{8'd212,8'd104} : s = 248;
	{8'd212,8'd105} : s = 411;
	{8'd212,8'd106} : s = 407;
	{8'd212,8'd107} : s = 491;
	{8'd212,8'd108} : s = 5;
	{8'd212,8'd109} : s = 38;
	{8'd212,8'd110} : s = 37;
	{8'd212,8'd111} : s = 135;
	{8'd212,8'd112} : s = 35;
	{8'd212,8'd113} : s = 120;
	{8'd212,8'd114} : s = 116;
	{8'd212,8'd115} : s = 244;
	{8'd212,8'd116} : s = 28;
	{8'd212,8'd117} : s = 114;
	{8'd212,8'd118} : s = 113;
	{8'd212,8'd119} : s = 242;
	{8'd212,8'd120} : s = 108;
	{8'd212,8'd121} : s = 241;
	{8'd212,8'd122} : s = 236;
	{8'd212,8'd123} : s = 399;
	{8'd212,8'd124} : s = 26;
	{8'd212,8'd125} : s = 106;
	{8'd212,8'd126} : s = 105;
	{8'd212,8'd127} : s = 234;
	{8'd212,8'd128} : s = 102;
	{8'd212,8'd129} : s = 233;
	{8'd212,8'd130} : s = 230;
	{8'd212,8'd131} : s = 380;
	{8'd212,8'd132} : s = 101;
	{8'd212,8'd133} : s = 229;
	{8'd212,8'd134} : s = 227;
	{8'd212,8'd135} : s = 378;
	{8'd212,8'd136} : s = 220;
	{8'd212,8'd137} : s = 377;
	{8'd212,8'd138} : s = 374;
	{8'd212,8'd139} : s = 487;
	{8'd212,8'd140} : s = 25;
	{8'd212,8'd141} : s = 99;
	{8'd212,8'd142} : s = 92;
	{8'd212,8'd143} : s = 218;
	{8'd212,8'd144} : s = 90;
	{8'd212,8'd145} : s = 217;
	{8'd212,8'd146} : s = 214;
	{8'd212,8'd147} : s = 373;
	{8'd212,8'd148} : s = 89;
	{8'd212,8'd149} : s = 213;
	{8'd212,8'd150} : s = 211;
	{8'd212,8'd151} : s = 371;
	{8'd212,8'd152} : s = 206;
	{8'd212,8'd153} : s = 366;
	{8'd212,8'd154} : s = 365;
	{8'd212,8'd155} : s = 478;
	{8'd212,8'd156} : s = 86;
	{8'd212,8'd157} : s = 205;
	{8'd212,8'd158} : s = 203;
	{8'd212,8'd159} : s = 363;
	{8'd212,8'd160} : s = 199;
	{8'd212,8'd161} : s = 359;
	{8'd212,8'd162} : s = 350;
	{8'd212,8'd163} : s = 477;
	{8'd212,8'd164} : s = 188;
	{8'd212,8'd165} : s = 349;
	{8'd212,8'd166} : s = 347;
	{8'd212,8'd167} : s = 475;
	{8'd212,8'd168} : s = 343;
	{8'd212,8'd169} : s = 471;
	{8'd212,8'd170} : s = 463;
	{8'd212,8'd171} : s = 509;
	{8'd212,8'd172} : s = 3;
	{8'd212,8'd173} : s = 22;
	{8'd212,8'd174} : s = 21;
	{8'd212,8'd175} : s = 85;
	{8'd212,8'd176} : s = 19;
	{8'd212,8'd177} : s = 83;
	{8'd212,8'd178} : s = 78;
	{8'd212,8'd179} : s = 186;
	{8'd212,8'd180} : s = 14;
	{8'd212,8'd181} : s = 77;
	{8'd212,8'd182} : s = 75;
	{8'd212,8'd183} : s = 185;
	{8'd212,8'd184} : s = 71;
	{8'd212,8'd185} : s = 182;
	{8'd212,8'd186} : s = 181;
	{8'd212,8'd187} : s = 335;
	{8'd212,8'd188} : s = 13;
	{8'd212,8'd189} : s = 60;
	{8'd212,8'd190} : s = 58;
	{8'd212,8'd191} : s = 179;
	{8'd212,8'd192} : s = 57;
	{8'd212,8'd193} : s = 174;
	{8'd212,8'd194} : s = 173;
	{8'd212,8'd195} : s = 318;
	{8'd212,8'd196} : s = 54;
	{8'd212,8'd197} : s = 171;
	{8'd212,8'd198} : s = 167;
	{8'd212,8'd199} : s = 317;
	{8'd212,8'd200} : s = 158;
	{8'd212,8'd201} : s = 315;
	{8'd212,8'd202} : s = 311;
	{8'd212,8'd203} : s = 446;
	{8'd212,8'd204} : s = 11;
	{8'd212,8'd205} : s = 53;
	{8'd212,8'd206} : s = 51;
	{8'd212,8'd207} : s = 157;
	{8'd212,8'd208} : s = 46;
	{8'd212,8'd209} : s = 155;
	{8'd212,8'd210} : s = 151;
	{8'd212,8'd211} : s = 303;
	{8'd212,8'd212} : s = 45;
	{8'd212,8'd213} : s = 143;
	{8'd212,8'd214} : s = 124;
	{8'd212,8'd215} : s = 287;
	{8'd212,8'd216} : s = 122;
	{8'd212,8'd217} : s = 252;
	{8'd212,8'd218} : s = 250;
	{8'd212,8'd219} : s = 445;
	{8'd212,8'd220} : s = 43;
	{8'd212,8'd221} : s = 121;
	{8'd212,8'd222} : s = 118;
	{8'd212,8'd223} : s = 249;
	{8'd212,8'd224} : s = 117;
	{8'd212,8'd225} : s = 246;
	{8'd212,8'd226} : s = 245;
	{8'd212,8'd227} : s = 443;
	{8'd212,8'd228} : s = 115;
	{8'd212,8'd229} : s = 243;
	{8'd212,8'd230} : s = 238;
	{8'd212,8'd231} : s = 439;
	{8'd212,8'd232} : s = 237;
	{8'd212,8'd233} : s = 431;
	{8'd212,8'd234} : s = 415;
	{8'd212,8'd235} : s = 507;
	{8'd212,8'd236} : s = 7;
	{8'd212,8'd237} : s = 39;
	{8'd212,8'd238} : s = 30;
	{8'd212,8'd239} : s = 110;
	{8'd212,8'd240} : s = 29;
	{8'd212,8'd241} : s = 109;
	{8'd212,8'd242} : s = 107;
	{8'd212,8'd243} : s = 235;
	{8'd212,8'd244} : s = 27;
	{8'd212,8'd245} : s = 103;
	{8'd212,8'd246} : s = 94;
	{8'd212,8'd247} : s = 231;
	{8'd212,8'd248} : s = 93;
	{8'd212,8'd249} : s = 222;
	{8'd212,8'd250} : s = 221;
	{8'd212,8'd251} : s = 382;
	{8'd212,8'd252} : s = 23;
	{8'd212,8'd253} : s = 91;
	{8'd212,8'd254} : s = 87;
	{8'd212,8'd255} : s = 219;
	{8'd213,8'd0} : s = 361;
	{8'd213,8'd1} : s = 358;
	{8'd213,8'd2} : s = 469;
	{8'd213,8'd3} : s = 209;
	{8'd213,8'd4} : s = 357;
	{8'd213,8'd5} : s = 355;
	{8'd213,8'd6} : s = 467;
	{8'd213,8'd7} : s = 348;
	{8'd213,8'd8} : s = 462;
	{8'd213,8'd9} : s = 461;
	{8'd213,8'd10} : s = 505;
	{8'd213,8'd11} : s = 84;
	{8'd213,8'd12} : s = 204;
	{8'd213,8'd13} : s = 202;
	{8'd213,8'd14} : s = 346;
	{8'd213,8'd15} : s = 201;
	{8'd213,8'd16} : s = 345;
	{8'd213,8'd17} : s = 342;
	{8'd213,8'd18} : s = 459;
	{8'd213,8'd19} : s = 198;
	{8'd213,8'd20} : s = 341;
	{8'd213,8'd21} : s = 339;
	{8'd213,8'd22} : s = 455;
	{8'd213,8'd23} : s = 334;
	{8'd213,8'd24} : s = 444;
	{8'd213,8'd25} : s = 442;
	{8'd213,8'd26} : s = 502;
	{8'd213,8'd27} : s = 197;
	{8'd213,8'd28} : s = 333;
	{8'd213,8'd29} : s = 331;
	{8'd213,8'd30} : s = 441;
	{8'd213,8'd31} : s = 327;
	{8'd213,8'd32} : s = 438;
	{8'd213,8'd33} : s = 437;
	{8'd213,8'd34} : s = 501;
	{8'd213,8'd35} : s = 316;
	{8'd213,8'd36} : s = 435;
	{8'd213,8'd37} : s = 430;
	{8'd213,8'd38} : s = 499;
	{8'd213,8'd39} : s = 429;
	{8'd213,8'd40} : s = 494;
	{8'd213,8'd41} : s = 493;
	{8'd213,8'd42} : s = 510;
	{8'd213,8'd43} : s = 1;
	{8'd213,8'd44} : s = 18;
	{8'd213,8'd45} : s = 17;
	{8'd213,8'd46} : s = 82;
	{8'd213,8'd47} : s = 12;
	{8'd213,8'd48} : s = 81;
	{8'd213,8'd49} : s = 76;
	{8'd213,8'd50} : s = 195;
	{8'd213,8'd51} : s = 10;
	{8'd213,8'd52} : s = 74;
	{8'd213,8'd53} : s = 73;
	{8'd213,8'd54} : s = 184;
	{8'd213,8'd55} : s = 70;
	{8'd213,8'd56} : s = 180;
	{8'd213,8'd57} : s = 178;
	{8'd213,8'd58} : s = 314;
	{8'd213,8'd59} : s = 9;
	{8'd213,8'd60} : s = 69;
	{8'd213,8'd61} : s = 67;
	{8'd213,8'd62} : s = 177;
	{8'd213,8'd63} : s = 56;
	{8'd213,8'd64} : s = 172;
	{8'd213,8'd65} : s = 170;
	{8'd213,8'd66} : s = 313;
	{8'd213,8'd67} : s = 52;
	{8'd213,8'd68} : s = 169;
	{8'd213,8'd69} : s = 166;
	{8'd213,8'd70} : s = 310;
	{8'd213,8'd71} : s = 165;
	{8'd213,8'd72} : s = 309;
	{8'd213,8'd73} : s = 307;
	{8'd213,8'd74} : s = 427;
	{8'd213,8'd75} : s = 6;
	{8'd213,8'd76} : s = 50;
	{8'd213,8'd77} : s = 49;
	{8'd213,8'd78} : s = 163;
	{8'd213,8'd79} : s = 44;
	{8'd213,8'd80} : s = 156;
	{8'd213,8'd81} : s = 154;
	{8'd213,8'd82} : s = 302;
	{8'd213,8'd83} : s = 42;
	{8'd213,8'd84} : s = 153;
	{8'd213,8'd85} : s = 150;
	{8'd213,8'd86} : s = 301;
	{8'd213,8'd87} : s = 149;
	{8'd213,8'd88} : s = 299;
	{8'd213,8'd89} : s = 295;
	{8'd213,8'd90} : s = 423;
	{8'd213,8'd91} : s = 41;
	{8'd213,8'd92} : s = 147;
	{8'd213,8'd93} : s = 142;
	{8'd213,8'd94} : s = 286;
	{8'd213,8'd95} : s = 141;
	{8'd213,8'd96} : s = 285;
	{8'd213,8'd97} : s = 283;
	{8'd213,8'd98} : s = 414;
	{8'd213,8'd99} : s = 139;
	{8'd213,8'd100} : s = 279;
	{8'd213,8'd101} : s = 271;
	{8'd213,8'd102} : s = 413;
	{8'd213,8'd103} : s = 248;
	{8'd213,8'd104} : s = 411;
	{8'd213,8'd105} : s = 407;
	{8'd213,8'd106} : s = 491;
	{8'd213,8'd107} : s = 5;
	{8'd213,8'd108} : s = 38;
	{8'd213,8'd109} : s = 37;
	{8'd213,8'd110} : s = 135;
	{8'd213,8'd111} : s = 35;
	{8'd213,8'd112} : s = 120;
	{8'd213,8'd113} : s = 116;
	{8'd213,8'd114} : s = 244;
	{8'd213,8'd115} : s = 28;
	{8'd213,8'd116} : s = 114;
	{8'd213,8'd117} : s = 113;
	{8'd213,8'd118} : s = 242;
	{8'd213,8'd119} : s = 108;
	{8'd213,8'd120} : s = 241;
	{8'd213,8'd121} : s = 236;
	{8'd213,8'd122} : s = 399;
	{8'd213,8'd123} : s = 26;
	{8'd213,8'd124} : s = 106;
	{8'd213,8'd125} : s = 105;
	{8'd213,8'd126} : s = 234;
	{8'd213,8'd127} : s = 102;
	{8'd213,8'd128} : s = 233;
	{8'd213,8'd129} : s = 230;
	{8'd213,8'd130} : s = 380;
	{8'd213,8'd131} : s = 101;
	{8'd213,8'd132} : s = 229;
	{8'd213,8'd133} : s = 227;
	{8'd213,8'd134} : s = 378;
	{8'd213,8'd135} : s = 220;
	{8'd213,8'd136} : s = 377;
	{8'd213,8'd137} : s = 374;
	{8'd213,8'd138} : s = 487;
	{8'd213,8'd139} : s = 25;
	{8'd213,8'd140} : s = 99;
	{8'd213,8'd141} : s = 92;
	{8'd213,8'd142} : s = 218;
	{8'd213,8'd143} : s = 90;
	{8'd213,8'd144} : s = 217;
	{8'd213,8'd145} : s = 214;
	{8'd213,8'd146} : s = 373;
	{8'd213,8'd147} : s = 89;
	{8'd213,8'd148} : s = 213;
	{8'd213,8'd149} : s = 211;
	{8'd213,8'd150} : s = 371;
	{8'd213,8'd151} : s = 206;
	{8'd213,8'd152} : s = 366;
	{8'd213,8'd153} : s = 365;
	{8'd213,8'd154} : s = 478;
	{8'd213,8'd155} : s = 86;
	{8'd213,8'd156} : s = 205;
	{8'd213,8'd157} : s = 203;
	{8'd213,8'd158} : s = 363;
	{8'd213,8'd159} : s = 199;
	{8'd213,8'd160} : s = 359;
	{8'd213,8'd161} : s = 350;
	{8'd213,8'd162} : s = 477;
	{8'd213,8'd163} : s = 188;
	{8'd213,8'd164} : s = 349;
	{8'd213,8'd165} : s = 347;
	{8'd213,8'd166} : s = 475;
	{8'd213,8'd167} : s = 343;
	{8'd213,8'd168} : s = 471;
	{8'd213,8'd169} : s = 463;
	{8'd213,8'd170} : s = 509;
	{8'd213,8'd171} : s = 3;
	{8'd213,8'd172} : s = 22;
	{8'd213,8'd173} : s = 21;
	{8'd213,8'd174} : s = 85;
	{8'd213,8'd175} : s = 19;
	{8'd213,8'd176} : s = 83;
	{8'd213,8'd177} : s = 78;
	{8'd213,8'd178} : s = 186;
	{8'd213,8'd179} : s = 14;
	{8'd213,8'd180} : s = 77;
	{8'd213,8'd181} : s = 75;
	{8'd213,8'd182} : s = 185;
	{8'd213,8'd183} : s = 71;
	{8'd213,8'd184} : s = 182;
	{8'd213,8'd185} : s = 181;
	{8'd213,8'd186} : s = 335;
	{8'd213,8'd187} : s = 13;
	{8'd213,8'd188} : s = 60;
	{8'd213,8'd189} : s = 58;
	{8'd213,8'd190} : s = 179;
	{8'd213,8'd191} : s = 57;
	{8'd213,8'd192} : s = 174;
	{8'd213,8'd193} : s = 173;
	{8'd213,8'd194} : s = 318;
	{8'd213,8'd195} : s = 54;
	{8'd213,8'd196} : s = 171;
	{8'd213,8'd197} : s = 167;
	{8'd213,8'd198} : s = 317;
	{8'd213,8'd199} : s = 158;
	{8'd213,8'd200} : s = 315;
	{8'd213,8'd201} : s = 311;
	{8'd213,8'd202} : s = 446;
	{8'd213,8'd203} : s = 11;
	{8'd213,8'd204} : s = 53;
	{8'd213,8'd205} : s = 51;
	{8'd213,8'd206} : s = 157;
	{8'd213,8'd207} : s = 46;
	{8'd213,8'd208} : s = 155;
	{8'd213,8'd209} : s = 151;
	{8'd213,8'd210} : s = 303;
	{8'd213,8'd211} : s = 45;
	{8'd213,8'd212} : s = 143;
	{8'd213,8'd213} : s = 124;
	{8'd213,8'd214} : s = 287;
	{8'd213,8'd215} : s = 122;
	{8'd213,8'd216} : s = 252;
	{8'd213,8'd217} : s = 250;
	{8'd213,8'd218} : s = 445;
	{8'd213,8'd219} : s = 43;
	{8'd213,8'd220} : s = 121;
	{8'd213,8'd221} : s = 118;
	{8'd213,8'd222} : s = 249;
	{8'd213,8'd223} : s = 117;
	{8'd213,8'd224} : s = 246;
	{8'd213,8'd225} : s = 245;
	{8'd213,8'd226} : s = 443;
	{8'd213,8'd227} : s = 115;
	{8'd213,8'd228} : s = 243;
	{8'd213,8'd229} : s = 238;
	{8'd213,8'd230} : s = 439;
	{8'd213,8'd231} : s = 237;
	{8'd213,8'd232} : s = 431;
	{8'd213,8'd233} : s = 415;
	{8'd213,8'd234} : s = 507;
	{8'd213,8'd235} : s = 7;
	{8'd213,8'd236} : s = 39;
	{8'd213,8'd237} : s = 30;
	{8'd213,8'd238} : s = 110;
	{8'd213,8'd239} : s = 29;
	{8'd213,8'd240} : s = 109;
	{8'd213,8'd241} : s = 107;
	{8'd213,8'd242} : s = 235;
	{8'd213,8'd243} : s = 27;
	{8'd213,8'd244} : s = 103;
	{8'd213,8'd245} : s = 94;
	{8'd213,8'd246} : s = 231;
	{8'd213,8'd247} : s = 93;
	{8'd213,8'd248} : s = 222;
	{8'd213,8'd249} : s = 221;
	{8'd213,8'd250} : s = 382;
	{8'd213,8'd251} : s = 23;
	{8'd213,8'd252} : s = 91;
	{8'd213,8'd253} : s = 87;
	{8'd213,8'd254} : s = 219;
	{8'd213,8'd255} : s = 79;
	{8'd214,8'd0} : s = 358;
	{8'd214,8'd1} : s = 469;
	{8'd214,8'd2} : s = 209;
	{8'd214,8'd3} : s = 357;
	{8'd214,8'd4} : s = 355;
	{8'd214,8'd5} : s = 467;
	{8'd214,8'd6} : s = 348;
	{8'd214,8'd7} : s = 462;
	{8'd214,8'd8} : s = 461;
	{8'd214,8'd9} : s = 505;
	{8'd214,8'd10} : s = 84;
	{8'd214,8'd11} : s = 204;
	{8'd214,8'd12} : s = 202;
	{8'd214,8'd13} : s = 346;
	{8'd214,8'd14} : s = 201;
	{8'd214,8'd15} : s = 345;
	{8'd214,8'd16} : s = 342;
	{8'd214,8'd17} : s = 459;
	{8'd214,8'd18} : s = 198;
	{8'd214,8'd19} : s = 341;
	{8'd214,8'd20} : s = 339;
	{8'd214,8'd21} : s = 455;
	{8'd214,8'd22} : s = 334;
	{8'd214,8'd23} : s = 444;
	{8'd214,8'd24} : s = 442;
	{8'd214,8'd25} : s = 502;
	{8'd214,8'd26} : s = 197;
	{8'd214,8'd27} : s = 333;
	{8'd214,8'd28} : s = 331;
	{8'd214,8'd29} : s = 441;
	{8'd214,8'd30} : s = 327;
	{8'd214,8'd31} : s = 438;
	{8'd214,8'd32} : s = 437;
	{8'd214,8'd33} : s = 501;
	{8'd214,8'd34} : s = 316;
	{8'd214,8'd35} : s = 435;
	{8'd214,8'd36} : s = 430;
	{8'd214,8'd37} : s = 499;
	{8'd214,8'd38} : s = 429;
	{8'd214,8'd39} : s = 494;
	{8'd214,8'd40} : s = 493;
	{8'd214,8'd41} : s = 510;
	{8'd214,8'd42} : s = 1;
	{8'd214,8'd43} : s = 18;
	{8'd214,8'd44} : s = 17;
	{8'd214,8'd45} : s = 82;
	{8'd214,8'd46} : s = 12;
	{8'd214,8'd47} : s = 81;
	{8'd214,8'd48} : s = 76;
	{8'd214,8'd49} : s = 195;
	{8'd214,8'd50} : s = 10;
	{8'd214,8'd51} : s = 74;
	{8'd214,8'd52} : s = 73;
	{8'd214,8'd53} : s = 184;
	{8'd214,8'd54} : s = 70;
	{8'd214,8'd55} : s = 180;
	{8'd214,8'd56} : s = 178;
	{8'd214,8'd57} : s = 314;
	{8'd214,8'd58} : s = 9;
	{8'd214,8'd59} : s = 69;
	{8'd214,8'd60} : s = 67;
	{8'd214,8'd61} : s = 177;
	{8'd214,8'd62} : s = 56;
	{8'd214,8'd63} : s = 172;
	{8'd214,8'd64} : s = 170;
	{8'd214,8'd65} : s = 313;
	{8'd214,8'd66} : s = 52;
	{8'd214,8'd67} : s = 169;
	{8'd214,8'd68} : s = 166;
	{8'd214,8'd69} : s = 310;
	{8'd214,8'd70} : s = 165;
	{8'd214,8'd71} : s = 309;
	{8'd214,8'd72} : s = 307;
	{8'd214,8'd73} : s = 427;
	{8'd214,8'd74} : s = 6;
	{8'd214,8'd75} : s = 50;
	{8'd214,8'd76} : s = 49;
	{8'd214,8'd77} : s = 163;
	{8'd214,8'd78} : s = 44;
	{8'd214,8'd79} : s = 156;
	{8'd214,8'd80} : s = 154;
	{8'd214,8'd81} : s = 302;
	{8'd214,8'd82} : s = 42;
	{8'd214,8'd83} : s = 153;
	{8'd214,8'd84} : s = 150;
	{8'd214,8'd85} : s = 301;
	{8'd214,8'd86} : s = 149;
	{8'd214,8'd87} : s = 299;
	{8'd214,8'd88} : s = 295;
	{8'd214,8'd89} : s = 423;
	{8'd214,8'd90} : s = 41;
	{8'd214,8'd91} : s = 147;
	{8'd214,8'd92} : s = 142;
	{8'd214,8'd93} : s = 286;
	{8'd214,8'd94} : s = 141;
	{8'd214,8'd95} : s = 285;
	{8'd214,8'd96} : s = 283;
	{8'd214,8'd97} : s = 414;
	{8'd214,8'd98} : s = 139;
	{8'd214,8'd99} : s = 279;
	{8'd214,8'd100} : s = 271;
	{8'd214,8'd101} : s = 413;
	{8'd214,8'd102} : s = 248;
	{8'd214,8'd103} : s = 411;
	{8'd214,8'd104} : s = 407;
	{8'd214,8'd105} : s = 491;
	{8'd214,8'd106} : s = 5;
	{8'd214,8'd107} : s = 38;
	{8'd214,8'd108} : s = 37;
	{8'd214,8'd109} : s = 135;
	{8'd214,8'd110} : s = 35;
	{8'd214,8'd111} : s = 120;
	{8'd214,8'd112} : s = 116;
	{8'd214,8'd113} : s = 244;
	{8'd214,8'd114} : s = 28;
	{8'd214,8'd115} : s = 114;
	{8'd214,8'd116} : s = 113;
	{8'd214,8'd117} : s = 242;
	{8'd214,8'd118} : s = 108;
	{8'd214,8'd119} : s = 241;
	{8'd214,8'd120} : s = 236;
	{8'd214,8'd121} : s = 399;
	{8'd214,8'd122} : s = 26;
	{8'd214,8'd123} : s = 106;
	{8'd214,8'd124} : s = 105;
	{8'd214,8'd125} : s = 234;
	{8'd214,8'd126} : s = 102;
	{8'd214,8'd127} : s = 233;
	{8'd214,8'd128} : s = 230;
	{8'd214,8'd129} : s = 380;
	{8'd214,8'd130} : s = 101;
	{8'd214,8'd131} : s = 229;
	{8'd214,8'd132} : s = 227;
	{8'd214,8'd133} : s = 378;
	{8'd214,8'd134} : s = 220;
	{8'd214,8'd135} : s = 377;
	{8'd214,8'd136} : s = 374;
	{8'd214,8'd137} : s = 487;
	{8'd214,8'd138} : s = 25;
	{8'd214,8'd139} : s = 99;
	{8'd214,8'd140} : s = 92;
	{8'd214,8'd141} : s = 218;
	{8'd214,8'd142} : s = 90;
	{8'd214,8'd143} : s = 217;
	{8'd214,8'd144} : s = 214;
	{8'd214,8'd145} : s = 373;
	{8'd214,8'd146} : s = 89;
	{8'd214,8'd147} : s = 213;
	{8'd214,8'd148} : s = 211;
	{8'd214,8'd149} : s = 371;
	{8'd214,8'd150} : s = 206;
	{8'd214,8'd151} : s = 366;
	{8'd214,8'd152} : s = 365;
	{8'd214,8'd153} : s = 478;
	{8'd214,8'd154} : s = 86;
	{8'd214,8'd155} : s = 205;
	{8'd214,8'd156} : s = 203;
	{8'd214,8'd157} : s = 363;
	{8'd214,8'd158} : s = 199;
	{8'd214,8'd159} : s = 359;
	{8'd214,8'd160} : s = 350;
	{8'd214,8'd161} : s = 477;
	{8'd214,8'd162} : s = 188;
	{8'd214,8'd163} : s = 349;
	{8'd214,8'd164} : s = 347;
	{8'd214,8'd165} : s = 475;
	{8'd214,8'd166} : s = 343;
	{8'd214,8'd167} : s = 471;
	{8'd214,8'd168} : s = 463;
	{8'd214,8'd169} : s = 509;
	{8'd214,8'd170} : s = 3;
	{8'd214,8'd171} : s = 22;
	{8'd214,8'd172} : s = 21;
	{8'd214,8'd173} : s = 85;
	{8'd214,8'd174} : s = 19;
	{8'd214,8'd175} : s = 83;
	{8'd214,8'd176} : s = 78;
	{8'd214,8'd177} : s = 186;
	{8'd214,8'd178} : s = 14;
	{8'd214,8'd179} : s = 77;
	{8'd214,8'd180} : s = 75;
	{8'd214,8'd181} : s = 185;
	{8'd214,8'd182} : s = 71;
	{8'd214,8'd183} : s = 182;
	{8'd214,8'd184} : s = 181;
	{8'd214,8'd185} : s = 335;
	{8'd214,8'd186} : s = 13;
	{8'd214,8'd187} : s = 60;
	{8'd214,8'd188} : s = 58;
	{8'd214,8'd189} : s = 179;
	{8'd214,8'd190} : s = 57;
	{8'd214,8'd191} : s = 174;
	{8'd214,8'd192} : s = 173;
	{8'd214,8'd193} : s = 318;
	{8'd214,8'd194} : s = 54;
	{8'd214,8'd195} : s = 171;
	{8'd214,8'd196} : s = 167;
	{8'd214,8'd197} : s = 317;
	{8'd214,8'd198} : s = 158;
	{8'd214,8'd199} : s = 315;
	{8'd214,8'd200} : s = 311;
	{8'd214,8'd201} : s = 446;
	{8'd214,8'd202} : s = 11;
	{8'd214,8'd203} : s = 53;
	{8'd214,8'd204} : s = 51;
	{8'd214,8'd205} : s = 157;
	{8'd214,8'd206} : s = 46;
	{8'd214,8'd207} : s = 155;
	{8'd214,8'd208} : s = 151;
	{8'd214,8'd209} : s = 303;
	{8'd214,8'd210} : s = 45;
	{8'd214,8'd211} : s = 143;
	{8'd214,8'd212} : s = 124;
	{8'd214,8'd213} : s = 287;
	{8'd214,8'd214} : s = 122;
	{8'd214,8'd215} : s = 252;
	{8'd214,8'd216} : s = 250;
	{8'd214,8'd217} : s = 445;
	{8'd214,8'd218} : s = 43;
	{8'd214,8'd219} : s = 121;
	{8'd214,8'd220} : s = 118;
	{8'd214,8'd221} : s = 249;
	{8'd214,8'd222} : s = 117;
	{8'd214,8'd223} : s = 246;
	{8'd214,8'd224} : s = 245;
	{8'd214,8'd225} : s = 443;
	{8'd214,8'd226} : s = 115;
	{8'd214,8'd227} : s = 243;
	{8'd214,8'd228} : s = 238;
	{8'd214,8'd229} : s = 439;
	{8'd214,8'd230} : s = 237;
	{8'd214,8'd231} : s = 431;
	{8'd214,8'd232} : s = 415;
	{8'd214,8'd233} : s = 507;
	{8'd214,8'd234} : s = 7;
	{8'd214,8'd235} : s = 39;
	{8'd214,8'd236} : s = 30;
	{8'd214,8'd237} : s = 110;
	{8'd214,8'd238} : s = 29;
	{8'd214,8'd239} : s = 109;
	{8'd214,8'd240} : s = 107;
	{8'd214,8'd241} : s = 235;
	{8'd214,8'd242} : s = 27;
	{8'd214,8'd243} : s = 103;
	{8'd214,8'd244} : s = 94;
	{8'd214,8'd245} : s = 231;
	{8'd214,8'd246} : s = 93;
	{8'd214,8'd247} : s = 222;
	{8'd214,8'd248} : s = 221;
	{8'd214,8'd249} : s = 382;
	{8'd214,8'd250} : s = 23;
	{8'd214,8'd251} : s = 91;
	{8'd214,8'd252} : s = 87;
	{8'd214,8'd253} : s = 219;
	{8'd214,8'd254} : s = 79;
	{8'd214,8'd255} : s = 215;
	{8'd215,8'd0} : s = 469;
	{8'd215,8'd1} : s = 209;
	{8'd215,8'd2} : s = 357;
	{8'd215,8'd3} : s = 355;
	{8'd215,8'd4} : s = 467;
	{8'd215,8'd5} : s = 348;
	{8'd215,8'd6} : s = 462;
	{8'd215,8'd7} : s = 461;
	{8'd215,8'd8} : s = 505;
	{8'd215,8'd9} : s = 84;
	{8'd215,8'd10} : s = 204;
	{8'd215,8'd11} : s = 202;
	{8'd215,8'd12} : s = 346;
	{8'd215,8'd13} : s = 201;
	{8'd215,8'd14} : s = 345;
	{8'd215,8'd15} : s = 342;
	{8'd215,8'd16} : s = 459;
	{8'd215,8'd17} : s = 198;
	{8'd215,8'd18} : s = 341;
	{8'd215,8'd19} : s = 339;
	{8'd215,8'd20} : s = 455;
	{8'd215,8'd21} : s = 334;
	{8'd215,8'd22} : s = 444;
	{8'd215,8'd23} : s = 442;
	{8'd215,8'd24} : s = 502;
	{8'd215,8'd25} : s = 197;
	{8'd215,8'd26} : s = 333;
	{8'd215,8'd27} : s = 331;
	{8'd215,8'd28} : s = 441;
	{8'd215,8'd29} : s = 327;
	{8'd215,8'd30} : s = 438;
	{8'd215,8'd31} : s = 437;
	{8'd215,8'd32} : s = 501;
	{8'd215,8'd33} : s = 316;
	{8'd215,8'd34} : s = 435;
	{8'd215,8'd35} : s = 430;
	{8'd215,8'd36} : s = 499;
	{8'd215,8'd37} : s = 429;
	{8'd215,8'd38} : s = 494;
	{8'd215,8'd39} : s = 493;
	{8'd215,8'd40} : s = 510;
	{8'd215,8'd41} : s = 1;
	{8'd215,8'd42} : s = 18;
	{8'd215,8'd43} : s = 17;
	{8'd215,8'd44} : s = 82;
	{8'd215,8'd45} : s = 12;
	{8'd215,8'd46} : s = 81;
	{8'd215,8'd47} : s = 76;
	{8'd215,8'd48} : s = 195;
	{8'd215,8'd49} : s = 10;
	{8'd215,8'd50} : s = 74;
	{8'd215,8'd51} : s = 73;
	{8'd215,8'd52} : s = 184;
	{8'd215,8'd53} : s = 70;
	{8'd215,8'd54} : s = 180;
	{8'd215,8'd55} : s = 178;
	{8'd215,8'd56} : s = 314;
	{8'd215,8'd57} : s = 9;
	{8'd215,8'd58} : s = 69;
	{8'd215,8'd59} : s = 67;
	{8'd215,8'd60} : s = 177;
	{8'd215,8'd61} : s = 56;
	{8'd215,8'd62} : s = 172;
	{8'd215,8'd63} : s = 170;
	{8'd215,8'd64} : s = 313;
	{8'd215,8'd65} : s = 52;
	{8'd215,8'd66} : s = 169;
	{8'd215,8'd67} : s = 166;
	{8'd215,8'd68} : s = 310;
	{8'd215,8'd69} : s = 165;
	{8'd215,8'd70} : s = 309;
	{8'd215,8'd71} : s = 307;
	{8'd215,8'd72} : s = 427;
	{8'd215,8'd73} : s = 6;
	{8'd215,8'd74} : s = 50;
	{8'd215,8'd75} : s = 49;
	{8'd215,8'd76} : s = 163;
	{8'd215,8'd77} : s = 44;
	{8'd215,8'd78} : s = 156;
	{8'd215,8'd79} : s = 154;
	{8'd215,8'd80} : s = 302;
	{8'd215,8'd81} : s = 42;
	{8'd215,8'd82} : s = 153;
	{8'd215,8'd83} : s = 150;
	{8'd215,8'd84} : s = 301;
	{8'd215,8'd85} : s = 149;
	{8'd215,8'd86} : s = 299;
	{8'd215,8'd87} : s = 295;
	{8'd215,8'd88} : s = 423;
	{8'd215,8'd89} : s = 41;
	{8'd215,8'd90} : s = 147;
	{8'd215,8'd91} : s = 142;
	{8'd215,8'd92} : s = 286;
	{8'd215,8'd93} : s = 141;
	{8'd215,8'd94} : s = 285;
	{8'd215,8'd95} : s = 283;
	{8'd215,8'd96} : s = 414;
	{8'd215,8'd97} : s = 139;
	{8'd215,8'd98} : s = 279;
	{8'd215,8'd99} : s = 271;
	{8'd215,8'd100} : s = 413;
	{8'd215,8'd101} : s = 248;
	{8'd215,8'd102} : s = 411;
	{8'd215,8'd103} : s = 407;
	{8'd215,8'd104} : s = 491;
	{8'd215,8'd105} : s = 5;
	{8'd215,8'd106} : s = 38;
	{8'd215,8'd107} : s = 37;
	{8'd215,8'd108} : s = 135;
	{8'd215,8'd109} : s = 35;
	{8'd215,8'd110} : s = 120;
	{8'd215,8'd111} : s = 116;
	{8'd215,8'd112} : s = 244;
	{8'd215,8'd113} : s = 28;
	{8'd215,8'd114} : s = 114;
	{8'd215,8'd115} : s = 113;
	{8'd215,8'd116} : s = 242;
	{8'd215,8'd117} : s = 108;
	{8'd215,8'd118} : s = 241;
	{8'd215,8'd119} : s = 236;
	{8'd215,8'd120} : s = 399;
	{8'd215,8'd121} : s = 26;
	{8'd215,8'd122} : s = 106;
	{8'd215,8'd123} : s = 105;
	{8'd215,8'd124} : s = 234;
	{8'd215,8'd125} : s = 102;
	{8'd215,8'd126} : s = 233;
	{8'd215,8'd127} : s = 230;
	{8'd215,8'd128} : s = 380;
	{8'd215,8'd129} : s = 101;
	{8'd215,8'd130} : s = 229;
	{8'd215,8'd131} : s = 227;
	{8'd215,8'd132} : s = 378;
	{8'd215,8'd133} : s = 220;
	{8'd215,8'd134} : s = 377;
	{8'd215,8'd135} : s = 374;
	{8'd215,8'd136} : s = 487;
	{8'd215,8'd137} : s = 25;
	{8'd215,8'd138} : s = 99;
	{8'd215,8'd139} : s = 92;
	{8'd215,8'd140} : s = 218;
	{8'd215,8'd141} : s = 90;
	{8'd215,8'd142} : s = 217;
	{8'd215,8'd143} : s = 214;
	{8'd215,8'd144} : s = 373;
	{8'd215,8'd145} : s = 89;
	{8'd215,8'd146} : s = 213;
	{8'd215,8'd147} : s = 211;
	{8'd215,8'd148} : s = 371;
	{8'd215,8'd149} : s = 206;
	{8'd215,8'd150} : s = 366;
	{8'd215,8'd151} : s = 365;
	{8'd215,8'd152} : s = 478;
	{8'd215,8'd153} : s = 86;
	{8'd215,8'd154} : s = 205;
	{8'd215,8'd155} : s = 203;
	{8'd215,8'd156} : s = 363;
	{8'd215,8'd157} : s = 199;
	{8'd215,8'd158} : s = 359;
	{8'd215,8'd159} : s = 350;
	{8'd215,8'd160} : s = 477;
	{8'd215,8'd161} : s = 188;
	{8'd215,8'd162} : s = 349;
	{8'd215,8'd163} : s = 347;
	{8'd215,8'd164} : s = 475;
	{8'd215,8'd165} : s = 343;
	{8'd215,8'd166} : s = 471;
	{8'd215,8'd167} : s = 463;
	{8'd215,8'd168} : s = 509;
	{8'd215,8'd169} : s = 3;
	{8'd215,8'd170} : s = 22;
	{8'd215,8'd171} : s = 21;
	{8'd215,8'd172} : s = 85;
	{8'd215,8'd173} : s = 19;
	{8'd215,8'd174} : s = 83;
	{8'd215,8'd175} : s = 78;
	{8'd215,8'd176} : s = 186;
	{8'd215,8'd177} : s = 14;
	{8'd215,8'd178} : s = 77;
	{8'd215,8'd179} : s = 75;
	{8'd215,8'd180} : s = 185;
	{8'd215,8'd181} : s = 71;
	{8'd215,8'd182} : s = 182;
	{8'd215,8'd183} : s = 181;
	{8'd215,8'd184} : s = 335;
	{8'd215,8'd185} : s = 13;
	{8'd215,8'd186} : s = 60;
	{8'd215,8'd187} : s = 58;
	{8'd215,8'd188} : s = 179;
	{8'd215,8'd189} : s = 57;
	{8'd215,8'd190} : s = 174;
	{8'd215,8'd191} : s = 173;
	{8'd215,8'd192} : s = 318;
	{8'd215,8'd193} : s = 54;
	{8'd215,8'd194} : s = 171;
	{8'd215,8'd195} : s = 167;
	{8'd215,8'd196} : s = 317;
	{8'd215,8'd197} : s = 158;
	{8'd215,8'd198} : s = 315;
	{8'd215,8'd199} : s = 311;
	{8'd215,8'd200} : s = 446;
	{8'd215,8'd201} : s = 11;
	{8'd215,8'd202} : s = 53;
	{8'd215,8'd203} : s = 51;
	{8'd215,8'd204} : s = 157;
	{8'd215,8'd205} : s = 46;
	{8'd215,8'd206} : s = 155;
	{8'd215,8'd207} : s = 151;
	{8'd215,8'd208} : s = 303;
	{8'd215,8'd209} : s = 45;
	{8'd215,8'd210} : s = 143;
	{8'd215,8'd211} : s = 124;
	{8'd215,8'd212} : s = 287;
	{8'd215,8'd213} : s = 122;
	{8'd215,8'd214} : s = 252;
	{8'd215,8'd215} : s = 250;
	{8'd215,8'd216} : s = 445;
	{8'd215,8'd217} : s = 43;
	{8'd215,8'd218} : s = 121;
	{8'd215,8'd219} : s = 118;
	{8'd215,8'd220} : s = 249;
	{8'd215,8'd221} : s = 117;
	{8'd215,8'd222} : s = 246;
	{8'd215,8'd223} : s = 245;
	{8'd215,8'd224} : s = 443;
	{8'd215,8'd225} : s = 115;
	{8'd215,8'd226} : s = 243;
	{8'd215,8'd227} : s = 238;
	{8'd215,8'd228} : s = 439;
	{8'd215,8'd229} : s = 237;
	{8'd215,8'd230} : s = 431;
	{8'd215,8'd231} : s = 415;
	{8'd215,8'd232} : s = 507;
	{8'd215,8'd233} : s = 7;
	{8'd215,8'd234} : s = 39;
	{8'd215,8'd235} : s = 30;
	{8'd215,8'd236} : s = 110;
	{8'd215,8'd237} : s = 29;
	{8'd215,8'd238} : s = 109;
	{8'd215,8'd239} : s = 107;
	{8'd215,8'd240} : s = 235;
	{8'd215,8'd241} : s = 27;
	{8'd215,8'd242} : s = 103;
	{8'd215,8'd243} : s = 94;
	{8'd215,8'd244} : s = 231;
	{8'd215,8'd245} : s = 93;
	{8'd215,8'd246} : s = 222;
	{8'd215,8'd247} : s = 221;
	{8'd215,8'd248} : s = 382;
	{8'd215,8'd249} : s = 23;
	{8'd215,8'd250} : s = 91;
	{8'd215,8'd251} : s = 87;
	{8'd215,8'd252} : s = 219;
	{8'd215,8'd253} : s = 79;
	{8'd215,8'd254} : s = 215;
	{8'd215,8'd255} : s = 207;
	{8'd216,8'd0} : s = 209;
	{8'd216,8'd1} : s = 357;
	{8'd216,8'd2} : s = 355;
	{8'd216,8'd3} : s = 467;
	{8'd216,8'd4} : s = 348;
	{8'd216,8'd5} : s = 462;
	{8'd216,8'd6} : s = 461;
	{8'd216,8'd7} : s = 505;
	{8'd216,8'd8} : s = 84;
	{8'd216,8'd9} : s = 204;
	{8'd216,8'd10} : s = 202;
	{8'd216,8'd11} : s = 346;
	{8'd216,8'd12} : s = 201;
	{8'd216,8'd13} : s = 345;
	{8'd216,8'd14} : s = 342;
	{8'd216,8'd15} : s = 459;
	{8'd216,8'd16} : s = 198;
	{8'd216,8'd17} : s = 341;
	{8'd216,8'd18} : s = 339;
	{8'd216,8'd19} : s = 455;
	{8'd216,8'd20} : s = 334;
	{8'd216,8'd21} : s = 444;
	{8'd216,8'd22} : s = 442;
	{8'd216,8'd23} : s = 502;
	{8'd216,8'd24} : s = 197;
	{8'd216,8'd25} : s = 333;
	{8'd216,8'd26} : s = 331;
	{8'd216,8'd27} : s = 441;
	{8'd216,8'd28} : s = 327;
	{8'd216,8'd29} : s = 438;
	{8'd216,8'd30} : s = 437;
	{8'd216,8'd31} : s = 501;
	{8'd216,8'd32} : s = 316;
	{8'd216,8'd33} : s = 435;
	{8'd216,8'd34} : s = 430;
	{8'd216,8'd35} : s = 499;
	{8'd216,8'd36} : s = 429;
	{8'd216,8'd37} : s = 494;
	{8'd216,8'd38} : s = 493;
	{8'd216,8'd39} : s = 510;
	{8'd216,8'd40} : s = 1;
	{8'd216,8'd41} : s = 18;
	{8'd216,8'd42} : s = 17;
	{8'd216,8'd43} : s = 82;
	{8'd216,8'd44} : s = 12;
	{8'd216,8'd45} : s = 81;
	{8'd216,8'd46} : s = 76;
	{8'd216,8'd47} : s = 195;
	{8'd216,8'd48} : s = 10;
	{8'd216,8'd49} : s = 74;
	{8'd216,8'd50} : s = 73;
	{8'd216,8'd51} : s = 184;
	{8'd216,8'd52} : s = 70;
	{8'd216,8'd53} : s = 180;
	{8'd216,8'd54} : s = 178;
	{8'd216,8'd55} : s = 314;
	{8'd216,8'd56} : s = 9;
	{8'd216,8'd57} : s = 69;
	{8'd216,8'd58} : s = 67;
	{8'd216,8'd59} : s = 177;
	{8'd216,8'd60} : s = 56;
	{8'd216,8'd61} : s = 172;
	{8'd216,8'd62} : s = 170;
	{8'd216,8'd63} : s = 313;
	{8'd216,8'd64} : s = 52;
	{8'd216,8'd65} : s = 169;
	{8'd216,8'd66} : s = 166;
	{8'd216,8'd67} : s = 310;
	{8'd216,8'd68} : s = 165;
	{8'd216,8'd69} : s = 309;
	{8'd216,8'd70} : s = 307;
	{8'd216,8'd71} : s = 427;
	{8'd216,8'd72} : s = 6;
	{8'd216,8'd73} : s = 50;
	{8'd216,8'd74} : s = 49;
	{8'd216,8'd75} : s = 163;
	{8'd216,8'd76} : s = 44;
	{8'd216,8'd77} : s = 156;
	{8'd216,8'd78} : s = 154;
	{8'd216,8'd79} : s = 302;
	{8'd216,8'd80} : s = 42;
	{8'd216,8'd81} : s = 153;
	{8'd216,8'd82} : s = 150;
	{8'd216,8'd83} : s = 301;
	{8'd216,8'd84} : s = 149;
	{8'd216,8'd85} : s = 299;
	{8'd216,8'd86} : s = 295;
	{8'd216,8'd87} : s = 423;
	{8'd216,8'd88} : s = 41;
	{8'd216,8'd89} : s = 147;
	{8'd216,8'd90} : s = 142;
	{8'd216,8'd91} : s = 286;
	{8'd216,8'd92} : s = 141;
	{8'd216,8'd93} : s = 285;
	{8'd216,8'd94} : s = 283;
	{8'd216,8'd95} : s = 414;
	{8'd216,8'd96} : s = 139;
	{8'd216,8'd97} : s = 279;
	{8'd216,8'd98} : s = 271;
	{8'd216,8'd99} : s = 413;
	{8'd216,8'd100} : s = 248;
	{8'd216,8'd101} : s = 411;
	{8'd216,8'd102} : s = 407;
	{8'd216,8'd103} : s = 491;
	{8'd216,8'd104} : s = 5;
	{8'd216,8'd105} : s = 38;
	{8'd216,8'd106} : s = 37;
	{8'd216,8'd107} : s = 135;
	{8'd216,8'd108} : s = 35;
	{8'd216,8'd109} : s = 120;
	{8'd216,8'd110} : s = 116;
	{8'd216,8'd111} : s = 244;
	{8'd216,8'd112} : s = 28;
	{8'd216,8'd113} : s = 114;
	{8'd216,8'd114} : s = 113;
	{8'd216,8'd115} : s = 242;
	{8'd216,8'd116} : s = 108;
	{8'd216,8'd117} : s = 241;
	{8'd216,8'd118} : s = 236;
	{8'd216,8'd119} : s = 399;
	{8'd216,8'd120} : s = 26;
	{8'd216,8'd121} : s = 106;
	{8'd216,8'd122} : s = 105;
	{8'd216,8'd123} : s = 234;
	{8'd216,8'd124} : s = 102;
	{8'd216,8'd125} : s = 233;
	{8'd216,8'd126} : s = 230;
	{8'd216,8'd127} : s = 380;
	{8'd216,8'd128} : s = 101;
	{8'd216,8'd129} : s = 229;
	{8'd216,8'd130} : s = 227;
	{8'd216,8'd131} : s = 378;
	{8'd216,8'd132} : s = 220;
	{8'd216,8'd133} : s = 377;
	{8'd216,8'd134} : s = 374;
	{8'd216,8'd135} : s = 487;
	{8'd216,8'd136} : s = 25;
	{8'd216,8'd137} : s = 99;
	{8'd216,8'd138} : s = 92;
	{8'd216,8'd139} : s = 218;
	{8'd216,8'd140} : s = 90;
	{8'd216,8'd141} : s = 217;
	{8'd216,8'd142} : s = 214;
	{8'd216,8'd143} : s = 373;
	{8'd216,8'd144} : s = 89;
	{8'd216,8'd145} : s = 213;
	{8'd216,8'd146} : s = 211;
	{8'd216,8'd147} : s = 371;
	{8'd216,8'd148} : s = 206;
	{8'd216,8'd149} : s = 366;
	{8'd216,8'd150} : s = 365;
	{8'd216,8'd151} : s = 478;
	{8'd216,8'd152} : s = 86;
	{8'd216,8'd153} : s = 205;
	{8'd216,8'd154} : s = 203;
	{8'd216,8'd155} : s = 363;
	{8'd216,8'd156} : s = 199;
	{8'd216,8'd157} : s = 359;
	{8'd216,8'd158} : s = 350;
	{8'd216,8'd159} : s = 477;
	{8'd216,8'd160} : s = 188;
	{8'd216,8'd161} : s = 349;
	{8'd216,8'd162} : s = 347;
	{8'd216,8'd163} : s = 475;
	{8'd216,8'd164} : s = 343;
	{8'd216,8'd165} : s = 471;
	{8'd216,8'd166} : s = 463;
	{8'd216,8'd167} : s = 509;
	{8'd216,8'd168} : s = 3;
	{8'd216,8'd169} : s = 22;
	{8'd216,8'd170} : s = 21;
	{8'd216,8'd171} : s = 85;
	{8'd216,8'd172} : s = 19;
	{8'd216,8'd173} : s = 83;
	{8'd216,8'd174} : s = 78;
	{8'd216,8'd175} : s = 186;
	{8'd216,8'd176} : s = 14;
	{8'd216,8'd177} : s = 77;
	{8'd216,8'd178} : s = 75;
	{8'd216,8'd179} : s = 185;
	{8'd216,8'd180} : s = 71;
	{8'd216,8'd181} : s = 182;
	{8'd216,8'd182} : s = 181;
	{8'd216,8'd183} : s = 335;
	{8'd216,8'd184} : s = 13;
	{8'd216,8'd185} : s = 60;
	{8'd216,8'd186} : s = 58;
	{8'd216,8'd187} : s = 179;
	{8'd216,8'd188} : s = 57;
	{8'd216,8'd189} : s = 174;
	{8'd216,8'd190} : s = 173;
	{8'd216,8'd191} : s = 318;
	{8'd216,8'd192} : s = 54;
	{8'd216,8'd193} : s = 171;
	{8'd216,8'd194} : s = 167;
	{8'd216,8'd195} : s = 317;
	{8'd216,8'd196} : s = 158;
	{8'd216,8'd197} : s = 315;
	{8'd216,8'd198} : s = 311;
	{8'd216,8'd199} : s = 446;
	{8'd216,8'd200} : s = 11;
	{8'd216,8'd201} : s = 53;
	{8'd216,8'd202} : s = 51;
	{8'd216,8'd203} : s = 157;
	{8'd216,8'd204} : s = 46;
	{8'd216,8'd205} : s = 155;
	{8'd216,8'd206} : s = 151;
	{8'd216,8'd207} : s = 303;
	{8'd216,8'd208} : s = 45;
	{8'd216,8'd209} : s = 143;
	{8'd216,8'd210} : s = 124;
	{8'd216,8'd211} : s = 287;
	{8'd216,8'd212} : s = 122;
	{8'd216,8'd213} : s = 252;
	{8'd216,8'd214} : s = 250;
	{8'd216,8'd215} : s = 445;
	{8'd216,8'd216} : s = 43;
	{8'd216,8'd217} : s = 121;
	{8'd216,8'd218} : s = 118;
	{8'd216,8'd219} : s = 249;
	{8'd216,8'd220} : s = 117;
	{8'd216,8'd221} : s = 246;
	{8'd216,8'd222} : s = 245;
	{8'd216,8'd223} : s = 443;
	{8'd216,8'd224} : s = 115;
	{8'd216,8'd225} : s = 243;
	{8'd216,8'd226} : s = 238;
	{8'd216,8'd227} : s = 439;
	{8'd216,8'd228} : s = 237;
	{8'd216,8'd229} : s = 431;
	{8'd216,8'd230} : s = 415;
	{8'd216,8'd231} : s = 507;
	{8'd216,8'd232} : s = 7;
	{8'd216,8'd233} : s = 39;
	{8'd216,8'd234} : s = 30;
	{8'd216,8'd235} : s = 110;
	{8'd216,8'd236} : s = 29;
	{8'd216,8'd237} : s = 109;
	{8'd216,8'd238} : s = 107;
	{8'd216,8'd239} : s = 235;
	{8'd216,8'd240} : s = 27;
	{8'd216,8'd241} : s = 103;
	{8'd216,8'd242} : s = 94;
	{8'd216,8'd243} : s = 231;
	{8'd216,8'd244} : s = 93;
	{8'd216,8'd245} : s = 222;
	{8'd216,8'd246} : s = 221;
	{8'd216,8'd247} : s = 382;
	{8'd216,8'd248} : s = 23;
	{8'd216,8'd249} : s = 91;
	{8'd216,8'd250} : s = 87;
	{8'd216,8'd251} : s = 219;
	{8'd216,8'd252} : s = 79;
	{8'd216,8'd253} : s = 215;
	{8'd216,8'd254} : s = 207;
	{8'd216,8'd255} : s = 381;
	{8'd217,8'd0} : s = 357;
	{8'd217,8'd1} : s = 355;
	{8'd217,8'd2} : s = 467;
	{8'd217,8'd3} : s = 348;
	{8'd217,8'd4} : s = 462;
	{8'd217,8'd5} : s = 461;
	{8'd217,8'd6} : s = 505;
	{8'd217,8'd7} : s = 84;
	{8'd217,8'd8} : s = 204;
	{8'd217,8'd9} : s = 202;
	{8'd217,8'd10} : s = 346;
	{8'd217,8'd11} : s = 201;
	{8'd217,8'd12} : s = 345;
	{8'd217,8'd13} : s = 342;
	{8'd217,8'd14} : s = 459;
	{8'd217,8'd15} : s = 198;
	{8'd217,8'd16} : s = 341;
	{8'd217,8'd17} : s = 339;
	{8'd217,8'd18} : s = 455;
	{8'd217,8'd19} : s = 334;
	{8'd217,8'd20} : s = 444;
	{8'd217,8'd21} : s = 442;
	{8'd217,8'd22} : s = 502;
	{8'd217,8'd23} : s = 197;
	{8'd217,8'd24} : s = 333;
	{8'd217,8'd25} : s = 331;
	{8'd217,8'd26} : s = 441;
	{8'd217,8'd27} : s = 327;
	{8'd217,8'd28} : s = 438;
	{8'd217,8'd29} : s = 437;
	{8'd217,8'd30} : s = 501;
	{8'd217,8'd31} : s = 316;
	{8'd217,8'd32} : s = 435;
	{8'd217,8'd33} : s = 430;
	{8'd217,8'd34} : s = 499;
	{8'd217,8'd35} : s = 429;
	{8'd217,8'd36} : s = 494;
	{8'd217,8'd37} : s = 493;
	{8'd217,8'd38} : s = 510;
	{8'd217,8'd39} : s = 1;
	{8'd217,8'd40} : s = 18;
	{8'd217,8'd41} : s = 17;
	{8'd217,8'd42} : s = 82;
	{8'd217,8'd43} : s = 12;
	{8'd217,8'd44} : s = 81;
	{8'd217,8'd45} : s = 76;
	{8'd217,8'd46} : s = 195;
	{8'd217,8'd47} : s = 10;
	{8'd217,8'd48} : s = 74;
	{8'd217,8'd49} : s = 73;
	{8'd217,8'd50} : s = 184;
	{8'd217,8'd51} : s = 70;
	{8'd217,8'd52} : s = 180;
	{8'd217,8'd53} : s = 178;
	{8'd217,8'd54} : s = 314;
	{8'd217,8'd55} : s = 9;
	{8'd217,8'd56} : s = 69;
	{8'd217,8'd57} : s = 67;
	{8'd217,8'd58} : s = 177;
	{8'd217,8'd59} : s = 56;
	{8'd217,8'd60} : s = 172;
	{8'd217,8'd61} : s = 170;
	{8'd217,8'd62} : s = 313;
	{8'd217,8'd63} : s = 52;
	{8'd217,8'd64} : s = 169;
	{8'd217,8'd65} : s = 166;
	{8'd217,8'd66} : s = 310;
	{8'd217,8'd67} : s = 165;
	{8'd217,8'd68} : s = 309;
	{8'd217,8'd69} : s = 307;
	{8'd217,8'd70} : s = 427;
	{8'd217,8'd71} : s = 6;
	{8'd217,8'd72} : s = 50;
	{8'd217,8'd73} : s = 49;
	{8'd217,8'd74} : s = 163;
	{8'd217,8'd75} : s = 44;
	{8'd217,8'd76} : s = 156;
	{8'd217,8'd77} : s = 154;
	{8'd217,8'd78} : s = 302;
	{8'd217,8'd79} : s = 42;
	{8'd217,8'd80} : s = 153;
	{8'd217,8'd81} : s = 150;
	{8'd217,8'd82} : s = 301;
	{8'd217,8'd83} : s = 149;
	{8'd217,8'd84} : s = 299;
	{8'd217,8'd85} : s = 295;
	{8'd217,8'd86} : s = 423;
	{8'd217,8'd87} : s = 41;
	{8'd217,8'd88} : s = 147;
	{8'd217,8'd89} : s = 142;
	{8'd217,8'd90} : s = 286;
	{8'd217,8'd91} : s = 141;
	{8'd217,8'd92} : s = 285;
	{8'd217,8'd93} : s = 283;
	{8'd217,8'd94} : s = 414;
	{8'd217,8'd95} : s = 139;
	{8'd217,8'd96} : s = 279;
	{8'd217,8'd97} : s = 271;
	{8'd217,8'd98} : s = 413;
	{8'd217,8'd99} : s = 248;
	{8'd217,8'd100} : s = 411;
	{8'd217,8'd101} : s = 407;
	{8'd217,8'd102} : s = 491;
	{8'd217,8'd103} : s = 5;
	{8'd217,8'd104} : s = 38;
	{8'd217,8'd105} : s = 37;
	{8'd217,8'd106} : s = 135;
	{8'd217,8'd107} : s = 35;
	{8'd217,8'd108} : s = 120;
	{8'd217,8'd109} : s = 116;
	{8'd217,8'd110} : s = 244;
	{8'd217,8'd111} : s = 28;
	{8'd217,8'd112} : s = 114;
	{8'd217,8'd113} : s = 113;
	{8'd217,8'd114} : s = 242;
	{8'd217,8'd115} : s = 108;
	{8'd217,8'd116} : s = 241;
	{8'd217,8'd117} : s = 236;
	{8'd217,8'd118} : s = 399;
	{8'd217,8'd119} : s = 26;
	{8'd217,8'd120} : s = 106;
	{8'd217,8'd121} : s = 105;
	{8'd217,8'd122} : s = 234;
	{8'd217,8'd123} : s = 102;
	{8'd217,8'd124} : s = 233;
	{8'd217,8'd125} : s = 230;
	{8'd217,8'd126} : s = 380;
	{8'd217,8'd127} : s = 101;
	{8'd217,8'd128} : s = 229;
	{8'd217,8'd129} : s = 227;
	{8'd217,8'd130} : s = 378;
	{8'd217,8'd131} : s = 220;
	{8'd217,8'd132} : s = 377;
	{8'd217,8'd133} : s = 374;
	{8'd217,8'd134} : s = 487;
	{8'd217,8'd135} : s = 25;
	{8'd217,8'd136} : s = 99;
	{8'd217,8'd137} : s = 92;
	{8'd217,8'd138} : s = 218;
	{8'd217,8'd139} : s = 90;
	{8'd217,8'd140} : s = 217;
	{8'd217,8'd141} : s = 214;
	{8'd217,8'd142} : s = 373;
	{8'd217,8'd143} : s = 89;
	{8'd217,8'd144} : s = 213;
	{8'd217,8'd145} : s = 211;
	{8'd217,8'd146} : s = 371;
	{8'd217,8'd147} : s = 206;
	{8'd217,8'd148} : s = 366;
	{8'd217,8'd149} : s = 365;
	{8'd217,8'd150} : s = 478;
	{8'd217,8'd151} : s = 86;
	{8'd217,8'd152} : s = 205;
	{8'd217,8'd153} : s = 203;
	{8'd217,8'd154} : s = 363;
	{8'd217,8'd155} : s = 199;
	{8'd217,8'd156} : s = 359;
	{8'd217,8'd157} : s = 350;
	{8'd217,8'd158} : s = 477;
	{8'd217,8'd159} : s = 188;
	{8'd217,8'd160} : s = 349;
	{8'd217,8'd161} : s = 347;
	{8'd217,8'd162} : s = 475;
	{8'd217,8'd163} : s = 343;
	{8'd217,8'd164} : s = 471;
	{8'd217,8'd165} : s = 463;
	{8'd217,8'd166} : s = 509;
	{8'd217,8'd167} : s = 3;
	{8'd217,8'd168} : s = 22;
	{8'd217,8'd169} : s = 21;
	{8'd217,8'd170} : s = 85;
	{8'd217,8'd171} : s = 19;
	{8'd217,8'd172} : s = 83;
	{8'd217,8'd173} : s = 78;
	{8'd217,8'd174} : s = 186;
	{8'd217,8'd175} : s = 14;
	{8'd217,8'd176} : s = 77;
	{8'd217,8'd177} : s = 75;
	{8'd217,8'd178} : s = 185;
	{8'd217,8'd179} : s = 71;
	{8'd217,8'd180} : s = 182;
	{8'd217,8'd181} : s = 181;
	{8'd217,8'd182} : s = 335;
	{8'd217,8'd183} : s = 13;
	{8'd217,8'd184} : s = 60;
	{8'd217,8'd185} : s = 58;
	{8'd217,8'd186} : s = 179;
	{8'd217,8'd187} : s = 57;
	{8'd217,8'd188} : s = 174;
	{8'd217,8'd189} : s = 173;
	{8'd217,8'd190} : s = 318;
	{8'd217,8'd191} : s = 54;
	{8'd217,8'd192} : s = 171;
	{8'd217,8'd193} : s = 167;
	{8'd217,8'd194} : s = 317;
	{8'd217,8'd195} : s = 158;
	{8'd217,8'd196} : s = 315;
	{8'd217,8'd197} : s = 311;
	{8'd217,8'd198} : s = 446;
	{8'd217,8'd199} : s = 11;
	{8'd217,8'd200} : s = 53;
	{8'd217,8'd201} : s = 51;
	{8'd217,8'd202} : s = 157;
	{8'd217,8'd203} : s = 46;
	{8'd217,8'd204} : s = 155;
	{8'd217,8'd205} : s = 151;
	{8'd217,8'd206} : s = 303;
	{8'd217,8'd207} : s = 45;
	{8'd217,8'd208} : s = 143;
	{8'd217,8'd209} : s = 124;
	{8'd217,8'd210} : s = 287;
	{8'd217,8'd211} : s = 122;
	{8'd217,8'd212} : s = 252;
	{8'd217,8'd213} : s = 250;
	{8'd217,8'd214} : s = 445;
	{8'd217,8'd215} : s = 43;
	{8'd217,8'd216} : s = 121;
	{8'd217,8'd217} : s = 118;
	{8'd217,8'd218} : s = 249;
	{8'd217,8'd219} : s = 117;
	{8'd217,8'd220} : s = 246;
	{8'd217,8'd221} : s = 245;
	{8'd217,8'd222} : s = 443;
	{8'd217,8'd223} : s = 115;
	{8'd217,8'd224} : s = 243;
	{8'd217,8'd225} : s = 238;
	{8'd217,8'd226} : s = 439;
	{8'd217,8'd227} : s = 237;
	{8'd217,8'd228} : s = 431;
	{8'd217,8'd229} : s = 415;
	{8'd217,8'd230} : s = 507;
	{8'd217,8'd231} : s = 7;
	{8'd217,8'd232} : s = 39;
	{8'd217,8'd233} : s = 30;
	{8'd217,8'd234} : s = 110;
	{8'd217,8'd235} : s = 29;
	{8'd217,8'd236} : s = 109;
	{8'd217,8'd237} : s = 107;
	{8'd217,8'd238} : s = 235;
	{8'd217,8'd239} : s = 27;
	{8'd217,8'd240} : s = 103;
	{8'd217,8'd241} : s = 94;
	{8'd217,8'd242} : s = 231;
	{8'd217,8'd243} : s = 93;
	{8'd217,8'd244} : s = 222;
	{8'd217,8'd245} : s = 221;
	{8'd217,8'd246} : s = 382;
	{8'd217,8'd247} : s = 23;
	{8'd217,8'd248} : s = 91;
	{8'd217,8'd249} : s = 87;
	{8'd217,8'd250} : s = 219;
	{8'd217,8'd251} : s = 79;
	{8'd217,8'd252} : s = 215;
	{8'd217,8'd253} : s = 207;
	{8'd217,8'd254} : s = 381;
	{8'd217,8'd255} : s = 62;
	{8'd218,8'd0} : s = 355;
	{8'd218,8'd1} : s = 467;
	{8'd218,8'd2} : s = 348;
	{8'd218,8'd3} : s = 462;
	{8'd218,8'd4} : s = 461;
	{8'd218,8'd5} : s = 505;
	{8'd218,8'd6} : s = 84;
	{8'd218,8'd7} : s = 204;
	{8'd218,8'd8} : s = 202;
	{8'd218,8'd9} : s = 346;
	{8'd218,8'd10} : s = 201;
	{8'd218,8'd11} : s = 345;
	{8'd218,8'd12} : s = 342;
	{8'd218,8'd13} : s = 459;
	{8'd218,8'd14} : s = 198;
	{8'd218,8'd15} : s = 341;
	{8'd218,8'd16} : s = 339;
	{8'd218,8'd17} : s = 455;
	{8'd218,8'd18} : s = 334;
	{8'd218,8'd19} : s = 444;
	{8'd218,8'd20} : s = 442;
	{8'd218,8'd21} : s = 502;
	{8'd218,8'd22} : s = 197;
	{8'd218,8'd23} : s = 333;
	{8'd218,8'd24} : s = 331;
	{8'd218,8'd25} : s = 441;
	{8'd218,8'd26} : s = 327;
	{8'd218,8'd27} : s = 438;
	{8'd218,8'd28} : s = 437;
	{8'd218,8'd29} : s = 501;
	{8'd218,8'd30} : s = 316;
	{8'd218,8'd31} : s = 435;
	{8'd218,8'd32} : s = 430;
	{8'd218,8'd33} : s = 499;
	{8'd218,8'd34} : s = 429;
	{8'd218,8'd35} : s = 494;
	{8'd218,8'd36} : s = 493;
	{8'd218,8'd37} : s = 510;
	{8'd218,8'd38} : s = 1;
	{8'd218,8'd39} : s = 18;
	{8'd218,8'd40} : s = 17;
	{8'd218,8'd41} : s = 82;
	{8'd218,8'd42} : s = 12;
	{8'd218,8'd43} : s = 81;
	{8'd218,8'd44} : s = 76;
	{8'd218,8'd45} : s = 195;
	{8'd218,8'd46} : s = 10;
	{8'd218,8'd47} : s = 74;
	{8'd218,8'd48} : s = 73;
	{8'd218,8'd49} : s = 184;
	{8'd218,8'd50} : s = 70;
	{8'd218,8'd51} : s = 180;
	{8'd218,8'd52} : s = 178;
	{8'd218,8'd53} : s = 314;
	{8'd218,8'd54} : s = 9;
	{8'd218,8'd55} : s = 69;
	{8'd218,8'd56} : s = 67;
	{8'd218,8'd57} : s = 177;
	{8'd218,8'd58} : s = 56;
	{8'd218,8'd59} : s = 172;
	{8'd218,8'd60} : s = 170;
	{8'd218,8'd61} : s = 313;
	{8'd218,8'd62} : s = 52;
	{8'd218,8'd63} : s = 169;
	{8'd218,8'd64} : s = 166;
	{8'd218,8'd65} : s = 310;
	{8'd218,8'd66} : s = 165;
	{8'd218,8'd67} : s = 309;
	{8'd218,8'd68} : s = 307;
	{8'd218,8'd69} : s = 427;
	{8'd218,8'd70} : s = 6;
	{8'd218,8'd71} : s = 50;
	{8'd218,8'd72} : s = 49;
	{8'd218,8'd73} : s = 163;
	{8'd218,8'd74} : s = 44;
	{8'd218,8'd75} : s = 156;
	{8'd218,8'd76} : s = 154;
	{8'd218,8'd77} : s = 302;
	{8'd218,8'd78} : s = 42;
	{8'd218,8'd79} : s = 153;
	{8'd218,8'd80} : s = 150;
	{8'd218,8'd81} : s = 301;
	{8'd218,8'd82} : s = 149;
	{8'd218,8'd83} : s = 299;
	{8'd218,8'd84} : s = 295;
	{8'd218,8'd85} : s = 423;
	{8'd218,8'd86} : s = 41;
	{8'd218,8'd87} : s = 147;
	{8'd218,8'd88} : s = 142;
	{8'd218,8'd89} : s = 286;
	{8'd218,8'd90} : s = 141;
	{8'd218,8'd91} : s = 285;
	{8'd218,8'd92} : s = 283;
	{8'd218,8'd93} : s = 414;
	{8'd218,8'd94} : s = 139;
	{8'd218,8'd95} : s = 279;
	{8'd218,8'd96} : s = 271;
	{8'd218,8'd97} : s = 413;
	{8'd218,8'd98} : s = 248;
	{8'd218,8'd99} : s = 411;
	{8'd218,8'd100} : s = 407;
	{8'd218,8'd101} : s = 491;
	{8'd218,8'd102} : s = 5;
	{8'd218,8'd103} : s = 38;
	{8'd218,8'd104} : s = 37;
	{8'd218,8'd105} : s = 135;
	{8'd218,8'd106} : s = 35;
	{8'd218,8'd107} : s = 120;
	{8'd218,8'd108} : s = 116;
	{8'd218,8'd109} : s = 244;
	{8'd218,8'd110} : s = 28;
	{8'd218,8'd111} : s = 114;
	{8'd218,8'd112} : s = 113;
	{8'd218,8'd113} : s = 242;
	{8'd218,8'd114} : s = 108;
	{8'd218,8'd115} : s = 241;
	{8'd218,8'd116} : s = 236;
	{8'd218,8'd117} : s = 399;
	{8'd218,8'd118} : s = 26;
	{8'd218,8'd119} : s = 106;
	{8'd218,8'd120} : s = 105;
	{8'd218,8'd121} : s = 234;
	{8'd218,8'd122} : s = 102;
	{8'd218,8'd123} : s = 233;
	{8'd218,8'd124} : s = 230;
	{8'd218,8'd125} : s = 380;
	{8'd218,8'd126} : s = 101;
	{8'd218,8'd127} : s = 229;
	{8'd218,8'd128} : s = 227;
	{8'd218,8'd129} : s = 378;
	{8'd218,8'd130} : s = 220;
	{8'd218,8'd131} : s = 377;
	{8'd218,8'd132} : s = 374;
	{8'd218,8'd133} : s = 487;
	{8'd218,8'd134} : s = 25;
	{8'd218,8'd135} : s = 99;
	{8'd218,8'd136} : s = 92;
	{8'd218,8'd137} : s = 218;
	{8'd218,8'd138} : s = 90;
	{8'd218,8'd139} : s = 217;
	{8'd218,8'd140} : s = 214;
	{8'd218,8'd141} : s = 373;
	{8'd218,8'd142} : s = 89;
	{8'd218,8'd143} : s = 213;
	{8'd218,8'd144} : s = 211;
	{8'd218,8'd145} : s = 371;
	{8'd218,8'd146} : s = 206;
	{8'd218,8'd147} : s = 366;
	{8'd218,8'd148} : s = 365;
	{8'd218,8'd149} : s = 478;
	{8'd218,8'd150} : s = 86;
	{8'd218,8'd151} : s = 205;
	{8'd218,8'd152} : s = 203;
	{8'd218,8'd153} : s = 363;
	{8'd218,8'd154} : s = 199;
	{8'd218,8'd155} : s = 359;
	{8'd218,8'd156} : s = 350;
	{8'd218,8'd157} : s = 477;
	{8'd218,8'd158} : s = 188;
	{8'd218,8'd159} : s = 349;
	{8'd218,8'd160} : s = 347;
	{8'd218,8'd161} : s = 475;
	{8'd218,8'd162} : s = 343;
	{8'd218,8'd163} : s = 471;
	{8'd218,8'd164} : s = 463;
	{8'd218,8'd165} : s = 509;
	{8'd218,8'd166} : s = 3;
	{8'd218,8'd167} : s = 22;
	{8'd218,8'd168} : s = 21;
	{8'd218,8'd169} : s = 85;
	{8'd218,8'd170} : s = 19;
	{8'd218,8'd171} : s = 83;
	{8'd218,8'd172} : s = 78;
	{8'd218,8'd173} : s = 186;
	{8'd218,8'd174} : s = 14;
	{8'd218,8'd175} : s = 77;
	{8'd218,8'd176} : s = 75;
	{8'd218,8'd177} : s = 185;
	{8'd218,8'd178} : s = 71;
	{8'd218,8'd179} : s = 182;
	{8'd218,8'd180} : s = 181;
	{8'd218,8'd181} : s = 335;
	{8'd218,8'd182} : s = 13;
	{8'd218,8'd183} : s = 60;
	{8'd218,8'd184} : s = 58;
	{8'd218,8'd185} : s = 179;
	{8'd218,8'd186} : s = 57;
	{8'd218,8'd187} : s = 174;
	{8'd218,8'd188} : s = 173;
	{8'd218,8'd189} : s = 318;
	{8'd218,8'd190} : s = 54;
	{8'd218,8'd191} : s = 171;
	{8'd218,8'd192} : s = 167;
	{8'd218,8'd193} : s = 317;
	{8'd218,8'd194} : s = 158;
	{8'd218,8'd195} : s = 315;
	{8'd218,8'd196} : s = 311;
	{8'd218,8'd197} : s = 446;
	{8'd218,8'd198} : s = 11;
	{8'd218,8'd199} : s = 53;
	{8'd218,8'd200} : s = 51;
	{8'd218,8'd201} : s = 157;
	{8'd218,8'd202} : s = 46;
	{8'd218,8'd203} : s = 155;
	{8'd218,8'd204} : s = 151;
	{8'd218,8'd205} : s = 303;
	{8'd218,8'd206} : s = 45;
	{8'd218,8'd207} : s = 143;
	{8'd218,8'd208} : s = 124;
	{8'd218,8'd209} : s = 287;
	{8'd218,8'd210} : s = 122;
	{8'd218,8'd211} : s = 252;
	{8'd218,8'd212} : s = 250;
	{8'd218,8'd213} : s = 445;
	{8'd218,8'd214} : s = 43;
	{8'd218,8'd215} : s = 121;
	{8'd218,8'd216} : s = 118;
	{8'd218,8'd217} : s = 249;
	{8'd218,8'd218} : s = 117;
	{8'd218,8'd219} : s = 246;
	{8'd218,8'd220} : s = 245;
	{8'd218,8'd221} : s = 443;
	{8'd218,8'd222} : s = 115;
	{8'd218,8'd223} : s = 243;
	{8'd218,8'd224} : s = 238;
	{8'd218,8'd225} : s = 439;
	{8'd218,8'd226} : s = 237;
	{8'd218,8'd227} : s = 431;
	{8'd218,8'd228} : s = 415;
	{8'd218,8'd229} : s = 507;
	{8'd218,8'd230} : s = 7;
	{8'd218,8'd231} : s = 39;
	{8'd218,8'd232} : s = 30;
	{8'd218,8'd233} : s = 110;
	{8'd218,8'd234} : s = 29;
	{8'd218,8'd235} : s = 109;
	{8'd218,8'd236} : s = 107;
	{8'd218,8'd237} : s = 235;
	{8'd218,8'd238} : s = 27;
	{8'd218,8'd239} : s = 103;
	{8'd218,8'd240} : s = 94;
	{8'd218,8'd241} : s = 231;
	{8'd218,8'd242} : s = 93;
	{8'd218,8'd243} : s = 222;
	{8'd218,8'd244} : s = 221;
	{8'd218,8'd245} : s = 382;
	{8'd218,8'd246} : s = 23;
	{8'd218,8'd247} : s = 91;
	{8'd218,8'd248} : s = 87;
	{8'd218,8'd249} : s = 219;
	{8'd218,8'd250} : s = 79;
	{8'd218,8'd251} : s = 215;
	{8'd218,8'd252} : s = 207;
	{8'd218,8'd253} : s = 381;
	{8'd218,8'd254} : s = 62;
	{8'd218,8'd255} : s = 190;
	{8'd219,8'd0} : s = 467;
	{8'd219,8'd1} : s = 348;
	{8'd219,8'd2} : s = 462;
	{8'd219,8'd3} : s = 461;
	{8'd219,8'd4} : s = 505;
	{8'd219,8'd5} : s = 84;
	{8'd219,8'd6} : s = 204;
	{8'd219,8'd7} : s = 202;
	{8'd219,8'd8} : s = 346;
	{8'd219,8'd9} : s = 201;
	{8'd219,8'd10} : s = 345;
	{8'd219,8'd11} : s = 342;
	{8'd219,8'd12} : s = 459;
	{8'd219,8'd13} : s = 198;
	{8'd219,8'd14} : s = 341;
	{8'd219,8'd15} : s = 339;
	{8'd219,8'd16} : s = 455;
	{8'd219,8'd17} : s = 334;
	{8'd219,8'd18} : s = 444;
	{8'd219,8'd19} : s = 442;
	{8'd219,8'd20} : s = 502;
	{8'd219,8'd21} : s = 197;
	{8'd219,8'd22} : s = 333;
	{8'd219,8'd23} : s = 331;
	{8'd219,8'd24} : s = 441;
	{8'd219,8'd25} : s = 327;
	{8'd219,8'd26} : s = 438;
	{8'd219,8'd27} : s = 437;
	{8'd219,8'd28} : s = 501;
	{8'd219,8'd29} : s = 316;
	{8'd219,8'd30} : s = 435;
	{8'd219,8'd31} : s = 430;
	{8'd219,8'd32} : s = 499;
	{8'd219,8'd33} : s = 429;
	{8'd219,8'd34} : s = 494;
	{8'd219,8'd35} : s = 493;
	{8'd219,8'd36} : s = 510;
	{8'd219,8'd37} : s = 1;
	{8'd219,8'd38} : s = 18;
	{8'd219,8'd39} : s = 17;
	{8'd219,8'd40} : s = 82;
	{8'd219,8'd41} : s = 12;
	{8'd219,8'd42} : s = 81;
	{8'd219,8'd43} : s = 76;
	{8'd219,8'd44} : s = 195;
	{8'd219,8'd45} : s = 10;
	{8'd219,8'd46} : s = 74;
	{8'd219,8'd47} : s = 73;
	{8'd219,8'd48} : s = 184;
	{8'd219,8'd49} : s = 70;
	{8'd219,8'd50} : s = 180;
	{8'd219,8'd51} : s = 178;
	{8'd219,8'd52} : s = 314;
	{8'd219,8'd53} : s = 9;
	{8'd219,8'd54} : s = 69;
	{8'd219,8'd55} : s = 67;
	{8'd219,8'd56} : s = 177;
	{8'd219,8'd57} : s = 56;
	{8'd219,8'd58} : s = 172;
	{8'd219,8'd59} : s = 170;
	{8'd219,8'd60} : s = 313;
	{8'd219,8'd61} : s = 52;
	{8'd219,8'd62} : s = 169;
	{8'd219,8'd63} : s = 166;
	{8'd219,8'd64} : s = 310;
	{8'd219,8'd65} : s = 165;
	{8'd219,8'd66} : s = 309;
	{8'd219,8'd67} : s = 307;
	{8'd219,8'd68} : s = 427;
	{8'd219,8'd69} : s = 6;
	{8'd219,8'd70} : s = 50;
	{8'd219,8'd71} : s = 49;
	{8'd219,8'd72} : s = 163;
	{8'd219,8'd73} : s = 44;
	{8'd219,8'd74} : s = 156;
	{8'd219,8'd75} : s = 154;
	{8'd219,8'd76} : s = 302;
	{8'd219,8'd77} : s = 42;
	{8'd219,8'd78} : s = 153;
	{8'd219,8'd79} : s = 150;
	{8'd219,8'd80} : s = 301;
	{8'd219,8'd81} : s = 149;
	{8'd219,8'd82} : s = 299;
	{8'd219,8'd83} : s = 295;
	{8'd219,8'd84} : s = 423;
	{8'd219,8'd85} : s = 41;
	{8'd219,8'd86} : s = 147;
	{8'd219,8'd87} : s = 142;
	{8'd219,8'd88} : s = 286;
	{8'd219,8'd89} : s = 141;
	{8'd219,8'd90} : s = 285;
	{8'd219,8'd91} : s = 283;
	{8'd219,8'd92} : s = 414;
	{8'd219,8'd93} : s = 139;
	{8'd219,8'd94} : s = 279;
	{8'd219,8'd95} : s = 271;
	{8'd219,8'd96} : s = 413;
	{8'd219,8'd97} : s = 248;
	{8'd219,8'd98} : s = 411;
	{8'd219,8'd99} : s = 407;
	{8'd219,8'd100} : s = 491;
	{8'd219,8'd101} : s = 5;
	{8'd219,8'd102} : s = 38;
	{8'd219,8'd103} : s = 37;
	{8'd219,8'd104} : s = 135;
	{8'd219,8'd105} : s = 35;
	{8'd219,8'd106} : s = 120;
	{8'd219,8'd107} : s = 116;
	{8'd219,8'd108} : s = 244;
	{8'd219,8'd109} : s = 28;
	{8'd219,8'd110} : s = 114;
	{8'd219,8'd111} : s = 113;
	{8'd219,8'd112} : s = 242;
	{8'd219,8'd113} : s = 108;
	{8'd219,8'd114} : s = 241;
	{8'd219,8'd115} : s = 236;
	{8'd219,8'd116} : s = 399;
	{8'd219,8'd117} : s = 26;
	{8'd219,8'd118} : s = 106;
	{8'd219,8'd119} : s = 105;
	{8'd219,8'd120} : s = 234;
	{8'd219,8'd121} : s = 102;
	{8'd219,8'd122} : s = 233;
	{8'd219,8'd123} : s = 230;
	{8'd219,8'd124} : s = 380;
	{8'd219,8'd125} : s = 101;
	{8'd219,8'd126} : s = 229;
	{8'd219,8'd127} : s = 227;
	{8'd219,8'd128} : s = 378;
	{8'd219,8'd129} : s = 220;
	{8'd219,8'd130} : s = 377;
	{8'd219,8'd131} : s = 374;
	{8'd219,8'd132} : s = 487;
	{8'd219,8'd133} : s = 25;
	{8'd219,8'd134} : s = 99;
	{8'd219,8'd135} : s = 92;
	{8'd219,8'd136} : s = 218;
	{8'd219,8'd137} : s = 90;
	{8'd219,8'd138} : s = 217;
	{8'd219,8'd139} : s = 214;
	{8'd219,8'd140} : s = 373;
	{8'd219,8'd141} : s = 89;
	{8'd219,8'd142} : s = 213;
	{8'd219,8'd143} : s = 211;
	{8'd219,8'd144} : s = 371;
	{8'd219,8'd145} : s = 206;
	{8'd219,8'd146} : s = 366;
	{8'd219,8'd147} : s = 365;
	{8'd219,8'd148} : s = 478;
	{8'd219,8'd149} : s = 86;
	{8'd219,8'd150} : s = 205;
	{8'd219,8'd151} : s = 203;
	{8'd219,8'd152} : s = 363;
	{8'd219,8'd153} : s = 199;
	{8'd219,8'd154} : s = 359;
	{8'd219,8'd155} : s = 350;
	{8'd219,8'd156} : s = 477;
	{8'd219,8'd157} : s = 188;
	{8'd219,8'd158} : s = 349;
	{8'd219,8'd159} : s = 347;
	{8'd219,8'd160} : s = 475;
	{8'd219,8'd161} : s = 343;
	{8'd219,8'd162} : s = 471;
	{8'd219,8'd163} : s = 463;
	{8'd219,8'd164} : s = 509;
	{8'd219,8'd165} : s = 3;
	{8'd219,8'd166} : s = 22;
	{8'd219,8'd167} : s = 21;
	{8'd219,8'd168} : s = 85;
	{8'd219,8'd169} : s = 19;
	{8'd219,8'd170} : s = 83;
	{8'd219,8'd171} : s = 78;
	{8'd219,8'd172} : s = 186;
	{8'd219,8'd173} : s = 14;
	{8'd219,8'd174} : s = 77;
	{8'd219,8'd175} : s = 75;
	{8'd219,8'd176} : s = 185;
	{8'd219,8'd177} : s = 71;
	{8'd219,8'd178} : s = 182;
	{8'd219,8'd179} : s = 181;
	{8'd219,8'd180} : s = 335;
	{8'd219,8'd181} : s = 13;
	{8'd219,8'd182} : s = 60;
	{8'd219,8'd183} : s = 58;
	{8'd219,8'd184} : s = 179;
	{8'd219,8'd185} : s = 57;
	{8'd219,8'd186} : s = 174;
	{8'd219,8'd187} : s = 173;
	{8'd219,8'd188} : s = 318;
	{8'd219,8'd189} : s = 54;
	{8'd219,8'd190} : s = 171;
	{8'd219,8'd191} : s = 167;
	{8'd219,8'd192} : s = 317;
	{8'd219,8'd193} : s = 158;
	{8'd219,8'd194} : s = 315;
	{8'd219,8'd195} : s = 311;
	{8'd219,8'd196} : s = 446;
	{8'd219,8'd197} : s = 11;
	{8'd219,8'd198} : s = 53;
	{8'd219,8'd199} : s = 51;
	{8'd219,8'd200} : s = 157;
	{8'd219,8'd201} : s = 46;
	{8'd219,8'd202} : s = 155;
	{8'd219,8'd203} : s = 151;
	{8'd219,8'd204} : s = 303;
	{8'd219,8'd205} : s = 45;
	{8'd219,8'd206} : s = 143;
	{8'd219,8'd207} : s = 124;
	{8'd219,8'd208} : s = 287;
	{8'd219,8'd209} : s = 122;
	{8'd219,8'd210} : s = 252;
	{8'd219,8'd211} : s = 250;
	{8'd219,8'd212} : s = 445;
	{8'd219,8'd213} : s = 43;
	{8'd219,8'd214} : s = 121;
	{8'd219,8'd215} : s = 118;
	{8'd219,8'd216} : s = 249;
	{8'd219,8'd217} : s = 117;
	{8'd219,8'd218} : s = 246;
	{8'd219,8'd219} : s = 245;
	{8'd219,8'd220} : s = 443;
	{8'd219,8'd221} : s = 115;
	{8'd219,8'd222} : s = 243;
	{8'd219,8'd223} : s = 238;
	{8'd219,8'd224} : s = 439;
	{8'd219,8'd225} : s = 237;
	{8'd219,8'd226} : s = 431;
	{8'd219,8'd227} : s = 415;
	{8'd219,8'd228} : s = 507;
	{8'd219,8'd229} : s = 7;
	{8'd219,8'd230} : s = 39;
	{8'd219,8'd231} : s = 30;
	{8'd219,8'd232} : s = 110;
	{8'd219,8'd233} : s = 29;
	{8'd219,8'd234} : s = 109;
	{8'd219,8'd235} : s = 107;
	{8'd219,8'd236} : s = 235;
	{8'd219,8'd237} : s = 27;
	{8'd219,8'd238} : s = 103;
	{8'd219,8'd239} : s = 94;
	{8'd219,8'd240} : s = 231;
	{8'd219,8'd241} : s = 93;
	{8'd219,8'd242} : s = 222;
	{8'd219,8'd243} : s = 221;
	{8'd219,8'd244} : s = 382;
	{8'd219,8'd245} : s = 23;
	{8'd219,8'd246} : s = 91;
	{8'd219,8'd247} : s = 87;
	{8'd219,8'd248} : s = 219;
	{8'd219,8'd249} : s = 79;
	{8'd219,8'd250} : s = 215;
	{8'd219,8'd251} : s = 207;
	{8'd219,8'd252} : s = 381;
	{8'd219,8'd253} : s = 62;
	{8'd219,8'd254} : s = 190;
	{8'd219,8'd255} : s = 189;
	{8'd220,8'd0} : s = 348;
	{8'd220,8'd1} : s = 462;
	{8'd220,8'd2} : s = 461;
	{8'd220,8'd3} : s = 505;
	{8'd220,8'd4} : s = 84;
	{8'd220,8'd5} : s = 204;
	{8'd220,8'd6} : s = 202;
	{8'd220,8'd7} : s = 346;
	{8'd220,8'd8} : s = 201;
	{8'd220,8'd9} : s = 345;
	{8'd220,8'd10} : s = 342;
	{8'd220,8'd11} : s = 459;
	{8'd220,8'd12} : s = 198;
	{8'd220,8'd13} : s = 341;
	{8'd220,8'd14} : s = 339;
	{8'd220,8'd15} : s = 455;
	{8'd220,8'd16} : s = 334;
	{8'd220,8'd17} : s = 444;
	{8'd220,8'd18} : s = 442;
	{8'd220,8'd19} : s = 502;
	{8'd220,8'd20} : s = 197;
	{8'd220,8'd21} : s = 333;
	{8'd220,8'd22} : s = 331;
	{8'd220,8'd23} : s = 441;
	{8'd220,8'd24} : s = 327;
	{8'd220,8'd25} : s = 438;
	{8'd220,8'd26} : s = 437;
	{8'd220,8'd27} : s = 501;
	{8'd220,8'd28} : s = 316;
	{8'd220,8'd29} : s = 435;
	{8'd220,8'd30} : s = 430;
	{8'd220,8'd31} : s = 499;
	{8'd220,8'd32} : s = 429;
	{8'd220,8'd33} : s = 494;
	{8'd220,8'd34} : s = 493;
	{8'd220,8'd35} : s = 510;
	{8'd220,8'd36} : s = 1;
	{8'd220,8'd37} : s = 18;
	{8'd220,8'd38} : s = 17;
	{8'd220,8'd39} : s = 82;
	{8'd220,8'd40} : s = 12;
	{8'd220,8'd41} : s = 81;
	{8'd220,8'd42} : s = 76;
	{8'd220,8'd43} : s = 195;
	{8'd220,8'd44} : s = 10;
	{8'd220,8'd45} : s = 74;
	{8'd220,8'd46} : s = 73;
	{8'd220,8'd47} : s = 184;
	{8'd220,8'd48} : s = 70;
	{8'd220,8'd49} : s = 180;
	{8'd220,8'd50} : s = 178;
	{8'd220,8'd51} : s = 314;
	{8'd220,8'd52} : s = 9;
	{8'd220,8'd53} : s = 69;
	{8'd220,8'd54} : s = 67;
	{8'd220,8'd55} : s = 177;
	{8'd220,8'd56} : s = 56;
	{8'd220,8'd57} : s = 172;
	{8'd220,8'd58} : s = 170;
	{8'd220,8'd59} : s = 313;
	{8'd220,8'd60} : s = 52;
	{8'd220,8'd61} : s = 169;
	{8'd220,8'd62} : s = 166;
	{8'd220,8'd63} : s = 310;
	{8'd220,8'd64} : s = 165;
	{8'd220,8'd65} : s = 309;
	{8'd220,8'd66} : s = 307;
	{8'd220,8'd67} : s = 427;
	{8'd220,8'd68} : s = 6;
	{8'd220,8'd69} : s = 50;
	{8'd220,8'd70} : s = 49;
	{8'd220,8'd71} : s = 163;
	{8'd220,8'd72} : s = 44;
	{8'd220,8'd73} : s = 156;
	{8'd220,8'd74} : s = 154;
	{8'd220,8'd75} : s = 302;
	{8'd220,8'd76} : s = 42;
	{8'd220,8'd77} : s = 153;
	{8'd220,8'd78} : s = 150;
	{8'd220,8'd79} : s = 301;
	{8'd220,8'd80} : s = 149;
	{8'd220,8'd81} : s = 299;
	{8'd220,8'd82} : s = 295;
	{8'd220,8'd83} : s = 423;
	{8'd220,8'd84} : s = 41;
	{8'd220,8'd85} : s = 147;
	{8'd220,8'd86} : s = 142;
	{8'd220,8'd87} : s = 286;
	{8'd220,8'd88} : s = 141;
	{8'd220,8'd89} : s = 285;
	{8'd220,8'd90} : s = 283;
	{8'd220,8'd91} : s = 414;
	{8'd220,8'd92} : s = 139;
	{8'd220,8'd93} : s = 279;
	{8'd220,8'd94} : s = 271;
	{8'd220,8'd95} : s = 413;
	{8'd220,8'd96} : s = 248;
	{8'd220,8'd97} : s = 411;
	{8'd220,8'd98} : s = 407;
	{8'd220,8'd99} : s = 491;
	{8'd220,8'd100} : s = 5;
	{8'd220,8'd101} : s = 38;
	{8'd220,8'd102} : s = 37;
	{8'd220,8'd103} : s = 135;
	{8'd220,8'd104} : s = 35;
	{8'd220,8'd105} : s = 120;
	{8'd220,8'd106} : s = 116;
	{8'd220,8'd107} : s = 244;
	{8'd220,8'd108} : s = 28;
	{8'd220,8'd109} : s = 114;
	{8'd220,8'd110} : s = 113;
	{8'd220,8'd111} : s = 242;
	{8'd220,8'd112} : s = 108;
	{8'd220,8'd113} : s = 241;
	{8'd220,8'd114} : s = 236;
	{8'd220,8'd115} : s = 399;
	{8'd220,8'd116} : s = 26;
	{8'd220,8'd117} : s = 106;
	{8'd220,8'd118} : s = 105;
	{8'd220,8'd119} : s = 234;
	{8'd220,8'd120} : s = 102;
	{8'd220,8'd121} : s = 233;
	{8'd220,8'd122} : s = 230;
	{8'd220,8'd123} : s = 380;
	{8'd220,8'd124} : s = 101;
	{8'd220,8'd125} : s = 229;
	{8'd220,8'd126} : s = 227;
	{8'd220,8'd127} : s = 378;
	{8'd220,8'd128} : s = 220;
	{8'd220,8'd129} : s = 377;
	{8'd220,8'd130} : s = 374;
	{8'd220,8'd131} : s = 487;
	{8'd220,8'd132} : s = 25;
	{8'd220,8'd133} : s = 99;
	{8'd220,8'd134} : s = 92;
	{8'd220,8'd135} : s = 218;
	{8'd220,8'd136} : s = 90;
	{8'd220,8'd137} : s = 217;
	{8'd220,8'd138} : s = 214;
	{8'd220,8'd139} : s = 373;
	{8'd220,8'd140} : s = 89;
	{8'd220,8'd141} : s = 213;
	{8'd220,8'd142} : s = 211;
	{8'd220,8'd143} : s = 371;
	{8'd220,8'd144} : s = 206;
	{8'd220,8'd145} : s = 366;
	{8'd220,8'd146} : s = 365;
	{8'd220,8'd147} : s = 478;
	{8'd220,8'd148} : s = 86;
	{8'd220,8'd149} : s = 205;
	{8'd220,8'd150} : s = 203;
	{8'd220,8'd151} : s = 363;
	{8'd220,8'd152} : s = 199;
	{8'd220,8'd153} : s = 359;
	{8'd220,8'd154} : s = 350;
	{8'd220,8'd155} : s = 477;
	{8'd220,8'd156} : s = 188;
	{8'd220,8'd157} : s = 349;
	{8'd220,8'd158} : s = 347;
	{8'd220,8'd159} : s = 475;
	{8'd220,8'd160} : s = 343;
	{8'd220,8'd161} : s = 471;
	{8'd220,8'd162} : s = 463;
	{8'd220,8'd163} : s = 509;
	{8'd220,8'd164} : s = 3;
	{8'd220,8'd165} : s = 22;
	{8'd220,8'd166} : s = 21;
	{8'd220,8'd167} : s = 85;
	{8'd220,8'd168} : s = 19;
	{8'd220,8'd169} : s = 83;
	{8'd220,8'd170} : s = 78;
	{8'd220,8'd171} : s = 186;
	{8'd220,8'd172} : s = 14;
	{8'd220,8'd173} : s = 77;
	{8'd220,8'd174} : s = 75;
	{8'd220,8'd175} : s = 185;
	{8'd220,8'd176} : s = 71;
	{8'd220,8'd177} : s = 182;
	{8'd220,8'd178} : s = 181;
	{8'd220,8'd179} : s = 335;
	{8'd220,8'd180} : s = 13;
	{8'd220,8'd181} : s = 60;
	{8'd220,8'd182} : s = 58;
	{8'd220,8'd183} : s = 179;
	{8'd220,8'd184} : s = 57;
	{8'd220,8'd185} : s = 174;
	{8'd220,8'd186} : s = 173;
	{8'd220,8'd187} : s = 318;
	{8'd220,8'd188} : s = 54;
	{8'd220,8'd189} : s = 171;
	{8'd220,8'd190} : s = 167;
	{8'd220,8'd191} : s = 317;
	{8'd220,8'd192} : s = 158;
	{8'd220,8'd193} : s = 315;
	{8'd220,8'd194} : s = 311;
	{8'd220,8'd195} : s = 446;
	{8'd220,8'd196} : s = 11;
	{8'd220,8'd197} : s = 53;
	{8'd220,8'd198} : s = 51;
	{8'd220,8'd199} : s = 157;
	{8'd220,8'd200} : s = 46;
	{8'd220,8'd201} : s = 155;
	{8'd220,8'd202} : s = 151;
	{8'd220,8'd203} : s = 303;
	{8'd220,8'd204} : s = 45;
	{8'd220,8'd205} : s = 143;
	{8'd220,8'd206} : s = 124;
	{8'd220,8'd207} : s = 287;
	{8'd220,8'd208} : s = 122;
	{8'd220,8'd209} : s = 252;
	{8'd220,8'd210} : s = 250;
	{8'd220,8'd211} : s = 445;
	{8'd220,8'd212} : s = 43;
	{8'd220,8'd213} : s = 121;
	{8'd220,8'd214} : s = 118;
	{8'd220,8'd215} : s = 249;
	{8'd220,8'd216} : s = 117;
	{8'd220,8'd217} : s = 246;
	{8'd220,8'd218} : s = 245;
	{8'd220,8'd219} : s = 443;
	{8'd220,8'd220} : s = 115;
	{8'd220,8'd221} : s = 243;
	{8'd220,8'd222} : s = 238;
	{8'd220,8'd223} : s = 439;
	{8'd220,8'd224} : s = 237;
	{8'd220,8'd225} : s = 431;
	{8'd220,8'd226} : s = 415;
	{8'd220,8'd227} : s = 507;
	{8'd220,8'd228} : s = 7;
	{8'd220,8'd229} : s = 39;
	{8'd220,8'd230} : s = 30;
	{8'd220,8'd231} : s = 110;
	{8'd220,8'd232} : s = 29;
	{8'd220,8'd233} : s = 109;
	{8'd220,8'd234} : s = 107;
	{8'd220,8'd235} : s = 235;
	{8'd220,8'd236} : s = 27;
	{8'd220,8'd237} : s = 103;
	{8'd220,8'd238} : s = 94;
	{8'd220,8'd239} : s = 231;
	{8'd220,8'd240} : s = 93;
	{8'd220,8'd241} : s = 222;
	{8'd220,8'd242} : s = 221;
	{8'd220,8'd243} : s = 382;
	{8'd220,8'd244} : s = 23;
	{8'd220,8'd245} : s = 91;
	{8'd220,8'd246} : s = 87;
	{8'd220,8'd247} : s = 219;
	{8'd220,8'd248} : s = 79;
	{8'd220,8'd249} : s = 215;
	{8'd220,8'd250} : s = 207;
	{8'd220,8'd251} : s = 381;
	{8'd220,8'd252} : s = 62;
	{8'd220,8'd253} : s = 190;
	{8'd220,8'd254} : s = 189;
	{8'd220,8'd255} : s = 379;
	{8'd221,8'd0} : s = 462;
	{8'd221,8'd1} : s = 461;
	{8'd221,8'd2} : s = 505;
	{8'd221,8'd3} : s = 84;
	{8'd221,8'd4} : s = 204;
	{8'd221,8'd5} : s = 202;
	{8'd221,8'd6} : s = 346;
	{8'd221,8'd7} : s = 201;
	{8'd221,8'd8} : s = 345;
	{8'd221,8'd9} : s = 342;
	{8'd221,8'd10} : s = 459;
	{8'd221,8'd11} : s = 198;
	{8'd221,8'd12} : s = 341;
	{8'd221,8'd13} : s = 339;
	{8'd221,8'd14} : s = 455;
	{8'd221,8'd15} : s = 334;
	{8'd221,8'd16} : s = 444;
	{8'd221,8'd17} : s = 442;
	{8'd221,8'd18} : s = 502;
	{8'd221,8'd19} : s = 197;
	{8'd221,8'd20} : s = 333;
	{8'd221,8'd21} : s = 331;
	{8'd221,8'd22} : s = 441;
	{8'd221,8'd23} : s = 327;
	{8'd221,8'd24} : s = 438;
	{8'd221,8'd25} : s = 437;
	{8'd221,8'd26} : s = 501;
	{8'd221,8'd27} : s = 316;
	{8'd221,8'd28} : s = 435;
	{8'd221,8'd29} : s = 430;
	{8'd221,8'd30} : s = 499;
	{8'd221,8'd31} : s = 429;
	{8'd221,8'd32} : s = 494;
	{8'd221,8'd33} : s = 493;
	{8'd221,8'd34} : s = 510;
	{8'd221,8'd35} : s = 1;
	{8'd221,8'd36} : s = 18;
	{8'd221,8'd37} : s = 17;
	{8'd221,8'd38} : s = 82;
	{8'd221,8'd39} : s = 12;
	{8'd221,8'd40} : s = 81;
	{8'd221,8'd41} : s = 76;
	{8'd221,8'd42} : s = 195;
	{8'd221,8'd43} : s = 10;
	{8'd221,8'd44} : s = 74;
	{8'd221,8'd45} : s = 73;
	{8'd221,8'd46} : s = 184;
	{8'd221,8'd47} : s = 70;
	{8'd221,8'd48} : s = 180;
	{8'd221,8'd49} : s = 178;
	{8'd221,8'd50} : s = 314;
	{8'd221,8'd51} : s = 9;
	{8'd221,8'd52} : s = 69;
	{8'd221,8'd53} : s = 67;
	{8'd221,8'd54} : s = 177;
	{8'd221,8'd55} : s = 56;
	{8'd221,8'd56} : s = 172;
	{8'd221,8'd57} : s = 170;
	{8'd221,8'd58} : s = 313;
	{8'd221,8'd59} : s = 52;
	{8'd221,8'd60} : s = 169;
	{8'd221,8'd61} : s = 166;
	{8'd221,8'd62} : s = 310;
	{8'd221,8'd63} : s = 165;
	{8'd221,8'd64} : s = 309;
	{8'd221,8'd65} : s = 307;
	{8'd221,8'd66} : s = 427;
	{8'd221,8'd67} : s = 6;
	{8'd221,8'd68} : s = 50;
	{8'd221,8'd69} : s = 49;
	{8'd221,8'd70} : s = 163;
	{8'd221,8'd71} : s = 44;
	{8'd221,8'd72} : s = 156;
	{8'd221,8'd73} : s = 154;
	{8'd221,8'd74} : s = 302;
	{8'd221,8'd75} : s = 42;
	{8'd221,8'd76} : s = 153;
	{8'd221,8'd77} : s = 150;
	{8'd221,8'd78} : s = 301;
	{8'd221,8'd79} : s = 149;
	{8'd221,8'd80} : s = 299;
	{8'd221,8'd81} : s = 295;
	{8'd221,8'd82} : s = 423;
	{8'd221,8'd83} : s = 41;
	{8'd221,8'd84} : s = 147;
	{8'd221,8'd85} : s = 142;
	{8'd221,8'd86} : s = 286;
	{8'd221,8'd87} : s = 141;
	{8'd221,8'd88} : s = 285;
	{8'd221,8'd89} : s = 283;
	{8'd221,8'd90} : s = 414;
	{8'd221,8'd91} : s = 139;
	{8'd221,8'd92} : s = 279;
	{8'd221,8'd93} : s = 271;
	{8'd221,8'd94} : s = 413;
	{8'd221,8'd95} : s = 248;
	{8'd221,8'd96} : s = 411;
	{8'd221,8'd97} : s = 407;
	{8'd221,8'd98} : s = 491;
	{8'd221,8'd99} : s = 5;
	{8'd221,8'd100} : s = 38;
	{8'd221,8'd101} : s = 37;
	{8'd221,8'd102} : s = 135;
	{8'd221,8'd103} : s = 35;
	{8'd221,8'd104} : s = 120;
	{8'd221,8'd105} : s = 116;
	{8'd221,8'd106} : s = 244;
	{8'd221,8'd107} : s = 28;
	{8'd221,8'd108} : s = 114;
	{8'd221,8'd109} : s = 113;
	{8'd221,8'd110} : s = 242;
	{8'd221,8'd111} : s = 108;
	{8'd221,8'd112} : s = 241;
	{8'd221,8'd113} : s = 236;
	{8'd221,8'd114} : s = 399;
	{8'd221,8'd115} : s = 26;
	{8'd221,8'd116} : s = 106;
	{8'd221,8'd117} : s = 105;
	{8'd221,8'd118} : s = 234;
	{8'd221,8'd119} : s = 102;
	{8'd221,8'd120} : s = 233;
	{8'd221,8'd121} : s = 230;
	{8'd221,8'd122} : s = 380;
	{8'd221,8'd123} : s = 101;
	{8'd221,8'd124} : s = 229;
	{8'd221,8'd125} : s = 227;
	{8'd221,8'd126} : s = 378;
	{8'd221,8'd127} : s = 220;
	{8'd221,8'd128} : s = 377;
	{8'd221,8'd129} : s = 374;
	{8'd221,8'd130} : s = 487;
	{8'd221,8'd131} : s = 25;
	{8'd221,8'd132} : s = 99;
	{8'd221,8'd133} : s = 92;
	{8'd221,8'd134} : s = 218;
	{8'd221,8'd135} : s = 90;
	{8'd221,8'd136} : s = 217;
	{8'd221,8'd137} : s = 214;
	{8'd221,8'd138} : s = 373;
	{8'd221,8'd139} : s = 89;
	{8'd221,8'd140} : s = 213;
	{8'd221,8'd141} : s = 211;
	{8'd221,8'd142} : s = 371;
	{8'd221,8'd143} : s = 206;
	{8'd221,8'd144} : s = 366;
	{8'd221,8'd145} : s = 365;
	{8'd221,8'd146} : s = 478;
	{8'd221,8'd147} : s = 86;
	{8'd221,8'd148} : s = 205;
	{8'd221,8'd149} : s = 203;
	{8'd221,8'd150} : s = 363;
	{8'd221,8'd151} : s = 199;
	{8'd221,8'd152} : s = 359;
	{8'd221,8'd153} : s = 350;
	{8'd221,8'd154} : s = 477;
	{8'd221,8'd155} : s = 188;
	{8'd221,8'd156} : s = 349;
	{8'd221,8'd157} : s = 347;
	{8'd221,8'd158} : s = 475;
	{8'd221,8'd159} : s = 343;
	{8'd221,8'd160} : s = 471;
	{8'd221,8'd161} : s = 463;
	{8'd221,8'd162} : s = 509;
	{8'd221,8'd163} : s = 3;
	{8'd221,8'd164} : s = 22;
	{8'd221,8'd165} : s = 21;
	{8'd221,8'd166} : s = 85;
	{8'd221,8'd167} : s = 19;
	{8'd221,8'd168} : s = 83;
	{8'd221,8'd169} : s = 78;
	{8'd221,8'd170} : s = 186;
	{8'd221,8'd171} : s = 14;
	{8'd221,8'd172} : s = 77;
	{8'd221,8'd173} : s = 75;
	{8'd221,8'd174} : s = 185;
	{8'd221,8'd175} : s = 71;
	{8'd221,8'd176} : s = 182;
	{8'd221,8'd177} : s = 181;
	{8'd221,8'd178} : s = 335;
	{8'd221,8'd179} : s = 13;
	{8'd221,8'd180} : s = 60;
	{8'd221,8'd181} : s = 58;
	{8'd221,8'd182} : s = 179;
	{8'd221,8'd183} : s = 57;
	{8'd221,8'd184} : s = 174;
	{8'd221,8'd185} : s = 173;
	{8'd221,8'd186} : s = 318;
	{8'd221,8'd187} : s = 54;
	{8'd221,8'd188} : s = 171;
	{8'd221,8'd189} : s = 167;
	{8'd221,8'd190} : s = 317;
	{8'd221,8'd191} : s = 158;
	{8'd221,8'd192} : s = 315;
	{8'd221,8'd193} : s = 311;
	{8'd221,8'd194} : s = 446;
	{8'd221,8'd195} : s = 11;
	{8'd221,8'd196} : s = 53;
	{8'd221,8'd197} : s = 51;
	{8'd221,8'd198} : s = 157;
	{8'd221,8'd199} : s = 46;
	{8'd221,8'd200} : s = 155;
	{8'd221,8'd201} : s = 151;
	{8'd221,8'd202} : s = 303;
	{8'd221,8'd203} : s = 45;
	{8'd221,8'd204} : s = 143;
	{8'd221,8'd205} : s = 124;
	{8'd221,8'd206} : s = 287;
	{8'd221,8'd207} : s = 122;
	{8'd221,8'd208} : s = 252;
	{8'd221,8'd209} : s = 250;
	{8'd221,8'd210} : s = 445;
	{8'd221,8'd211} : s = 43;
	{8'd221,8'd212} : s = 121;
	{8'd221,8'd213} : s = 118;
	{8'd221,8'd214} : s = 249;
	{8'd221,8'd215} : s = 117;
	{8'd221,8'd216} : s = 246;
	{8'd221,8'd217} : s = 245;
	{8'd221,8'd218} : s = 443;
	{8'd221,8'd219} : s = 115;
	{8'd221,8'd220} : s = 243;
	{8'd221,8'd221} : s = 238;
	{8'd221,8'd222} : s = 439;
	{8'd221,8'd223} : s = 237;
	{8'd221,8'd224} : s = 431;
	{8'd221,8'd225} : s = 415;
	{8'd221,8'd226} : s = 507;
	{8'd221,8'd227} : s = 7;
	{8'd221,8'd228} : s = 39;
	{8'd221,8'd229} : s = 30;
	{8'd221,8'd230} : s = 110;
	{8'd221,8'd231} : s = 29;
	{8'd221,8'd232} : s = 109;
	{8'd221,8'd233} : s = 107;
	{8'd221,8'd234} : s = 235;
	{8'd221,8'd235} : s = 27;
	{8'd221,8'd236} : s = 103;
	{8'd221,8'd237} : s = 94;
	{8'd221,8'd238} : s = 231;
	{8'd221,8'd239} : s = 93;
	{8'd221,8'd240} : s = 222;
	{8'd221,8'd241} : s = 221;
	{8'd221,8'd242} : s = 382;
	{8'd221,8'd243} : s = 23;
	{8'd221,8'd244} : s = 91;
	{8'd221,8'd245} : s = 87;
	{8'd221,8'd246} : s = 219;
	{8'd221,8'd247} : s = 79;
	{8'd221,8'd248} : s = 215;
	{8'd221,8'd249} : s = 207;
	{8'd221,8'd250} : s = 381;
	{8'd221,8'd251} : s = 62;
	{8'd221,8'd252} : s = 190;
	{8'd221,8'd253} : s = 189;
	{8'd221,8'd254} : s = 379;
	{8'd221,8'd255} : s = 187;
	{8'd222,8'd0} : s = 461;
	{8'd222,8'd1} : s = 505;
	{8'd222,8'd2} : s = 84;
	{8'd222,8'd3} : s = 204;
	{8'd222,8'd4} : s = 202;
	{8'd222,8'd5} : s = 346;
	{8'd222,8'd6} : s = 201;
	{8'd222,8'd7} : s = 345;
	{8'd222,8'd8} : s = 342;
	{8'd222,8'd9} : s = 459;
	{8'd222,8'd10} : s = 198;
	{8'd222,8'd11} : s = 341;
	{8'd222,8'd12} : s = 339;
	{8'd222,8'd13} : s = 455;
	{8'd222,8'd14} : s = 334;
	{8'd222,8'd15} : s = 444;
	{8'd222,8'd16} : s = 442;
	{8'd222,8'd17} : s = 502;
	{8'd222,8'd18} : s = 197;
	{8'd222,8'd19} : s = 333;
	{8'd222,8'd20} : s = 331;
	{8'd222,8'd21} : s = 441;
	{8'd222,8'd22} : s = 327;
	{8'd222,8'd23} : s = 438;
	{8'd222,8'd24} : s = 437;
	{8'd222,8'd25} : s = 501;
	{8'd222,8'd26} : s = 316;
	{8'd222,8'd27} : s = 435;
	{8'd222,8'd28} : s = 430;
	{8'd222,8'd29} : s = 499;
	{8'd222,8'd30} : s = 429;
	{8'd222,8'd31} : s = 494;
	{8'd222,8'd32} : s = 493;
	{8'd222,8'd33} : s = 510;
	{8'd222,8'd34} : s = 1;
	{8'd222,8'd35} : s = 18;
	{8'd222,8'd36} : s = 17;
	{8'd222,8'd37} : s = 82;
	{8'd222,8'd38} : s = 12;
	{8'd222,8'd39} : s = 81;
	{8'd222,8'd40} : s = 76;
	{8'd222,8'd41} : s = 195;
	{8'd222,8'd42} : s = 10;
	{8'd222,8'd43} : s = 74;
	{8'd222,8'd44} : s = 73;
	{8'd222,8'd45} : s = 184;
	{8'd222,8'd46} : s = 70;
	{8'd222,8'd47} : s = 180;
	{8'd222,8'd48} : s = 178;
	{8'd222,8'd49} : s = 314;
	{8'd222,8'd50} : s = 9;
	{8'd222,8'd51} : s = 69;
	{8'd222,8'd52} : s = 67;
	{8'd222,8'd53} : s = 177;
	{8'd222,8'd54} : s = 56;
	{8'd222,8'd55} : s = 172;
	{8'd222,8'd56} : s = 170;
	{8'd222,8'd57} : s = 313;
	{8'd222,8'd58} : s = 52;
	{8'd222,8'd59} : s = 169;
	{8'd222,8'd60} : s = 166;
	{8'd222,8'd61} : s = 310;
	{8'd222,8'd62} : s = 165;
	{8'd222,8'd63} : s = 309;
	{8'd222,8'd64} : s = 307;
	{8'd222,8'd65} : s = 427;
	{8'd222,8'd66} : s = 6;
	{8'd222,8'd67} : s = 50;
	{8'd222,8'd68} : s = 49;
	{8'd222,8'd69} : s = 163;
	{8'd222,8'd70} : s = 44;
	{8'd222,8'd71} : s = 156;
	{8'd222,8'd72} : s = 154;
	{8'd222,8'd73} : s = 302;
	{8'd222,8'd74} : s = 42;
	{8'd222,8'd75} : s = 153;
	{8'd222,8'd76} : s = 150;
	{8'd222,8'd77} : s = 301;
	{8'd222,8'd78} : s = 149;
	{8'd222,8'd79} : s = 299;
	{8'd222,8'd80} : s = 295;
	{8'd222,8'd81} : s = 423;
	{8'd222,8'd82} : s = 41;
	{8'd222,8'd83} : s = 147;
	{8'd222,8'd84} : s = 142;
	{8'd222,8'd85} : s = 286;
	{8'd222,8'd86} : s = 141;
	{8'd222,8'd87} : s = 285;
	{8'd222,8'd88} : s = 283;
	{8'd222,8'd89} : s = 414;
	{8'd222,8'd90} : s = 139;
	{8'd222,8'd91} : s = 279;
	{8'd222,8'd92} : s = 271;
	{8'd222,8'd93} : s = 413;
	{8'd222,8'd94} : s = 248;
	{8'd222,8'd95} : s = 411;
	{8'd222,8'd96} : s = 407;
	{8'd222,8'd97} : s = 491;
	{8'd222,8'd98} : s = 5;
	{8'd222,8'd99} : s = 38;
	{8'd222,8'd100} : s = 37;
	{8'd222,8'd101} : s = 135;
	{8'd222,8'd102} : s = 35;
	{8'd222,8'd103} : s = 120;
	{8'd222,8'd104} : s = 116;
	{8'd222,8'd105} : s = 244;
	{8'd222,8'd106} : s = 28;
	{8'd222,8'd107} : s = 114;
	{8'd222,8'd108} : s = 113;
	{8'd222,8'd109} : s = 242;
	{8'd222,8'd110} : s = 108;
	{8'd222,8'd111} : s = 241;
	{8'd222,8'd112} : s = 236;
	{8'd222,8'd113} : s = 399;
	{8'd222,8'd114} : s = 26;
	{8'd222,8'd115} : s = 106;
	{8'd222,8'd116} : s = 105;
	{8'd222,8'd117} : s = 234;
	{8'd222,8'd118} : s = 102;
	{8'd222,8'd119} : s = 233;
	{8'd222,8'd120} : s = 230;
	{8'd222,8'd121} : s = 380;
	{8'd222,8'd122} : s = 101;
	{8'd222,8'd123} : s = 229;
	{8'd222,8'd124} : s = 227;
	{8'd222,8'd125} : s = 378;
	{8'd222,8'd126} : s = 220;
	{8'd222,8'd127} : s = 377;
	{8'd222,8'd128} : s = 374;
	{8'd222,8'd129} : s = 487;
	{8'd222,8'd130} : s = 25;
	{8'd222,8'd131} : s = 99;
	{8'd222,8'd132} : s = 92;
	{8'd222,8'd133} : s = 218;
	{8'd222,8'd134} : s = 90;
	{8'd222,8'd135} : s = 217;
	{8'd222,8'd136} : s = 214;
	{8'd222,8'd137} : s = 373;
	{8'd222,8'd138} : s = 89;
	{8'd222,8'd139} : s = 213;
	{8'd222,8'd140} : s = 211;
	{8'd222,8'd141} : s = 371;
	{8'd222,8'd142} : s = 206;
	{8'd222,8'd143} : s = 366;
	{8'd222,8'd144} : s = 365;
	{8'd222,8'd145} : s = 478;
	{8'd222,8'd146} : s = 86;
	{8'd222,8'd147} : s = 205;
	{8'd222,8'd148} : s = 203;
	{8'd222,8'd149} : s = 363;
	{8'd222,8'd150} : s = 199;
	{8'd222,8'd151} : s = 359;
	{8'd222,8'd152} : s = 350;
	{8'd222,8'd153} : s = 477;
	{8'd222,8'd154} : s = 188;
	{8'd222,8'd155} : s = 349;
	{8'd222,8'd156} : s = 347;
	{8'd222,8'd157} : s = 475;
	{8'd222,8'd158} : s = 343;
	{8'd222,8'd159} : s = 471;
	{8'd222,8'd160} : s = 463;
	{8'd222,8'd161} : s = 509;
	{8'd222,8'd162} : s = 3;
	{8'd222,8'd163} : s = 22;
	{8'd222,8'd164} : s = 21;
	{8'd222,8'd165} : s = 85;
	{8'd222,8'd166} : s = 19;
	{8'd222,8'd167} : s = 83;
	{8'd222,8'd168} : s = 78;
	{8'd222,8'd169} : s = 186;
	{8'd222,8'd170} : s = 14;
	{8'd222,8'd171} : s = 77;
	{8'd222,8'd172} : s = 75;
	{8'd222,8'd173} : s = 185;
	{8'd222,8'd174} : s = 71;
	{8'd222,8'd175} : s = 182;
	{8'd222,8'd176} : s = 181;
	{8'd222,8'd177} : s = 335;
	{8'd222,8'd178} : s = 13;
	{8'd222,8'd179} : s = 60;
	{8'd222,8'd180} : s = 58;
	{8'd222,8'd181} : s = 179;
	{8'd222,8'd182} : s = 57;
	{8'd222,8'd183} : s = 174;
	{8'd222,8'd184} : s = 173;
	{8'd222,8'd185} : s = 318;
	{8'd222,8'd186} : s = 54;
	{8'd222,8'd187} : s = 171;
	{8'd222,8'd188} : s = 167;
	{8'd222,8'd189} : s = 317;
	{8'd222,8'd190} : s = 158;
	{8'd222,8'd191} : s = 315;
	{8'd222,8'd192} : s = 311;
	{8'd222,8'd193} : s = 446;
	{8'd222,8'd194} : s = 11;
	{8'd222,8'd195} : s = 53;
	{8'd222,8'd196} : s = 51;
	{8'd222,8'd197} : s = 157;
	{8'd222,8'd198} : s = 46;
	{8'd222,8'd199} : s = 155;
	{8'd222,8'd200} : s = 151;
	{8'd222,8'd201} : s = 303;
	{8'd222,8'd202} : s = 45;
	{8'd222,8'd203} : s = 143;
	{8'd222,8'd204} : s = 124;
	{8'd222,8'd205} : s = 287;
	{8'd222,8'd206} : s = 122;
	{8'd222,8'd207} : s = 252;
	{8'd222,8'd208} : s = 250;
	{8'd222,8'd209} : s = 445;
	{8'd222,8'd210} : s = 43;
	{8'd222,8'd211} : s = 121;
	{8'd222,8'd212} : s = 118;
	{8'd222,8'd213} : s = 249;
	{8'd222,8'd214} : s = 117;
	{8'd222,8'd215} : s = 246;
	{8'd222,8'd216} : s = 245;
	{8'd222,8'd217} : s = 443;
	{8'd222,8'd218} : s = 115;
	{8'd222,8'd219} : s = 243;
	{8'd222,8'd220} : s = 238;
	{8'd222,8'd221} : s = 439;
	{8'd222,8'd222} : s = 237;
	{8'd222,8'd223} : s = 431;
	{8'd222,8'd224} : s = 415;
	{8'd222,8'd225} : s = 507;
	{8'd222,8'd226} : s = 7;
	{8'd222,8'd227} : s = 39;
	{8'd222,8'd228} : s = 30;
	{8'd222,8'd229} : s = 110;
	{8'd222,8'd230} : s = 29;
	{8'd222,8'd231} : s = 109;
	{8'd222,8'd232} : s = 107;
	{8'd222,8'd233} : s = 235;
	{8'd222,8'd234} : s = 27;
	{8'd222,8'd235} : s = 103;
	{8'd222,8'd236} : s = 94;
	{8'd222,8'd237} : s = 231;
	{8'd222,8'd238} : s = 93;
	{8'd222,8'd239} : s = 222;
	{8'd222,8'd240} : s = 221;
	{8'd222,8'd241} : s = 382;
	{8'd222,8'd242} : s = 23;
	{8'd222,8'd243} : s = 91;
	{8'd222,8'd244} : s = 87;
	{8'd222,8'd245} : s = 219;
	{8'd222,8'd246} : s = 79;
	{8'd222,8'd247} : s = 215;
	{8'd222,8'd248} : s = 207;
	{8'd222,8'd249} : s = 381;
	{8'd222,8'd250} : s = 62;
	{8'd222,8'd251} : s = 190;
	{8'd222,8'd252} : s = 189;
	{8'd222,8'd253} : s = 379;
	{8'd222,8'd254} : s = 187;
	{8'd222,8'd255} : s = 375;
	{8'd223,8'd0} : s = 505;
	{8'd223,8'd1} : s = 84;
	{8'd223,8'd2} : s = 204;
	{8'd223,8'd3} : s = 202;
	{8'd223,8'd4} : s = 346;
	{8'd223,8'd5} : s = 201;
	{8'd223,8'd6} : s = 345;
	{8'd223,8'd7} : s = 342;
	{8'd223,8'd8} : s = 459;
	{8'd223,8'd9} : s = 198;
	{8'd223,8'd10} : s = 341;
	{8'd223,8'd11} : s = 339;
	{8'd223,8'd12} : s = 455;
	{8'd223,8'd13} : s = 334;
	{8'd223,8'd14} : s = 444;
	{8'd223,8'd15} : s = 442;
	{8'd223,8'd16} : s = 502;
	{8'd223,8'd17} : s = 197;
	{8'd223,8'd18} : s = 333;
	{8'd223,8'd19} : s = 331;
	{8'd223,8'd20} : s = 441;
	{8'd223,8'd21} : s = 327;
	{8'd223,8'd22} : s = 438;
	{8'd223,8'd23} : s = 437;
	{8'd223,8'd24} : s = 501;
	{8'd223,8'd25} : s = 316;
	{8'd223,8'd26} : s = 435;
	{8'd223,8'd27} : s = 430;
	{8'd223,8'd28} : s = 499;
	{8'd223,8'd29} : s = 429;
	{8'd223,8'd30} : s = 494;
	{8'd223,8'd31} : s = 493;
	{8'd223,8'd32} : s = 510;
	{8'd223,8'd33} : s = 1;
	{8'd223,8'd34} : s = 18;
	{8'd223,8'd35} : s = 17;
	{8'd223,8'd36} : s = 82;
	{8'd223,8'd37} : s = 12;
	{8'd223,8'd38} : s = 81;
	{8'd223,8'd39} : s = 76;
	{8'd223,8'd40} : s = 195;
	{8'd223,8'd41} : s = 10;
	{8'd223,8'd42} : s = 74;
	{8'd223,8'd43} : s = 73;
	{8'd223,8'd44} : s = 184;
	{8'd223,8'd45} : s = 70;
	{8'd223,8'd46} : s = 180;
	{8'd223,8'd47} : s = 178;
	{8'd223,8'd48} : s = 314;
	{8'd223,8'd49} : s = 9;
	{8'd223,8'd50} : s = 69;
	{8'd223,8'd51} : s = 67;
	{8'd223,8'd52} : s = 177;
	{8'd223,8'd53} : s = 56;
	{8'd223,8'd54} : s = 172;
	{8'd223,8'd55} : s = 170;
	{8'd223,8'd56} : s = 313;
	{8'd223,8'd57} : s = 52;
	{8'd223,8'd58} : s = 169;
	{8'd223,8'd59} : s = 166;
	{8'd223,8'd60} : s = 310;
	{8'd223,8'd61} : s = 165;
	{8'd223,8'd62} : s = 309;
	{8'd223,8'd63} : s = 307;
	{8'd223,8'd64} : s = 427;
	{8'd223,8'd65} : s = 6;
	{8'd223,8'd66} : s = 50;
	{8'd223,8'd67} : s = 49;
	{8'd223,8'd68} : s = 163;
	{8'd223,8'd69} : s = 44;
	{8'd223,8'd70} : s = 156;
	{8'd223,8'd71} : s = 154;
	{8'd223,8'd72} : s = 302;
	{8'd223,8'd73} : s = 42;
	{8'd223,8'd74} : s = 153;
	{8'd223,8'd75} : s = 150;
	{8'd223,8'd76} : s = 301;
	{8'd223,8'd77} : s = 149;
	{8'd223,8'd78} : s = 299;
	{8'd223,8'd79} : s = 295;
	{8'd223,8'd80} : s = 423;
	{8'd223,8'd81} : s = 41;
	{8'd223,8'd82} : s = 147;
	{8'd223,8'd83} : s = 142;
	{8'd223,8'd84} : s = 286;
	{8'd223,8'd85} : s = 141;
	{8'd223,8'd86} : s = 285;
	{8'd223,8'd87} : s = 283;
	{8'd223,8'd88} : s = 414;
	{8'd223,8'd89} : s = 139;
	{8'd223,8'd90} : s = 279;
	{8'd223,8'd91} : s = 271;
	{8'd223,8'd92} : s = 413;
	{8'd223,8'd93} : s = 248;
	{8'd223,8'd94} : s = 411;
	{8'd223,8'd95} : s = 407;
	{8'd223,8'd96} : s = 491;
	{8'd223,8'd97} : s = 5;
	{8'd223,8'd98} : s = 38;
	{8'd223,8'd99} : s = 37;
	{8'd223,8'd100} : s = 135;
	{8'd223,8'd101} : s = 35;
	{8'd223,8'd102} : s = 120;
	{8'd223,8'd103} : s = 116;
	{8'd223,8'd104} : s = 244;
	{8'd223,8'd105} : s = 28;
	{8'd223,8'd106} : s = 114;
	{8'd223,8'd107} : s = 113;
	{8'd223,8'd108} : s = 242;
	{8'd223,8'd109} : s = 108;
	{8'd223,8'd110} : s = 241;
	{8'd223,8'd111} : s = 236;
	{8'd223,8'd112} : s = 399;
	{8'd223,8'd113} : s = 26;
	{8'd223,8'd114} : s = 106;
	{8'd223,8'd115} : s = 105;
	{8'd223,8'd116} : s = 234;
	{8'd223,8'd117} : s = 102;
	{8'd223,8'd118} : s = 233;
	{8'd223,8'd119} : s = 230;
	{8'd223,8'd120} : s = 380;
	{8'd223,8'd121} : s = 101;
	{8'd223,8'd122} : s = 229;
	{8'd223,8'd123} : s = 227;
	{8'd223,8'd124} : s = 378;
	{8'd223,8'd125} : s = 220;
	{8'd223,8'd126} : s = 377;
	{8'd223,8'd127} : s = 374;
	{8'd223,8'd128} : s = 487;
	{8'd223,8'd129} : s = 25;
	{8'd223,8'd130} : s = 99;
	{8'd223,8'd131} : s = 92;
	{8'd223,8'd132} : s = 218;
	{8'd223,8'd133} : s = 90;
	{8'd223,8'd134} : s = 217;
	{8'd223,8'd135} : s = 214;
	{8'd223,8'd136} : s = 373;
	{8'd223,8'd137} : s = 89;
	{8'd223,8'd138} : s = 213;
	{8'd223,8'd139} : s = 211;
	{8'd223,8'd140} : s = 371;
	{8'd223,8'd141} : s = 206;
	{8'd223,8'd142} : s = 366;
	{8'd223,8'd143} : s = 365;
	{8'd223,8'd144} : s = 478;
	{8'd223,8'd145} : s = 86;
	{8'd223,8'd146} : s = 205;
	{8'd223,8'd147} : s = 203;
	{8'd223,8'd148} : s = 363;
	{8'd223,8'd149} : s = 199;
	{8'd223,8'd150} : s = 359;
	{8'd223,8'd151} : s = 350;
	{8'd223,8'd152} : s = 477;
	{8'd223,8'd153} : s = 188;
	{8'd223,8'd154} : s = 349;
	{8'd223,8'd155} : s = 347;
	{8'd223,8'd156} : s = 475;
	{8'd223,8'd157} : s = 343;
	{8'd223,8'd158} : s = 471;
	{8'd223,8'd159} : s = 463;
	{8'd223,8'd160} : s = 509;
	{8'd223,8'd161} : s = 3;
	{8'd223,8'd162} : s = 22;
	{8'd223,8'd163} : s = 21;
	{8'd223,8'd164} : s = 85;
	{8'd223,8'd165} : s = 19;
	{8'd223,8'd166} : s = 83;
	{8'd223,8'd167} : s = 78;
	{8'd223,8'd168} : s = 186;
	{8'd223,8'd169} : s = 14;
	{8'd223,8'd170} : s = 77;
	{8'd223,8'd171} : s = 75;
	{8'd223,8'd172} : s = 185;
	{8'd223,8'd173} : s = 71;
	{8'd223,8'd174} : s = 182;
	{8'd223,8'd175} : s = 181;
	{8'd223,8'd176} : s = 335;
	{8'd223,8'd177} : s = 13;
	{8'd223,8'd178} : s = 60;
	{8'd223,8'd179} : s = 58;
	{8'd223,8'd180} : s = 179;
	{8'd223,8'd181} : s = 57;
	{8'd223,8'd182} : s = 174;
	{8'd223,8'd183} : s = 173;
	{8'd223,8'd184} : s = 318;
	{8'd223,8'd185} : s = 54;
	{8'd223,8'd186} : s = 171;
	{8'd223,8'd187} : s = 167;
	{8'd223,8'd188} : s = 317;
	{8'd223,8'd189} : s = 158;
	{8'd223,8'd190} : s = 315;
	{8'd223,8'd191} : s = 311;
	{8'd223,8'd192} : s = 446;
	{8'd223,8'd193} : s = 11;
	{8'd223,8'd194} : s = 53;
	{8'd223,8'd195} : s = 51;
	{8'd223,8'd196} : s = 157;
	{8'd223,8'd197} : s = 46;
	{8'd223,8'd198} : s = 155;
	{8'd223,8'd199} : s = 151;
	{8'd223,8'd200} : s = 303;
	{8'd223,8'd201} : s = 45;
	{8'd223,8'd202} : s = 143;
	{8'd223,8'd203} : s = 124;
	{8'd223,8'd204} : s = 287;
	{8'd223,8'd205} : s = 122;
	{8'd223,8'd206} : s = 252;
	{8'd223,8'd207} : s = 250;
	{8'd223,8'd208} : s = 445;
	{8'd223,8'd209} : s = 43;
	{8'd223,8'd210} : s = 121;
	{8'd223,8'd211} : s = 118;
	{8'd223,8'd212} : s = 249;
	{8'd223,8'd213} : s = 117;
	{8'd223,8'd214} : s = 246;
	{8'd223,8'd215} : s = 245;
	{8'd223,8'd216} : s = 443;
	{8'd223,8'd217} : s = 115;
	{8'd223,8'd218} : s = 243;
	{8'd223,8'd219} : s = 238;
	{8'd223,8'd220} : s = 439;
	{8'd223,8'd221} : s = 237;
	{8'd223,8'd222} : s = 431;
	{8'd223,8'd223} : s = 415;
	{8'd223,8'd224} : s = 507;
	{8'd223,8'd225} : s = 7;
	{8'd223,8'd226} : s = 39;
	{8'd223,8'd227} : s = 30;
	{8'd223,8'd228} : s = 110;
	{8'd223,8'd229} : s = 29;
	{8'd223,8'd230} : s = 109;
	{8'd223,8'd231} : s = 107;
	{8'd223,8'd232} : s = 235;
	{8'd223,8'd233} : s = 27;
	{8'd223,8'd234} : s = 103;
	{8'd223,8'd235} : s = 94;
	{8'd223,8'd236} : s = 231;
	{8'd223,8'd237} : s = 93;
	{8'd223,8'd238} : s = 222;
	{8'd223,8'd239} : s = 221;
	{8'd223,8'd240} : s = 382;
	{8'd223,8'd241} : s = 23;
	{8'd223,8'd242} : s = 91;
	{8'd223,8'd243} : s = 87;
	{8'd223,8'd244} : s = 219;
	{8'd223,8'd245} : s = 79;
	{8'd223,8'd246} : s = 215;
	{8'd223,8'd247} : s = 207;
	{8'd223,8'd248} : s = 381;
	{8'd223,8'd249} : s = 62;
	{8'd223,8'd250} : s = 190;
	{8'd223,8'd251} : s = 189;
	{8'd223,8'd252} : s = 379;
	{8'd223,8'd253} : s = 187;
	{8'd223,8'd254} : s = 375;
	{8'd223,8'd255} : s = 367;
	{8'd224,8'd0} : s = 84;
	{8'd224,8'd1} : s = 204;
	{8'd224,8'd2} : s = 202;
	{8'd224,8'd3} : s = 346;
	{8'd224,8'd4} : s = 201;
	{8'd224,8'd5} : s = 345;
	{8'd224,8'd6} : s = 342;
	{8'd224,8'd7} : s = 459;
	{8'd224,8'd8} : s = 198;
	{8'd224,8'd9} : s = 341;
	{8'd224,8'd10} : s = 339;
	{8'd224,8'd11} : s = 455;
	{8'd224,8'd12} : s = 334;
	{8'd224,8'd13} : s = 444;
	{8'd224,8'd14} : s = 442;
	{8'd224,8'd15} : s = 502;
	{8'd224,8'd16} : s = 197;
	{8'd224,8'd17} : s = 333;
	{8'd224,8'd18} : s = 331;
	{8'd224,8'd19} : s = 441;
	{8'd224,8'd20} : s = 327;
	{8'd224,8'd21} : s = 438;
	{8'd224,8'd22} : s = 437;
	{8'd224,8'd23} : s = 501;
	{8'd224,8'd24} : s = 316;
	{8'd224,8'd25} : s = 435;
	{8'd224,8'd26} : s = 430;
	{8'd224,8'd27} : s = 499;
	{8'd224,8'd28} : s = 429;
	{8'd224,8'd29} : s = 494;
	{8'd224,8'd30} : s = 493;
	{8'd224,8'd31} : s = 510;
	{8'd224,8'd32} : s = 1;
	{8'd224,8'd33} : s = 18;
	{8'd224,8'd34} : s = 17;
	{8'd224,8'd35} : s = 82;
	{8'd224,8'd36} : s = 12;
	{8'd224,8'd37} : s = 81;
	{8'd224,8'd38} : s = 76;
	{8'd224,8'd39} : s = 195;
	{8'd224,8'd40} : s = 10;
	{8'd224,8'd41} : s = 74;
	{8'd224,8'd42} : s = 73;
	{8'd224,8'd43} : s = 184;
	{8'd224,8'd44} : s = 70;
	{8'd224,8'd45} : s = 180;
	{8'd224,8'd46} : s = 178;
	{8'd224,8'd47} : s = 314;
	{8'd224,8'd48} : s = 9;
	{8'd224,8'd49} : s = 69;
	{8'd224,8'd50} : s = 67;
	{8'd224,8'd51} : s = 177;
	{8'd224,8'd52} : s = 56;
	{8'd224,8'd53} : s = 172;
	{8'd224,8'd54} : s = 170;
	{8'd224,8'd55} : s = 313;
	{8'd224,8'd56} : s = 52;
	{8'd224,8'd57} : s = 169;
	{8'd224,8'd58} : s = 166;
	{8'd224,8'd59} : s = 310;
	{8'd224,8'd60} : s = 165;
	{8'd224,8'd61} : s = 309;
	{8'd224,8'd62} : s = 307;
	{8'd224,8'd63} : s = 427;
	{8'd224,8'd64} : s = 6;
	{8'd224,8'd65} : s = 50;
	{8'd224,8'd66} : s = 49;
	{8'd224,8'd67} : s = 163;
	{8'd224,8'd68} : s = 44;
	{8'd224,8'd69} : s = 156;
	{8'd224,8'd70} : s = 154;
	{8'd224,8'd71} : s = 302;
	{8'd224,8'd72} : s = 42;
	{8'd224,8'd73} : s = 153;
	{8'd224,8'd74} : s = 150;
	{8'd224,8'd75} : s = 301;
	{8'd224,8'd76} : s = 149;
	{8'd224,8'd77} : s = 299;
	{8'd224,8'd78} : s = 295;
	{8'd224,8'd79} : s = 423;
	{8'd224,8'd80} : s = 41;
	{8'd224,8'd81} : s = 147;
	{8'd224,8'd82} : s = 142;
	{8'd224,8'd83} : s = 286;
	{8'd224,8'd84} : s = 141;
	{8'd224,8'd85} : s = 285;
	{8'd224,8'd86} : s = 283;
	{8'd224,8'd87} : s = 414;
	{8'd224,8'd88} : s = 139;
	{8'd224,8'd89} : s = 279;
	{8'd224,8'd90} : s = 271;
	{8'd224,8'd91} : s = 413;
	{8'd224,8'd92} : s = 248;
	{8'd224,8'd93} : s = 411;
	{8'd224,8'd94} : s = 407;
	{8'd224,8'd95} : s = 491;
	{8'd224,8'd96} : s = 5;
	{8'd224,8'd97} : s = 38;
	{8'd224,8'd98} : s = 37;
	{8'd224,8'd99} : s = 135;
	{8'd224,8'd100} : s = 35;
	{8'd224,8'd101} : s = 120;
	{8'd224,8'd102} : s = 116;
	{8'd224,8'd103} : s = 244;
	{8'd224,8'd104} : s = 28;
	{8'd224,8'd105} : s = 114;
	{8'd224,8'd106} : s = 113;
	{8'd224,8'd107} : s = 242;
	{8'd224,8'd108} : s = 108;
	{8'd224,8'd109} : s = 241;
	{8'd224,8'd110} : s = 236;
	{8'd224,8'd111} : s = 399;
	{8'd224,8'd112} : s = 26;
	{8'd224,8'd113} : s = 106;
	{8'd224,8'd114} : s = 105;
	{8'd224,8'd115} : s = 234;
	{8'd224,8'd116} : s = 102;
	{8'd224,8'd117} : s = 233;
	{8'd224,8'd118} : s = 230;
	{8'd224,8'd119} : s = 380;
	{8'd224,8'd120} : s = 101;
	{8'd224,8'd121} : s = 229;
	{8'd224,8'd122} : s = 227;
	{8'd224,8'd123} : s = 378;
	{8'd224,8'd124} : s = 220;
	{8'd224,8'd125} : s = 377;
	{8'd224,8'd126} : s = 374;
	{8'd224,8'd127} : s = 487;
	{8'd224,8'd128} : s = 25;
	{8'd224,8'd129} : s = 99;
	{8'd224,8'd130} : s = 92;
	{8'd224,8'd131} : s = 218;
	{8'd224,8'd132} : s = 90;
	{8'd224,8'd133} : s = 217;
	{8'd224,8'd134} : s = 214;
	{8'd224,8'd135} : s = 373;
	{8'd224,8'd136} : s = 89;
	{8'd224,8'd137} : s = 213;
	{8'd224,8'd138} : s = 211;
	{8'd224,8'd139} : s = 371;
	{8'd224,8'd140} : s = 206;
	{8'd224,8'd141} : s = 366;
	{8'd224,8'd142} : s = 365;
	{8'd224,8'd143} : s = 478;
	{8'd224,8'd144} : s = 86;
	{8'd224,8'd145} : s = 205;
	{8'd224,8'd146} : s = 203;
	{8'd224,8'd147} : s = 363;
	{8'd224,8'd148} : s = 199;
	{8'd224,8'd149} : s = 359;
	{8'd224,8'd150} : s = 350;
	{8'd224,8'd151} : s = 477;
	{8'd224,8'd152} : s = 188;
	{8'd224,8'd153} : s = 349;
	{8'd224,8'd154} : s = 347;
	{8'd224,8'd155} : s = 475;
	{8'd224,8'd156} : s = 343;
	{8'd224,8'd157} : s = 471;
	{8'd224,8'd158} : s = 463;
	{8'd224,8'd159} : s = 509;
	{8'd224,8'd160} : s = 3;
	{8'd224,8'd161} : s = 22;
	{8'd224,8'd162} : s = 21;
	{8'd224,8'd163} : s = 85;
	{8'd224,8'd164} : s = 19;
	{8'd224,8'd165} : s = 83;
	{8'd224,8'd166} : s = 78;
	{8'd224,8'd167} : s = 186;
	{8'd224,8'd168} : s = 14;
	{8'd224,8'd169} : s = 77;
	{8'd224,8'd170} : s = 75;
	{8'd224,8'd171} : s = 185;
	{8'd224,8'd172} : s = 71;
	{8'd224,8'd173} : s = 182;
	{8'd224,8'd174} : s = 181;
	{8'd224,8'd175} : s = 335;
	{8'd224,8'd176} : s = 13;
	{8'd224,8'd177} : s = 60;
	{8'd224,8'd178} : s = 58;
	{8'd224,8'd179} : s = 179;
	{8'd224,8'd180} : s = 57;
	{8'd224,8'd181} : s = 174;
	{8'd224,8'd182} : s = 173;
	{8'd224,8'd183} : s = 318;
	{8'd224,8'd184} : s = 54;
	{8'd224,8'd185} : s = 171;
	{8'd224,8'd186} : s = 167;
	{8'd224,8'd187} : s = 317;
	{8'd224,8'd188} : s = 158;
	{8'd224,8'd189} : s = 315;
	{8'd224,8'd190} : s = 311;
	{8'd224,8'd191} : s = 446;
	{8'd224,8'd192} : s = 11;
	{8'd224,8'd193} : s = 53;
	{8'd224,8'd194} : s = 51;
	{8'd224,8'd195} : s = 157;
	{8'd224,8'd196} : s = 46;
	{8'd224,8'd197} : s = 155;
	{8'd224,8'd198} : s = 151;
	{8'd224,8'd199} : s = 303;
	{8'd224,8'd200} : s = 45;
	{8'd224,8'd201} : s = 143;
	{8'd224,8'd202} : s = 124;
	{8'd224,8'd203} : s = 287;
	{8'd224,8'd204} : s = 122;
	{8'd224,8'd205} : s = 252;
	{8'd224,8'd206} : s = 250;
	{8'd224,8'd207} : s = 445;
	{8'd224,8'd208} : s = 43;
	{8'd224,8'd209} : s = 121;
	{8'd224,8'd210} : s = 118;
	{8'd224,8'd211} : s = 249;
	{8'd224,8'd212} : s = 117;
	{8'd224,8'd213} : s = 246;
	{8'd224,8'd214} : s = 245;
	{8'd224,8'd215} : s = 443;
	{8'd224,8'd216} : s = 115;
	{8'd224,8'd217} : s = 243;
	{8'd224,8'd218} : s = 238;
	{8'd224,8'd219} : s = 439;
	{8'd224,8'd220} : s = 237;
	{8'd224,8'd221} : s = 431;
	{8'd224,8'd222} : s = 415;
	{8'd224,8'd223} : s = 507;
	{8'd224,8'd224} : s = 7;
	{8'd224,8'd225} : s = 39;
	{8'd224,8'd226} : s = 30;
	{8'd224,8'd227} : s = 110;
	{8'd224,8'd228} : s = 29;
	{8'd224,8'd229} : s = 109;
	{8'd224,8'd230} : s = 107;
	{8'd224,8'd231} : s = 235;
	{8'd224,8'd232} : s = 27;
	{8'd224,8'd233} : s = 103;
	{8'd224,8'd234} : s = 94;
	{8'd224,8'd235} : s = 231;
	{8'd224,8'd236} : s = 93;
	{8'd224,8'd237} : s = 222;
	{8'd224,8'd238} : s = 221;
	{8'd224,8'd239} : s = 382;
	{8'd224,8'd240} : s = 23;
	{8'd224,8'd241} : s = 91;
	{8'd224,8'd242} : s = 87;
	{8'd224,8'd243} : s = 219;
	{8'd224,8'd244} : s = 79;
	{8'd224,8'd245} : s = 215;
	{8'd224,8'd246} : s = 207;
	{8'd224,8'd247} : s = 381;
	{8'd224,8'd248} : s = 62;
	{8'd224,8'd249} : s = 190;
	{8'd224,8'd250} : s = 189;
	{8'd224,8'd251} : s = 379;
	{8'd224,8'd252} : s = 187;
	{8'd224,8'd253} : s = 375;
	{8'd224,8'd254} : s = 367;
	{8'd224,8'd255} : s = 503;
	{8'd225,8'd0} : s = 204;
	{8'd225,8'd1} : s = 202;
	{8'd225,8'd2} : s = 346;
	{8'd225,8'd3} : s = 201;
	{8'd225,8'd4} : s = 345;
	{8'd225,8'd5} : s = 342;
	{8'd225,8'd6} : s = 459;
	{8'd225,8'd7} : s = 198;
	{8'd225,8'd8} : s = 341;
	{8'd225,8'd9} : s = 339;
	{8'd225,8'd10} : s = 455;
	{8'd225,8'd11} : s = 334;
	{8'd225,8'd12} : s = 444;
	{8'd225,8'd13} : s = 442;
	{8'd225,8'd14} : s = 502;
	{8'd225,8'd15} : s = 197;
	{8'd225,8'd16} : s = 333;
	{8'd225,8'd17} : s = 331;
	{8'd225,8'd18} : s = 441;
	{8'd225,8'd19} : s = 327;
	{8'd225,8'd20} : s = 438;
	{8'd225,8'd21} : s = 437;
	{8'd225,8'd22} : s = 501;
	{8'd225,8'd23} : s = 316;
	{8'd225,8'd24} : s = 435;
	{8'd225,8'd25} : s = 430;
	{8'd225,8'd26} : s = 499;
	{8'd225,8'd27} : s = 429;
	{8'd225,8'd28} : s = 494;
	{8'd225,8'd29} : s = 493;
	{8'd225,8'd30} : s = 510;
	{8'd225,8'd31} : s = 1;
	{8'd225,8'd32} : s = 18;
	{8'd225,8'd33} : s = 17;
	{8'd225,8'd34} : s = 82;
	{8'd225,8'd35} : s = 12;
	{8'd225,8'd36} : s = 81;
	{8'd225,8'd37} : s = 76;
	{8'd225,8'd38} : s = 195;
	{8'd225,8'd39} : s = 10;
	{8'd225,8'd40} : s = 74;
	{8'd225,8'd41} : s = 73;
	{8'd225,8'd42} : s = 184;
	{8'd225,8'd43} : s = 70;
	{8'd225,8'd44} : s = 180;
	{8'd225,8'd45} : s = 178;
	{8'd225,8'd46} : s = 314;
	{8'd225,8'd47} : s = 9;
	{8'd225,8'd48} : s = 69;
	{8'd225,8'd49} : s = 67;
	{8'd225,8'd50} : s = 177;
	{8'd225,8'd51} : s = 56;
	{8'd225,8'd52} : s = 172;
	{8'd225,8'd53} : s = 170;
	{8'd225,8'd54} : s = 313;
	{8'd225,8'd55} : s = 52;
	{8'd225,8'd56} : s = 169;
	{8'd225,8'd57} : s = 166;
	{8'd225,8'd58} : s = 310;
	{8'd225,8'd59} : s = 165;
	{8'd225,8'd60} : s = 309;
	{8'd225,8'd61} : s = 307;
	{8'd225,8'd62} : s = 427;
	{8'd225,8'd63} : s = 6;
	{8'd225,8'd64} : s = 50;
	{8'd225,8'd65} : s = 49;
	{8'd225,8'd66} : s = 163;
	{8'd225,8'd67} : s = 44;
	{8'd225,8'd68} : s = 156;
	{8'd225,8'd69} : s = 154;
	{8'd225,8'd70} : s = 302;
	{8'd225,8'd71} : s = 42;
	{8'd225,8'd72} : s = 153;
	{8'd225,8'd73} : s = 150;
	{8'd225,8'd74} : s = 301;
	{8'd225,8'd75} : s = 149;
	{8'd225,8'd76} : s = 299;
	{8'd225,8'd77} : s = 295;
	{8'd225,8'd78} : s = 423;
	{8'd225,8'd79} : s = 41;
	{8'd225,8'd80} : s = 147;
	{8'd225,8'd81} : s = 142;
	{8'd225,8'd82} : s = 286;
	{8'd225,8'd83} : s = 141;
	{8'd225,8'd84} : s = 285;
	{8'd225,8'd85} : s = 283;
	{8'd225,8'd86} : s = 414;
	{8'd225,8'd87} : s = 139;
	{8'd225,8'd88} : s = 279;
	{8'd225,8'd89} : s = 271;
	{8'd225,8'd90} : s = 413;
	{8'd225,8'd91} : s = 248;
	{8'd225,8'd92} : s = 411;
	{8'd225,8'd93} : s = 407;
	{8'd225,8'd94} : s = 491;
	{8'd225,8'd95} : s = 5;
	{8'd225,8'd96} : s = 38;
	{8'd225,8'd97} : s = 37;
	{8'd225,8'd98} : s = 135;
	{8'd225,8'd99} : s = 35;
	{8'd225,8'd100} : s = 120;
	{8'd225,8'd101} : s = 116;
	{8'd225,8'd102} : s = 244;
	{8'd225,8'd103} : s = 28;
	{8'd225,8'd104} : s = 114;
	{8'd225,8'd105} : s = 113;
	{8'd225,8'd106} : s = 242;
	{8'd225,8'd107} : s = 108;
	{8'd225,8'd108} : s = 241;
	{8'd225,8'd109} : s = 236;
	{8'd225,8'd110} : s = 399;
	{8'd225,8'd111} : s = 26;
	{8'd225,8'd112} : s = 106;
	{8'd225,8'd113} : s = 105;
	{8'd225,8'd114} : s = 234;
	{8'd225,8'd115} : s = 102;
	{8'd225,8'd116} : s = 233;
	{8'd225,8'd117} : s = 230;
	{8'd225,8'd118} : s = 380;
	{8'd225,8'd119} : s = 101;
	{8'd225,8'd120} : s = 229;
	{8'd225,8'd121} : s = 227;
	{8'd225,8'd122} : s = 378;
	{8'd225,8'd123} : s = 220;
	{8'd225,8'd124} : s = 377;
	{8'd225,8'd125} : s = 374;
	{8'd225,8'd126} : s = 487;
	{8'd225,8'd127} : s = 25;
	{8'd225,8'd128} : s = 99;
	{8'd225,8'd129} : s = 92;
	{8'd225,8'd130} : s = 218;
	{8'd225,8'd131} : s = 90;
	{8'd225,8'd132} : s = 217;
	{8'd225,8'd133} : s = 214;
	{8'd225,8'd134} : s = 373;
	{8'd225,8'd135} : s = 89;
	{8'd225,8'd136} : s = 213;
	{8'd225,8'd137} : s = 211;
	{8'd225,8'd138} : s = 371;
	{8'd225,8'd139} : s = 206;
	{8'd225,8'd140} : s = 366;
	{8'd225,8'd141} : s = 365;
	{8'd225,8'd142} : s = 478;
	{8'd225,8'd143} : s = 86;
	{8'd225,8'd144} : s = 205;
	{8'd225,8'd145} : s = 203;
	{8'd225,8'd146} : s = 363;
	{8'd225,8'd147} : s = 199;
	{8'd225,8'd148} : s = 359;
	{8'd225,8'd149} : s = 350;
	{8'd225,8'd150} : s = 477;
	{8'd225,8'd151} : s = 188;
	{8'd225,8'd152} : s = 349;
	{8'd225,8'd153} : s = 347;
	{8'd225,8'd154} : s = 475;
	{8'd225,8'd155} : s = 343;
	{8'd225,8'd156} : s = 471;
	{8'd225,8'd157} : s = 463;
	{8'd225,8'd158} : s = 509;
	{8'd225,8'd159} : s = 3;
	{8'd225,8'd160} : s = 22;
	{8'd225,8'd161} : s = 21;
	{8'd225,8'd162} : s = 85;
	{8'd225,8'd163} : s = 19;
	{8'd225,8'd164} : s = 83;
	{8'd225,8'd165} : s = 78;
	{8'd225,8'd166} : s = 186;
	{8'd225,8'd167} : s = 14;
	{8'd225,8'd168} : s = 77;
	{8'd225,8'd169} : s = 75;
	{8'd225,8'd170} : s = 185;
	{8'd225,8'd171} : s = 71;
	{8'd225,8'd172} : s = 182;
	{8'd225,8'd173} : s = 181;
	{8'd225,8'd174} : s = 335;
	{8'd225,8'd175} : s = 13;
	{8'd225,8'd176} : s = 60;
	{8'd225,8'd177} : s = 58;
	{8'd225,8'd178} : s = 179;
	{8'd225,8'd179} : s = 57;
	{8'd225,8'd180} : s = 174;
	{8'd225,8'd181} : s = 173;
	{8'd225,8'd182} : s = 318;
	{8'd225,8'd183} : s = 54;
	{8'd225,8'd184} : s = 171;
	{8'd225,8'd185} : s = 167;
	{8'd225,8'd186} : s = 317;
	{8'd225,8'd187} : s = 158;
	{8'd225,8'd188} : s = 315;
	{8'd225,8'd189} : s = 311;
	{8'd225,8'd190} : s = 446;
	{8'd225,8'd191} : s = 11;
	{8'd225,8'd192} : s = 53;
	{8'd225,8'd193} : s = 51;
	{8'd225,8'd194} : s = 157;
	{8'd225,8'd195} : s = 46;
	{8'd225,8'd196} : s = 155;
	{8'd225,8'd197} : s = 151;
	{8'd225,8'd198} : s = 303;
	{8'd225,8'd199} : s = 45;
	{8'd225,8'd200} : s = 143;
	{8'd225,8'd201} : s = 124;
	{8'd225,8'd202} : s = 287;
	{8'd225,8'd203} : s = 122;
	{8'd225,8'd204} : s = 252;
	{8'd225,8'd205} : s = 250;
	{8'd225,8'd206} : s = 445;
	{8'd225,8'd207} : s = 43;
	{8'd225,8'd208} : s = 121;
	{8'd225,8'd209} : s = 118;
	{8'd225,8'd210} : s = 249;
	{8'd225,8'd211} : s = 117;
	{8'd225,8'd212} : s = 246;
	{8'd225,8'd213} : s = 245;
	{8'd225,8'd214} : s = 443;
	{8'd225,8'd215} : s = 115;
	{8'd225,8'd216} : s = 243;
	{8'd225,8'd217} : s = 238;
	{8'd225,8'd218} : s = 439;
	{8'd225,8'd219} : s = 237;
	{8'd225,8'd220} : s = 431;
	{8'd225,8'd221} : s = 415;
	{8'd225,8'd222} : s = 507;
	{8'd225,8'd223} : s = 7;
	{8'd225,8'd224} : s = 39;
	{8'd225,8'd225} : s = 30;
	{8'd225,8'd226} : s = 110;
	{8'd225,8'd227} : s = 29;
	{8'd225,8'd228} : s = 109;
	{8'd225,8'd229} : s = 107;
	{8'd225,8'd230} : s = 235;
	{8'd225,8'd231} : s = 27;
	{8'd225,8'd232} : s = 103;
	{8'd225,8'd233} : s = 94;
	{8'd225,8'd234} : s = 231;
	{8'd225,8'd235} : s = 93;
	{8'd225,8'd236} : s = 222;
	{8'd225,8'd237} : s = 221;
	{8'd225,8'd238} : s = 382;
	{8'd225,8'd239} : s = 23;
	{8'd225,8'd240} : s = 91;
	{8'd225,8'd241} : s = 87;
	{8'd225,8'd242} : s = 219;
	{8'd225,8'd243} : s = 79;
	{8'd225,8'd244} : s = 215;
	{8'd225,8'd245} : s = 207;
	{8'd225,8'd246} : s = 381;
	{8'd225,8'd247} : s = 62;
	{8'd225,8'd248} : s = 190;
	{8'd225,8'd249} : s = 189;
	{8'd225,8'd250} : s = 379;
	{8'd225,8'd251} : s = 187;
	{8'd225,8'd252} : s = 375;
	{8'd225,8'd253} : s = 367;
	{8'd225,8'd254} : s = 503;
	{8'd225,8'd255} : s = 15;
	{8'd226,8'd0} : s = 202;
	{8'd226,8'd1} : s = 346;
	{8'd226,8'd2} : s = 201;
	{8'd226,8'd3} : s = 345;
	{8'd226,8'd4} : s = 342;
	{8'd226,8'd5} : s = 459;
	{8'd226,8'd6} : s = 198;
	{8'd226,8'd7} : s = 341;
	{8'd226,8'd8} : s = 339;
	{8'd226,8'd9} : s = 455;
	{8'd226,8'd10} : s = 334;
	{8'd226,8'd11} : s = 444;
	{8'd226,8'd12} : s = 442;
	{8'd226,8'd13} : s = 502;
	{8'd226,8'd14} : s = 197;
	{8'd226,8'd15} : s = 333;
	{8'd226,8'd16} : s = 331;
	{8'd226,8'd17} : s = 441;
	{8'd226,8'd18} : s = 327;
	{8'd226,8'd19} : s = 438;
	{8'd226,8'd20} : s = 437;
	{8'd226,8'd21} : s = 501;
	{8'd226,8'd22} : s = 316;
	{8'd226,8'd23} : s = 435;
	{8'd226,8'd24} : s = 430;
	{8'd226,8'd25} : s = 499;
	{8'd226,8'd26} : s = 429;
	{8'd226,8'd27} : s = 494;
	{8'd226,8'd28} : s = 493;
	{8'd226,8'd29} : s = 510;
	{8'd226,8'd30} : s = 1;
	{8'd226,8'd31} : s = 18;
	{8'd226,8'd32} : s = 17;
	{8'd226,8'd33} : s = 82;
	{8'd226,8'd34} : s = 12;
	{8'd226,8'd35} : s = 81;
	{8'd226,8'd36} : s = 76;
	{8'd226,8'd37} : s = 195;
	{8'd226,8'd38} : s = 10;
	{8'd226,8'd39} : s = 74;
	{8'd226,8'd40} : s = 73;
	{8'd226,8'd41} : s = 184;
	{8'd226,8'd42} : s = 70;
	{8'd226,8'd43} : s = 180;
	{8'd226,8'd44} : s = 178;
	{8'd226,8'd45} : s = 314;
	{8'd226,8'd46} : s = 9;
	{8'd226,8'd47} : s = 69;
	{8'd226,8'd48} : s = 67;
	{8'd226,8'd49} : s = 177;
	{8'd226,8'd50} : s = 56;
	{8'd226,8'd51} : s = 172;
	{8'd226,8'd52} : s = 170;
	{8'd226,8'd53} : s = 313;
	{8'd226,8'd54} : s = 52;
	{8'd226,8'd55} : s = 169;
	{8'd226,8'd56} : s = 166;
	{8'd226,8'd57} : s = 310;
	{8'd226,8'd58} : s = 165;
	{8'd226,8'd59} : s = 309;
	{8'd226,8'd60} : s = 307;
	{8'd226,8'd61} : s = 427;
	{8'd226,8'd62} : s = 6;
	{8'd226,8'd63} : s = 50;
	{8'd226,8'd64} : s = 49;
	{8'd226,8'd65} : s = 163;
	{8'd226,8'd66} : s = 44;
	{8'd226,8'd67} : s = 156;
	{8'd226,8'd68} : s = 154;
	{8'd226,8'd69} : s = 302;
	{8'd226,8'd70} : s = 42;
	{8'd226,8'd71} : s = 153;
	{8'd226,8'd72} : s = 150;
	{8'd226,8'd73} : s = 301;
	{8'd226,8'd74} : s = 149;
	{8'd226,8'd75} : s = 299;
	{8'd226,8'd76} : s = 295;
	{8'd226,8'd77} : s = 423;
	{8'd226,8'd78} : s = 41;
	{8'd226,8'd79} : s = 147;
	{8'd226,8'd80} : s = 142;
	{8'd226,8'd81} : s = 286;
	{8'd226,8'd82} : s = 141;
	{8'd226,8'd83} : s = 285;
	{8'd226,8'd84} : s = 283;
	{8'd226,8'd85} : s = 414;
	{8'd226,8'd86} : s = 139;
	{8'd226,8'd87} : s = 279;
	{8'd226,8'd88} : s = 271;
	{8'd226,8'd89} : s = 413;
	{8'd226,8'd90} : s = 248;
	{8'd226,8'd91} : s = 411;
	{8'd226,8'd92} : s = 407;
	{8'd226,8'd93} : s = 491;
	{8'd226,8'd94} : s = 5;
	{8'd226,8'd95} : s = 38;
	{8'd226,8'd96} : s = 37;
	{8'd226,8'd97} : s = 135;
	{8'd226,8'd98} : s = 35;
	{8'd226,8'd99} : s = 120;
	{8'd226,8'd100} : s = 116;
	{8'd226,8'd101} : s = 244;
	{8'd226,8'd102} : s = 28;
	{8'd226,8'd103} : s = 114;
	{8'd226,8'd104} : s = 113;
	{8'd226,8'd105} : s = 242;
	{8'd226,8'd106} : s = 108;
	{8'd226,8'd107} : s = 241;
	{8'd226,8'd108} : s = 236;
	{8'd226,8'd109} : s = 399;
	{8'd226,8'd110} : s = 26;
	{8'd226,8'd111} : s = 106;
	{8'd226,8'd112} : s = 105;
	{8'd226,8'd113} : s = 234;
	{8'd226,8'd114} : s = 102;
	{8'd226,8'd115} : s = 233;
	{8'd226,8'd116} : s = 230;
	{8'd226,8'd117} : s = 380;
	{8'd226,8'd118} : s = 101;
	{8'd226,8'd119} : s = 229;
	{8'd226,8'd120} : s = 227;
	{8'd226,8'd121} : s = 378;
	{8'd226,8'd122} : s = 220;
	{8'd226,8'd123} : s = 377;
	{8'd226,8'd124} : s = 374;
	{8'd226,8'd125} : s = 487;
	{8'd226,8'd126} : s = 25;
	{8'd226,8'd127} : s = 99;
	{8'd226,8'd128} : s = 92;
	{8'd226,8'd129} : s = 218;
	{8'd226,8'd130} : s = 90;
	{8'd226,8'd131} : s = 217;
	{8'd226,8'd132} : s = 214;
	{8'd226,8'd133} : s = 373;
	{8'd226,8'd134} : s = 89;
	{8'd226,8'd135} : s = 213;
	{8'd226,8'd136} : s = 211;
	{8'd226,8'd137} : s = 371;
	{8'd226,8'd138} : s = 206;
	{8'd226,8'd139} : s = 366;
	{8'd226,8'd140} : s = 365;
	{8'd226,8'd141} : s = 478;
	{8'd226,8'd142} : s = 86;
	{8'd226,8'd143} : s = 205;
	{8'd226,8'd144} : s = 203;
	{8'd226,8'd145} : s = 363;
	{8'd226,8'd146} : s = 199;
	{8'd226,8'd147} : s = 359;
	{8'd226,8'd148} : s = 350;
	{8'd226,8'd149} : s = 477;
	{8'd226,8'd150} : s = 188;
	{8'd226,8'd151} : s = 349;
	{8'd226,8'd152} : s = 347;
	{8'd226,8'd153} : s = 475;
	{8'd226,8'd154} : s = 343;
	{8'd226,8'd155} : s = 471;
	{8'd226,8'd156} : s = 463;
	{8'd226,8'd157} : s = 509;
	{8'd226,8'd158} : s = 3;
	{8'd226,8'd159} : s = 22;
	{8'd226,8'd160} : s = 21;
	{8'd226,8'd161} : s = 85;
	{8'd226,8'd162} : s = 19;
	{8'd226,8'd163} : s = 83;
	{8'd226,8'd164} : s = 78;
	{8'd226,8'd165} : s = 186;
	{8'd226,8'd166} : s = 14;
	{8'd226,8'd167} : s = 77;
	{8'd226,8'd168} : s = 75;
	{8'd226,8'd169} : s = 185;
	{8'd226,8'd170} : s = 71;
	{8'd226,8'd171} : s = 182;
	{8'd226,8'd172} : s = 181;
	{8'd226,8'd173} : s = 335;
	{8'd226,8'd174} : s = 13;
	{8'd226,8'd175} : s = 60;
	{8'd226,8'd176} : s = 58;
	{8'd226,8'd177} : s = 179;
	{8'd226,8'd178} : s = 57;
	{8'd226,8'd179} : s = 174;
	{8'd226,8'd180} : s = 173;
	{8'd226,8'd181} : s = 318;
	{8'd226,8'd182} : s = 54;
	{8'd226,8'd183} : s = 171;
	{8'd226,8'd184} : s = 167;
	{8'd226,8'd185} : s = 317;
	{8'd226,8'd186} : s = 158;
	{8'd226,8'd187} : s = 315;
	{8'd226,8'd188} : s = 311;
	{8'd226,8'd189} : s = 446;
	{8'd226,8'd190} : s = 11;
	{8'd226,8'd191} : s = 53;
	{8'd226,8'd192} : s = 51;
	{8'd226,8'd193} : s = 157;
	{8'd226,8'd194} : s = 46;
	{8'd226,8'd195} : s = 155;
	{8'd226,8'd196} : s = 151;
	{8'd226,8'd197} : s = 303;
	{8'd226,8'd198} : s = 45;
	{8'd226,8'd199} : s = 143;
	{8'd226,8'd200} : s = 124;
	{8'd226,8'd201} : s = 287;
	{8'd226,8'd202} : s = 122;
	{8'd226,8'd203} : s = 252;
	{8'd226,8'd204} : s = 250;
	{8'd226,8'd205} : s = 445;
	{8'd226,8'd206} : s = 43;
	{8'd226,8'd207} : s = 121;
	{8'd226,8'd208} : s = 118;
	{8'd226,8'd209} : s = 249;
	{8'd226,8'd210} : s = 117;
	{8'd226,8'd211} : s = 246;
	{8'd226,8'd212} : s = 245;
	{8'd226,8'd213} : s = 443;
	{8'd226,8'd214} : s = 115;
	{8'd226,8'd215} : s = 243;
	{8'd226,8'd216} : s = 238;
	{8'd226,8'd217} : s = 439;
	{8'd226,8'd218} : s = 237;
	{8'd226,8'd219} : s = 431;
	{8'd226,8'd220} : s = 415;
	{8'd226,8'd221} : s = 507;
	{8'd226,8'd222} : s = 7;
	{8'd226,8'd223} : s = 39;
	{8'd226,8'd224} : s = 30;
	{8'd226,8'd225} : s = 110;
	{8'd226,8'd226} : s = 29;
	{8'd226,8'd227} : s = 109;
	{8'd226,8'd228} : s = 107;
	{8'd226,8'd229} : s = 235;
	{8'd226,8'd230} : s = 27;
	{8'd226,8'd231} : s = 103;
	{8'd226,8'd232} : s = 94;
	{8'd226,8'd233} : s = 231;
	{8'd226,8'd234} : s = 93;
	{8'd226,8'd235} : s = 222;
	{8'd226,8'd236} : s = 221;
	{8'd226,8'd237} : s = 382;
	{8'd226,8'd238} : s = 23;
	{8'd226,8'd239} : s = 91;
	{8'd226,8'd240} : s = 87;
	{8'd226,8'd241} : s = 219;
	{8'd226,8'd242} : s = 79;
	{8'd226,8'd243} : s = 215;
	{8'd226,8'd244} : s = 207;
	{8'd226,8'd245} : s = 381;
	{8'd226,8'd246} : s = 62;
	{8'd226,8'd247} : s = 190;
	{8'd226,8'd248} : s = 189;
	{8'd226,8'd249} : s = 379;
	{8'd226,8'd250} : s = 187;
	{8'd226,8'd251} : s = 375;
	{8'd226,8'd252} : s = 367;
	{8'd226,8'd253} : s = 503;
	{8'd226,8'd254} : s = 15;
	{8'd226,8'd255} : s = 61;
	{8'd227,8'd0} : s = 346;
	{8'd227,8'd1} : s = 201;
	{8'd227,8'd2} : s = 345;
	{8'd227,8'd3} : s = 342;
	{8'd227,8'd4} : s = 459;
	{8'd227,8'd5} : s = 198;
	{8'd227,8'd6} : s = 341;
	{8'd227,8'd7} : s = 339;
	{8'd227,8'd8} : s = 455;
	{8'd227,8'd9} : s = 334;
	{8'd227,8'd10} : s = 444;
	{8'd227,8'd11} : s = 442;
	{8'd227,8'd12} : s = 502;
	{8'd227,8'd13} : s = 197;
	{8'd227,8'd14} : s = 333;
	{8'd227,8'd15} : s = 331;
	{8'd227,8'd16} : s = 441;
	{8'd227,8'd17} : s = 327;
	{8'd227,8'd18} : s = 438;
	{8'd227,8'd19} : s = 437;
	{8'd227,8'd20} : s = 501;
	{8'd227,8'd21} : s = 316;
	{8'd227,8'd22} : s = 435;
	{8'd227,8'd23} : s = 430;
	{8'd227,8'd24} : s = 499;
	{8'd227,8'd25} : s = 429;
	{8'd227,8'd26} : s = 494;
	{8'd227,8'd27} : s = 493;
	{8'd227,8'd28} : s = 510;
	{8'd227,8'd29} : s = 1;
	{8'd227,8'd30} : s = 18;
	{8'd227,8'd31} : s = 17;
	{8'd227,8'd32} : s = 82;
	{8'd227,8'd33} : s = 12;
	{8'd227,8'd34} : s = 81;
	{8'd227,8'd35} : s = 76;
	{8'd227,8'd36} : s = 195;
	{8'd227,8'd37} : s = 10;
	{8'd227,8'd38} : s = 74;
	{8'd227,8'd39} : s = 73;
	{8'd227,8'd40} : s = 184;
	{8'd227,8'd41} : s = 70;
	{8'd227,8'd42} : s = 180;
	{8'd227,8'd43} : s = 178;
	{8'd227,8'd44} : s = 314;
	{8'd227,8'd45} : s = 9;
	{8'd227,8'd46} : s = 69;
	{8'd227,8'd47} : s = 67;
	{8'd227,8'd48} : s = 177;
	{8'd227,8'd49} : s = 56;
	{8'd227,8'd50} : s = 172;
	{8'd227,8'd51} : s = 170;
	{8'd227,8'd52} : s = 313;
	{8'd227,8'd53} : s = 52;
	{8'd227,8'd54} : s = 169;
	{8'd227,8'd55} : s = 166;
	{8'd227,8'd56} : s = 310;
	{8'd227,8'd57} : s = 165;
	{8'd227,8'd58} : s = 309;
	{8'd227,8'd59} : s = 307;
	{8'd227,8'd60} : s = 427;
	{8'd227,8'd61} : s = 6;
	{8'd227,8'd62} : s = 50;
	{8'd227,8'd63} : s = 49;
	{8'd227,8'd64} : s = 163;
	{8'd227,8'd65} : s = 44;
	{8'd227,8'd66} : s = 156;
	{8'd227,8'd67} : s = 154;
	{8'd227,8'd68} : s = 302;
	{8'd227,8'd69} : s = 42;
	{8'd227,8'd70} : s = 153;
	{8'd227,8'd71} : s = 150;
	{8'd227,8'd72} : s = 301;
	{8'd227,8'd73} : s = 149;
	{8'd227,8'd74} : s = 299;
	{8'd227,8'd75} : s = 295;
	{8'd227,8'd76} : s = 423;
	{8'd227,8'd77} : s = 41;
	{8'd227,8'd78} : s = 147;
	{8'd227,8'd79} : s = 142;
	{8'd227,8'd80} : s = 286;
	{8'd227,8'd81} : s = 141;
	{8'd227,8'd82} : s = 285;
	{8'd227,8'd83} : s = 283;
	{8'd227,8'd84} : s = 414;
	{8'd227,8'd85} : s = 139;
	{8'd227,8'd86} : s = 279;
	{8'd227,8'd87} : s = 271;
	{8'd227,8'd88} : s = 413;
	{8'd227,8'd89} : s = 248;
	{8'd227,8'd90} : s = 411;
	{8'd227,8'd91} : s = 407;
	{8'd227,8'd92} : s = 491;
	{8'd227,8'd93} : s = 5;
	{8'd227,8'd94} : s = 38;
	{8'd227,8'd95} : s = 37;
	{8'd227,8'd96} : s = 135;
	{8'd227,8'd97} : s = 35;
	{8'd227,8'd98} : s = 120;
	{8'd227,8'd99} : s = 116;
	{8'd227,8'd100} : s = 244;
	{8'd227,8'd101} : s = 28;
	{8'd227,8'd102} : s = 114;
	{8'd227,8'd103} : s = 113;
	{8'd227,8'd104} : s = 242;
	{8'd227,8'd105} : s = 108;
	{8'd227,8'd106} : s = 241;
	{8'd227,8'd107} : s = 236;
	{8'd227,8'd108} : s = 399;
	{8'd227,8'd109} : s = 26;
	{8'd227,8'd110} : s = 106;
	{8'd227,8'd111} : s = 105;
	{8'd227,8'd112} : s = 234;
	{8'd227,8'd113} : s = 102;
	{8'd227,8'd114} : s = 233;
	{8'd227,8'd115} : s = 230;
	{8'd227,8'd116} : s = 380;
	{8'd227,8'd117} : s = 101;
	{8'd227,8'd118} : s = 229;
	{8'd227,8'd119} : s = 227;
	{8'd227,8'd120} : s = 378;
	{8'd227,8'd121} : s = 220;
	{8'd227,8'd122} : s = 377;
	{8'd227,8'd123} : s = 374;
	{8'd227,8'd124} : s = 487;
	{8'd227,8'd125} : s = 25;
	{8'd227,8'd126} : s = 99;
	{8'd227,8'd127} : s = 92;
	{8'd227,8'd128} : s = 218;
	{8'd227,8'd129} : s = 90;
	{8'd227,8'd130} : s = 217;
	{8'd227,8'd131} : s = 214;
	{8'd227,8'd132} : s = 373;
	{8'd227,8'd133} : s = 89;
	{8'd227,8'd134} : s = 213;
	{8'd227,8'd135} : s = 211;
	{8'd227,8'd136} : s = 371;
	{8'd227,8'd137} : s = 206;
	{8'd227,8'd138} : s = 366;
	{8'd227,8'd139} : s = 365;
	{8'd227,8'd140} : s = 478;
	{8'd227,8'd141} : s = 86;
	{8'd227,8'd142} : s = 205;
	{8'd227,8'd143} : s = 203;
	{8'd227,8'd144} : s = 363;
	{8'd227,8'd145} : s = 199;
	{8'd227,8'd146} : s = 359;
	{8'd227,8'd147} : s = 350;
	{8'd227,8'd148} : s = 477;
	{8'd227,8'd149} : s = 188;
	{8'd227,8'd150} : s = 349;
	{8'd227,8'd151} : s = 347;
	{8'd227,8'd152} : s = 475;
	{8'd227,8'd153} : s = 343;
	{8'd227,8'd154} : s = 471;
	{8'd227,8'd155} : s = 463;
	{8'd227,8'd156} : s = 509;
	{8'd227,8'd157} : s = 3;
	{8'd227,8'd158} : s = 22;
	{8'd227,8'd159} : s = 21;
	{8'd227,8'd160} : s = 85;
	{8'd227,8'd161} : s = 19;
	{8'd227,8'd162} : s = 83;
	{8'd227,8'd163} : s = 78;
	{8'd227,8'd164} : s = 186;
	{8'd227,8'd165} : s = 14;
	{8'd227,8'd166} : s = 77;
	{8'd227,8'd167} : s = 75;
	{8'd227,8'd168} : s = 185;
	{8'd227,8'd169} : s = 71;
	{8'd227,8'd170} : s = 182;
	{8'd227,8'd171} : s = 181;
	{8'd227,8'd172} : s = 335;
	{8'd227,8'd173} : s = 13;
	{8'd227,8'd174} : s = 60;
	{8'd227,8'd175} : s = 58;
	{8'd227,8'd176} : s = 179;
	{8'd227,8'd177} : s = 57;
	{8'd227,8'd178} : s = 174;
	{8'd227,8'd179} : s = 173;
	{8'd227,8'd180} : s = 318;
	{8'd227,8'd181} : s = 54;
	{8'd227,8'd182} : s = 171;
	{8'd227,8'd183} : s = 167;
	{8'd227,8'd184} : s = 317;
	{8'd227,8'd185} : s = 158;
	{8'd227,8'd186} : s = 315;
	{8'd227,8'd187} : s = 311;
	{8'd227,8'd188} : s = 446;
	{8'd227,8'd189} : s = 11;
	{8'd227,8'd190} : s = 53;
	{8'd227,8'd191} : s = 51;
	{8'd227,8'd192} : s = 157;
	{8'd227,8'd193} : s = 46;
	{8'd227,8'd194} : s = 155;
	{8'd227,8'd195} : s = 151;
	{8'd227,8'd196} : s = 303;
	{8'd227,8'd197} : s = 45;
	{8'd227,8'd198} : s = 143;
	{8'd227,8'd199} : s = 124;
	{8'd227,8'd200} : s = 287;
	{8'd227,8'd201} : s = 122;
	{8'd227,8'd202} : s = 252;
	{8'd227,8'd203} : s = 250;
	{8'd227,8'd204} : s = 445;
	{8'd227,8'd205} : s = 43;
	{8'd227,8'd206} : s = 121;
	{8'd227,8'd207} : s = 118;
	{8'd227,8'd208} : s = 249;
	{8'd227,8'd209} : s = 117;
	{8'd227,8'd210} : s = 246;
	{8'd227,8'd211} : s = 245;
	{8'd227,8'd212} : s = 443;
	{8'd227,8'd213} : s = 115;
	{8'd227,8'd214} : s = 243;
	{8'd227,8'd215} : s = 238;
	{8'd227,8'd216} : s = 439;
	{8'd227,8'd217} : s = 237;
	{8'd227,8'd218} : s = 431;
	{8'd227,8'd219} : s = 415;
	{8'd227,8'd220} : s = 507;
	{8'd227,8'd221} : s = 7;
	{8'd227,8'd222} : s = 39;
	{8'd227,8'd223} : s = 30;
	{8'd227,8'd224} : s = 110;
	{8'd227,8'd225} : s = 29;
	{8'd227,8'd226} : s = 109;
	{8'd227,8'd227} : s = 107;
	{8'd227,8'd228} : s = 235;
	{8'd227,8'd229} : s = 27;
	{8'd227,8'd230} : s = 103;
	{8'd227,8'd231} : s = 94;
	{8'd227,8'd232} : s = 231;
	{8'd227,8'd233} : s = 93;
	{8'd227,8'd234} : s = 222;
	{8'd227,8'd235} : s = 221;
	{8'd227,8'd236} : s = 382;
	{8'd227,8'd237} : s = 23;
	{8'd227,8'd238} : s = 91;
	{8'd227,8'd239} : s = 87;
	{8'd227,8'd240} : s = 219;
	{8'd227,8'd241} : s = 79;
	{8'd227,8'd242} : s = 215;
	{8'd227,8'd243} : s = 207;
	{8'd227,8'd244} : s = 381;
	{8'd227,8'd245} : s = 62;
	{8'd227,8'd246} : s = 190;
	{8'd227,8'd247} : s = 189;
	{8'd227,8'd248} : s = 379;
	{8'd227,8'd249} : s = 187;
	{8'd227,8'd250} : s = 375;
	{8'd227,8'd251} : s = 367;
	{8'd227,8'd252} : s = 503;
	{8'd227,8'd253} : s = 15;
	{8'd227,8'd254} : s = 61;
	{8'd227,8'd255} : s = 59;
	{8'd228,8'd0} : s = 201;
	{8'd228,8'd1} : s = 345;
	{8'd228,8'd2} : s = 342;
	{8'd228,8'd3} : s = 459;
	{8'd228,8'd4} : s = 198;
	{8'd228,8'd5} : s = 341;
	{8'd228,8'd6} : s = 339;
	{8'd228,8'd7} : s = 455;
	{8'd228,8'd8} : s = 334;
	{8'd228,8'd9} : s = 444;
	{8'd228,8'd10} : s = 442;
	{8'd228,8'd11} : s = 502;
	{8'd228,8'd12} : s = 197;
	{8'd228,8'd13} : s = 333;
	{8'd228,8'd14} : s = 331;
	{8'd228,8'd15} : s = 441;
	{8'd228,8'd16} : s = 327;
	{8'd228,8'd17} : s = 438;
	{8'd228,8'd18} : s = 437;
	{8'd228,8'd19} : s = 501;
	{8'd228,8'd20} : s = 316;
	{8'd228,8'd21} : s = 435;
	{8'd228,8'd22} : s = 430;
	{8'd228,8'd23} : s = 499;
	{8'd228,8'd24} : s = 429;
	{8'd228,8'd25} : s = 494;
	{8'd228,8'd26} : s = 493;
	{8'd228,8'd27} : s = 510;
	{8'd228,8'd28} : s = 1;
	{8'd228,8'd29} : s = 18;
	{8'd228,8'd30} : s = 17;
	{8'd228,8'd31} : s = 82;
	{8'd228,8'd32} : s = 12;
	{8'd228,8'd33} : s = 81;
	{8'd228,8'd34} : s = 76;
	{8'd228,8'd35} : s = 195;
	{8'd228,8'd36} : s = 10;
	{8'd228,8'd37} : s = 74;
	{8'd228,8'd38} : s = 73;
	{8'd228,8'd39} : s = 184;
	{8'd228,8'd40} : s = 70;
	{8'd228,8'd41} : s = 180;
	{8'd228,8'd42} : s = 178;
	{8'd228,8'd43} : s = 314;
	{8'd228,8'd44} : s = 9;
	{8'd228,8'd45} : s = 69;
	{8'd228,8'd46} : s = 67;
	{8'd228,8'd47} : s = 177;
	{8'd228,8'd48} : s = 56;
	{8'd228,8'd49} : s = 172;
	{8'd228,8'd50} : s = 170;
	{8'd228,8'd51} : s = 313;
	{8'd228,8'd52} : s = 52;
	{8'd228,8'd53} : s = 169;
	{8'd228,8'd54} : s = 166;
	{8'd228,8'd55} : s = 310;
	{8'd228,8'd56} : s = 165;
	{8'd228,8'd57} : s = 309;
	{8'd228,8'd58} : s = 307;
	{8'd228,8'd59} : s = 427;
	{8'd228,8'd60} : s = 6;
	{8'd228,8'd61} : s = 50;
	{8'd228,8'd62} : s = 49;
	{8'd228,8'd63} : s = 163;
	{8'd228,8'd64} : s = 44;
	{8'd228,8'd65} : s = 156;
	{8'd228,8'd66} : s = 154;
	{8'd228,8'd67} : s = 302;
	{8'd228,8'd68} : s = 42;
	{8'd228,8'd69} : s = 153;
	{8'd228,8'd70} : s = 150;
	{8'd228,8'd71} : s = 301;
	{8'd228,8'd72} : s = 149;
	{8'd228,8'd73} : s = 299;
	{8'd228,8'd74} : s = 295;
	{8'd228,8'd75} : s = 423;
	{8'd228,8'd76} : s = 41;
	{8'd228,8'd77} : s = 147;
	{8'd228,8'd78} : s = 142;
	{8'd228,8'd79} : s = 286;
	{8'd228,8'd80} : s = 141;
	{8'd228,8'd81} : s = 285;
	{8'd228,8'd82} : s = 283;
	{8'd228,8'd83} : s = 414;
	{8'd228,8'd84} : s = 139;
	{8'd228,8'd85} : s = 279;
	{8'd228,8'd86} : s = 271;
	{8'd228,8'd87} : s = 413;
	{8'd228,8'd88} : s = 248;
	{8'd228,8'd89} : s = 411;
	{8'd228,8'd90} : s = 407;
	{8'd228,8'd91} : s = 491;
	{8'd228,8'd92} : s = 5;
	{8'd228,8'd93} : s = 38;
	{8'd228,8'd94} : s = 37;
	{8'd228,8'd95} : s = 135;
	{8'd228,8'd96} : s = 35;
	{8'd228,8'd97} : s = 120;
	{8'd228,8'd98} : s = 116;
	{8'd228,8'd99} : s = 244;
	{8'd228,8'd100} : s = 28;
	{8'd228,8'd101} : s = 114;
	{8'd228,8'd102} : s = 113;
	{8'd228,8'd103} : s = 242;
	{8'd228,8'd104} : s = 108;
	{8'd228,8'd105} : s = 241;
	{8'd228,8'd106} : s = 236;
	{8'd228,8'd107} : s = 399;
	{8'd228,8'd108} : s = 26;
	{8'd228,8'd109} : s = 106;
	{8'd228,8'd110} : s = 105;
	{8'd228,8'd111} : s = 234;
	{8'd228,8'd112} : s = 102;
	{8'd228,8'd113} : s = 233;
	{8'd228,8'd114} : s = 230;
	{8'd228,8'd115} : s = 380;
	{8'd228,8'd116} : s = 101;
	{8'd228,8'd117} : s = 229;
	{8'd228,8'd118} : s = 227;
	{8'd228,8'd119} : s = 378;
	{8'd228,8'd120} : s = 220;
	{8'd228,8'd121} : s = 377;
	{8'd228,8'd122} : s = 374;
	{8'd228,8'd123} : s = 487;
	{8'd228,8'd124} : s = 25;
	{8'd228,8'd125} : s = 99;
	{8'd228,8'd126} : s = 92;
	{8'd228,8'd127} : s = 218;
	{8'd228,8'd128} : s = 90;
	{8'd228,8'd129} : s = 217;
	{8'd228,8'd130} : s = 214;
	{8'd228,8'd131} : s = 373;
	{8'd228,8'd132} : s = 89;
	{8'd228,8'd133} : s = 213;
	{8'd228,8'd134} : s = 211;
	{8'd228,8'd135} : s = 371;
	{8'd228,8'd136} : s = 206;
	{8'd228,8'd137} : s = 366;
	{8'd228,8'd138} : s = 365;
	{8'd228,8'd139} : s = 478;
	{8'd228,8'd140} : s = 86;
	{8'd228,8'd141} : s = 205;
	{8'd228,8'd142} : s = 203;
	{8'd228,8'd143} : s = 363;
	{8'd228,8'd144} : s = 199;
	{8'd228,8'd145} : s = 359;
	{8'd228,8'd146} : s = 350;
	{8'd228,8'd147} : s = 477;
	{8'd228,8'd148} : s = 188;
	{8'd228,8'd149} : s = 349;
	{8'd228,8'd150} : s = 347;
	{8'd228,8'd151} : s = 475;
	{8'd228,8'd152} : s = 343;
	{8'd228,8'd153} : s = 471;
	{8'd228,8'd154} : s = 463;
	{8'd228,8'd155} : s = 509;
	{8'd228,8'd156} : s = 3;
	{8'd228,8'd157} : s = 22;
	{8'd228,8'd158} : s = 21;
	{8'd228,8'd159} : s = 85;
	{8'd228,8'd160} : s = 19;
	{8'd228,8'd161} : s = 83;
	{8'd228,8'd162} : s = 78;
	{8'd228,8'd163} : s = 186;
	{8'd228,8'd164} : s = 14;
	{8'd228,8'd165} : s = 77;
	{8'd228,8'd166} : s = 75;
	{8'd228,8'd167} : s = 185;
	{8'd228,8'd168} : s = 71;
	{8'd228,8'd169} : s = 182;
	{8'd228,8'd170} : s = 181;
	{8'd228,8'd171} : s = 335;
	{8'd228,8'd172} : s = 13;
	{8'd228,8'd173} : s = 60;
	{8'd228,8'd174} : s = 58;
	{8'd228,8'd175} : s = 179;
	{8'd228,8'd176} : s = 57;
	{8'd228,8'd177} : s = 174;
	{8'd228,8'd178} : s = 173;
	{8'd228,8'd179} : s = 318;
	{8'd228,8'd180} : s = 54;
	{8'd228,8'd181} : s = 171;
	{8'd228,8'd182} : s = 167;
	{8'd228,8'd183} : s = 317;
	{8'd228,8'd184} : s = 158;
	{8'd228,8'd185} : s = 315;
	{8'd228,8'd186} : s = 311;
	{8'd228,8'd187} : s = 446;
	{8'd228,8'd188} : s = 11;
	{8'd228,8'd189} : s = 53;
	{8'd228,8'd190} : s = 51;
	{8'd228,8'd191} : s = 157;
	{8'd228,8'd192} : s = 46;
	{8'd228,8'd193} : s = 155;
	{8'd228,8'd194} : s = 151;
	{8'd228,8'd195} : s = 303;
	{8'd228,8'd196} : s = 45;
	{8'd228,8'd197} : s = 143;
	{8'd228,8'd198} : s = 124;
	{8'd228,8'd199} : s = 287;
	{8'd228,8'd200} : s = 122;
	{8'd228,8'd201} : s = 252;
	{8'd228,8'd202} : s = 250;
	{8'd228,8'd203} : s = 445;
	{8'd228,8'd204} : s = 43;
	{8'd228,8'd205} : s = 121;
	{8'd228,8'd206} : s = 118;
	{8'd228,8'd207} : s = 249;
	{8'd228,8'd208} : s = 117;
	{8'd228,8'd209} : s = 246;
	{8'd228,8'd210} : s = 245;
	{8'd228,8'd211} : s = 443;
	{8'd228,8'd212} : s = 115;
	{8'd228,8'd213} : s = 243;
	{8'd228,8'd214} : s = 238;
	{8'd228,8'd215} : s = 439;
	{8'd228,8'd216} : s = 237;
	{8'd228,8'd217} : s = 431;
	{8'd228,8'd218} : s = 415;
	{8'd228,8'd219} : s = 507;
	{8'd228,8'd220} : s = 7;
	{8'd228,8'd221} : s = 39;
	{8'd228,8'd222} : s = 30;
	{8'd228,8'd223} : s = 110;
	{8'd228,8'd224} : s = 29;
	{8'd228,8'd225} : s = 109;
	{8'd228,8'd226} : s = 107;
	{8'd228,8'd227} : s = 235;
	{8'd228,8'd228} : s = 27;
	{8'd228,8'd229} : s = 103;
	{8'd228,8'd230} : s = 94;
	{8'd228,8'd231} : s = 231;
	{8'd228,8'd232} : s = 93;
	{8'd228,8'd233} : s = 222;
	{8'd228,8'd234} : s = 221;
	{8'd228,8'd235} : s = 382;
	{8'd228,8'd236} : s = 23;
	{8'd228,8'd237} : s = 91;
	{8'd228,8'd238} : s = 87;
	{8'd228,8'd239} : s = 219;
	{8'd228,8'd240} : s = 79;
	{8'd228,8'd241} : s = 215;
	{8'd228,8'd242} : s = 207;
	{8'd228,8'd243} : s = 381;
	{8'd228,8'd244} : s = 62;
	{8'd228,8'd245} : s = 190;
	{8'd228,8'd246} : s = 189;
	{8'd228,8'd247} : s = 379;
	{8'd228,8'd248} : s = 187;
	{8'd228,8'd249} : s = 375;
	{8'd228,8'd250} : s = 367;
	{8'd228,8'd251} : s = 503;
	{8'd228,8'd252} : s = 15;
	{8'd228,8'd253} : s = 61;
	{8'd228,8'd254} : s = 59;
	{8'd228,8'd255} : s = 183;
	{8'd229,8'd0} : s = 345;
	{8'd229,8'd1} : s = 342;
	{8'd229,8'd2} : s = 459;
	{8'd229,8'd3} : s = 198;
	{8'd229,8'd4} : s = 341;
	{8'd229,8'd5} : s = 339;
	{8'd229,8'd6} : s = 455;
	{8'd229,8'd7} : s = 334;
	{8'd229,8'd8} : s = 444;
	{8'd229,8'd9} : s = 442;
	{8'd229,8'd10} : s = 502;
	{8'd229,8'd11} : s = 197;
	{8'd229,8'd12} : s = 333;
	{8'd229,8'd13} : s = 331;
	{8'd229,8'd14} : s = 441;
	{8'd229,8'd15} : s = 327;
	{8'd229,8'd16} : s = 438;
	{8'd229,8'd17} : s = 437;
	{8'd229,8'd18} : s = 501;
	{8'd229,8'd19} : s = 316;
	{8'd229,8'd20} : s = 435;
	{8'd229,8'd21} : s = 430;
	{8'd229,8'd22} : s = 499;
	{8'd229,8'd23} : s = 429;
	{8'd229,8'd24} : s = 494;
	{8'd229,8'd25} : s = 493;
	{8'd229,8'd26} : s = 510;
	{8'd229,8'd27} : s = 1;
	{8'd229,8'd28} : s = 18;
	{8'd229,8'd29} : s = 17;
	{8'd229,8'd30} : s = 82;
	{8'd229,8'd31} : s = 12;
	{8'd229,8'd32} : s = 81;
	{8'd229,8'd33} : s = 76;
	{8'd229,8'd34} : s = 195;
	{8'd229,8'd35} : s = 10;
	{8'd229,8'd36} : s = 74;
	{8'd229,8'd37} : s = 73;
	{8'd229,8'd38} : s = 184;
	{8'd229,8'd39} : s = 70;
	{8'd229,8'd40} : s = 180;
	{8'd229,8'd41} : s = 178;
	{8'd229,8'd42} : s = 314;
	{8'd229,8'd43} : s = 9;
	{8'd229,8'd44} : s = 69;
	{8'd229,8'd45} : s = 67;
	{8'd229,8'd46} : s = 177;
	{8'd229,8'd47} : s = 56;
	{8'd229,8'd48} : s = 172;
	{8'd229,8'd49} : s = 170;
	{8'd229,8'd50} : s = 313;
	{8'd229,8'd51} : s = 52;
	{8'd229,8'd52} : s = 169;
	{8'd229,8'd53} : s = 166;
	{8'd229,8'd54} : s = 310;
	{8'd229,8'd55} : s = 165;
	{8'd229,8'd56} : s = 309;
	{8'd229,8'd57} : s = 307;
	{8'd229,8'd58} : s = 427;
	{8'd229,8'd59} : s = 6;
	{8'd229,8'd60} : s = 50;
	{8'd229,8'd61} : s = 49;
	{8'd229,8'd62} : s = 163;
	{8'd229,8'd63} : s = 44;
	{8'd229,8'd64} : s = 156;
	{8'd229,8'd65} : s = 154;
	{8'd229,8'd66} : s = 302;
	{8'd229,8'd67} : s = 42;
	{8'd229,8'd68} : s = 153;
	{8'd229,8'd69} : s = 150;
	{8'd229,8'd70} : s = 301;
	{8'd229,8'd71} : s = 149;
	{8'd229,8'd72} : s = 299;
	{8'd229,8'd73} : s = 295;
	{8'd229,8'd74} : s = 423;
	{8'd229,8'd75} : s = 41;
	{8'd229,8'd76} : s = 147;
	{8'd229,8'd77} : s = 142;
	{8'd229,8'd78} : s = 286;
	{8'd229,8'd79} : s = 141;
	{8'd229,8'd80} : s = 285;
	{8'd229,8'd81} : s = 283;
	{8'd229,8'd82} : s = 414;
	{8'd229,8'd83} : s = 139;
	{8'd229,8'd84} : s = 279;
	{8'd229,8'd85} : s = 271;
	{8'd229,8'd86} : s = 413;
	{8'd229,8'd87} : s = 248;
	{8'd229,8'd88} : s = 411;
	{8'd229,8'd89} : s = 407;
	{8'd229,8'd90} : s = 491;
	{8'd229,8'd91} : s = 5;
	{8'd229,8'd92} : s = 38;
	{8'd229,8'd93} : s = 37;
	{8'd229,8'd94} : s = 135;
	{8'd229,8'd95} : s = 35;
	{8'd229,8'd96} : s = 120;
	{8'd229,8'd97} : s = 116;
	{8'd229,8'd98} : s = 244;
	{8'd229,8'd99} : s = 28;
	{8'd229,8'd100} : s = 114;
	{8'd229,8'd101} : s = 113;
	{8'd229,8'd102} : s = 242;
	{8'd229,8'd103} : s = 108;
	{8'd229,8'd104} : s = 241;
	{8'd229,8'd105} : s = 236;
	{8'd229,8'd106} : s = 399;
	{8'd229,8'd107} : s = 26;
	{8'd229,8'd108} : s = 106;
	{8'd229,8'd109} : s = 105;
	{8'd229,8'd110} : s = 234;
	{8'd229,8'd111} : s = 102;
	{8'd229,8'd112} : s = 233;
	{8'd229,8'd113} : s = 230;
	{8'd229,8'd114} : s = 380;
	{8'd229,8'd115} : s = 101;
	{8'd229,8'd116} : s = 229;
	{8'd229,8'd117} : s = 227;
	{8'd229,8'd118} : s = 378;
	{8'd229,8'd119} : s = 220;
	{8'd229,8'd120} : s = 377;
	{8'd229,8'd121} : s = 374;
	{8'd229,8'd122} : s = 487;
	{8'd229,8'd123} : s = 25;
	{8'd229,8'd124} : s = 99;
	{8'd229,8'd125} : s = 92;
	{8'd229,8'd126} : s = 218;
	{8'd229,8'd127} : s = 90;
	{8'd229,8'd128} : s = 217;
	{8'd229,8'd129} : s = 214;
	{8'd229,8'd130} : s = 373;
	{8'd229,8'd131} : s = 89;
	{8'd229,8'd132} : s = 213;
	{8'd229,8'd133} : s = 211;
	{8'd229,8'd134} : s = 371;
	{8'd229,8'd135} : s = 206;
	{8'd229,8'd136} : s = 366;
	{8'd229,8'd137} : s = 365;
	{8'd229,8'd138} : s = 478;
	{8'd229,8'd139} : s = 86;
	{8'd229,8'd140} : s = 205;
	{8'd229,8'd141} : s = 203;
	{8'd229,8'd142} : s = 363;
	{8'd229,8'd143} : s = 199;
	{8'd229,8'd144} : s = 359;
	{8'd229,8'd145} : s = 350;
	{8'd229,8'd146} : s = 477;
	{8'd229,8'd147} : s = 188;
	{8'd229,8'd148} : s = 349;
	{8'd229,8'd149} : s = 347;
	{8'd229,8'd150} : s = 475;
	{8'd229,8'd151} : s = 343;
	{8'd229,8'd152} : s = 471;
	{8'd229,8'd153} : s = 463;
	{8'd229,8'd154} : s = 509;
	{8'd229,8'd155} : s = 3;
	{8'd229,8'd156} : s = 22;
	{8'd229,8'd157} : s = 21;
	{8'd229,8'd158} : s = 85;
	{8'd229,8'd159} : s = 19;
	{8'd229,8'd160} : s = 83;
	{8'd229,8'd161} : s = 78;
	{8'd229,8'd162} : s = 186;
	{8'd229,8'd163} : s = 14;
	{8'd229,8'd164} : s = 77;
	{8'd229,8'd165} : s = 75;
	{8'd229,8'd166} : s = 185;
	{8'd229,8'd167} : s = 71;
	{8'd229,8'd168} : s = 182;
	{8'd229,8'd169} : s = 181;
	{8'd229,8'd170} : s = 335;
	{8'd229,8'd171} : s = 13;
	{8'd229,8'd172} : s = 60;
	{8'd229,8'd173} : s = 58;
	{8'd229,8'd174} : s = 179;
	{8'd229,8'd175} : s = 57;
	{8'd229,8'd176} : s = 174;
	{8'd229,8'd177} : s = 173;
	{8'd229,8'd178} : s = 318;
	{8'd229,8'd179} : s = 54;
	{8'd229,8'd180} : s = 171;
	{8'd229,8'd181} : s = 167;
	{8'd229,8'd182} : s = 317;
	{8'd229,8'd183} : s = 158;
	{8'd229,8'd184} : s = 315;
	{8'd229,8'd185} : s = 311;
	{8'd229,8'd186} : s = 446;
	{8'd229,8'd187} : s = 11;
	{8'd229,8'd188} : s = 53;
	{8'd229,8'd189} : s = 51;
	{8'd229,8'd190} : s = 157;
	{8'd229,8'd191} : s = 46;
	{8'd229,8'd192} : s = 155;
	{8'd229,8'd193} : s = 151;
	{8'd229,8'd194} : s = 303;
	{8'd229,8'd195} : s = 45;
	{8'd229,8'd196} : s = 143;
	{8'd229,8'd197} : s = 124;
	{8'd229,8'd198} : s = 287;
	{8'd229,8'd199} : s = 122;
	{8'd229,8'd200} : s = 252;
	{8'd229,8'd201} : s = 250;
	{8'd229,8'd202} : s = 445;
	{8'd229,8'd203} : s = 43;
	{8'd229,8'd204} : s = 121;
	{8'd229,8'd205} : s = 118;
	{8'd229,8'd206} : s = 249;
	{8'd229,8'd207} : s = 117;
	{8'd229,8'd208} : s = 246;
	{8'd229,8'd209} : s = 245;
	{8'd229,8'd210} : s = 443;
	{8'd229,8'd211} : s = 115;
	{8'd229,8'd212} : s = 243;
	{8'd229,8'd213} : s = 238;
	{8'd229,8'd214} : s = 439;
	{8'd229,8'd215} : s = 237;
	{8'd229,8'd216} : s = 431;
	{8'd229,8'd217} : s = 415;
	{8'd229,8'd218} : s = 507;
	{8'd229,8'd219} : s = 7;
	{8'd229,8'd220} : s = 39;
	{8'd229,8'd221} : s = 30;
	{8'd229,8'd222} : s = 110;
	{8'd229,8'd223} : s = 29;
	{8'd229,8'd224} : s = 109;
	{8'd229,8'd225} : s = 107;
	{8'd229,8'd226} : s = 235;
	{8'd229,8'd227} : s = 27;
	{8'd229,8'd228} : s = 103;
	{8'd229,8'd229} : s = 94;
	{8'd229,8'd230} : s = 231;
	{8'd229,8'd231} : s = 93;
	{8'd229,8'd232} : s = 222;
	{8'd229,8'd233} : s = 221;
	{8'd229,8'd234} : s = 382;
	{8'd229,8'd235} : s = 23;
	{8'd229,8'd236} : s = 91;
	{8'd229,8'd237} : s = 87;
	{8'd229,8'd238} : s = 219;
	{8'd229,8'd239} : s = 79;
	{8'd229,8'd240} : s = 215;
	{8'd229,8'd241} : s = 207;
	{8'd229,8'd242} : s = 381;
	{8'd229,8'd243} : s = 62;
	{8'd229,8'd244} : s = 190;
	{8'd229,8'd245} : s = 189;
	{8'd229,8'd246} : s = 379;
	{8'd229,8'd247} : s = 187;
	{8'd229,8'd248} : s = 375;
	{8'd229,8'd249} : s = 367;
	{8'd229,8'd250} : s = 503;
	{8'd229,8'd251} : s = 15;
	{8'd229,8'd252} : s = 61;
	{8'd229,8'd253} : s = 59;
	{8'd229,8'd254} : s = 183;
	{8'd229,8'd255} : s = 55;
	{8'd230,8'd0} : s = 342;
	{8'd230,8'd1} : s = 459;
	{8'd230,8'd2} : s = 198;
	{8'd230,8'd3} : s = 341;
	{8'd230,8'd4} : s = 339;
	{8'd230,8'd5} : s = 455;
	{8'd230,8'd6} : s = 334;
	{8'd230,8'd7} : s = 444;
	{8'd230,8'd8} : s = 442;
	{8'd230,8'd9} : s = 502;
	{8'd230,8'd10} : s = 197;
	{8'd230,8'd11} : s = 333;
	{8'd230,8'd12} : s = 331;
	{8'd230,8'd13} : s = 441;
	{8'd230,8'd14} : s = 327;
	{8'd230,8'd15} : s = 438;
	{8'd230,8'd16} : s = 437;
	{8'd230,8'd17} : s = 501;
	{8'd230,8'd18} : s = 316;
	{8'd230,8'd19} : s = 435;
	{8'd230,8'd20} : s = 430;
	{8'd230,8'd21} : s = 499;
	{8'd230,8'd22} : s = 429;
	{8'd230,8'd23} : s = 494;
	{8'd230,8'd24} : s = 493;
	{8'd230,8'd25} : s = 510;
	{8'd230,8'd26} : s = 1;
	{8'd230,8'd27} : s = 18;
	{8'd230,8'd28} : s = 17;
	{8'd230,8'd29} : s = 82;
	{8'd230,8'd30} : s = 12;
	{8'd230,8'd31} : s = 81;
	{8'd230,8'd32} : s = 76;
	{8'd230,8'd33} : s = 195;
	{8'd230,8'd34} : s = 10;
	{8'd230,8'd35} : s = 74;
	{8'd230,8'd36} : s = 73;
	{8'd230,8'd37} : s = 184;
	{8'd230,8'd38} : s = 70;
	{8'd230,8'd39} : s = 180;
	{8'd230,8'd40} : s = 178;
	{8'd230,8'd41} : s = 314;
	{8'd230,8'd42} : s = 9;
	{8'd230,8'd43} : s = 69;
	{8'd230,8'd44} : s = 67;
	{8'd230,8'd45} : s = 177;
	{8'd230,8'd46} : s = 56;
	{8'd230,8'd47} : s = 172;
	{8'd230,8'd48} : s = 170;
	{8'd230,8'd49} : s = 313;
	{8'd230,8'd50} : s = 52;
	{8'd230,8'd51} : s = 169;
	{8'd230,8'd52} : s = 166;
	{8'd230,8'd53} : s = 310;
	{8'd230,8'd54} : s = 165;
	{8'd230,8'd55} : s = 309;
	{8'd230,8'd56} : s = 307;
	{8'd230,8'd57} : s = 427;
	{8'd230,8'd58} : s = 6;
	{8'd230,8'd59} : s = 50;
	{8'd230,8'd60} : s = 49;
	{8'd230,8'd61} : s = 163;
	{8'd230,8'd62} : s = 44;
	{8'd230,8'd63} : s = 156;
	{8'd230,8'd64} : s = 154;
	{8'd230,8'd65} : s = 302;
	{8'd230,8'd66} : s = 42;
	{8'd230,8'd67} : s = 153;
	{8'd230,8'd68} : s = 150;
	{8'd230,8'd69} : s = 301;
	{8'd230,8'd70} : s = 149;
	{8'd230,8'd71} : s = 299;
	{8'd230,8'd72} : s = 295;
	{8'd230,8'd73} : s = 423;
	{8'd230,8'd74} : s = 41;
	{8'd230,8'd75} : s = 147;
	{8'd230,8'd76} : s = 142;
	{8'd230,8'd77} : s = 286;
	{8'd230,8'd78} : s = 141;
	{8'd230,8'd79} : s = 285;
	{8'd230,8'd80} : s = 283;
	{8'd230,8'd81} : s = 414;
	{8'd230,8'd82} : s = 139;
	{8'd230,8'd83} : s = 279;
	{8'd230,8'd84} : s = 271;
	{8'd230,8'd85} : s = 413;
	{8'd230,8'd86} : s = 248;
	{8'd230,8'd87} : s = 411;
	{8'd230,8'd88} : s = 407;
	{8'd230,8'd89} : s = 491;
	{8'd230,8'd90} : s = 5;
	{8'd230,8'd91} : s = 38;
	{8'd230,8'd92} : s = 37;
	{8'd230,8'd93} : s = 135;
	{8'd230,8'd94} : s = 35;
	{8'd230,8'd95} : s = 120;
	{8'd230,8'd96} : s = 116;
	{8'd230,8'd97} : s = 244;
	{8'd230,8'd98} : s = 28;
	{8'd230,8'd99} : s = 114;
	{8'd230,8'd100} : s = 113;
	{8'd230,8'd101} : s = 242;
	{8'd230,8'd102} : s = 108;
	{8'd230,8'd103} : s = 241;
	{8'd230,8'd104} : s = 236;
	{8'd230,8'd105} : s = 399;
	{8'd230,8'd106} : s = 26;
	{8'd230,8'd107} : s = 106;
	{8'd230,8'd108} : s = 105;
	{8'd230,8'd109} : s = 234;
	{8'd230,8'd110} : s = 102;
	{8'd230,8'd111} : s = 233;
	{8'd230,8'd112} : s = 230;
	{8'd230,8'd113} : s = 380;
	{8'd230,8'd114} : s = 101;
	{8'd230,8'd115} : s = 229;
	{8'd230,8'd116} : s = 227;
	{8'd230,8'd117} : s = 378;
	{8'd230,8'd118} : s = 220;
	{8'd230,8'd119} : s = 377;
	{8'd230,8'd120} : s = 374;
	{8'd230,8'd121} : s = 487;
	{8'd230,8'd122} : s = 25;
	{8'd230,8'd123} : s = 99;
	{8'd230,8'd124} : s = 92;
	{8'd230,8'd125} : s = 218;
	{8'd230,8'd126} : s = 90;
	{8'd230,8'd127} : s = 217;
	{8'd230,8'd128} : s = 214;
	{8'd230,8'd129} : s = 373;
	{8'd230,8'd130} : s = 89;
	{8'd230,8'd131} : s = 213;
	{8'd230,8'd132} : s = 211;
	{8'd230,8'd133} : s = 371;
	{8'd230,8'd134} : s = 206;
	{8'd230,8'd135} : s = 366;
	{8'd230,8'd136} : s = 365;
	{8'd230,8'd137} : s = 478;
	{8'd230,8'd138} : s = 86;
	{8'd230,8'd139} : s = 205;
	{8'd230,8'd140} : s = 203;
	{8'd230,8'd141} : s = 363;
	{8'd230,8'd142} : s = 199;
	{8'd230,8'd143} : s = 359;
	{8'd230,8'd144} : s = 350;
	{8'd230,8'd145} : s = 477;
	{8'd230,8'd146} : s = 188;
	{8'd230,8'd147} : s = 349;
	{8'd230,8'd148} : s = 347;
	{8'd230,8'd149} : s = 475;
	{8'd230,8'd150} : s = 343;
	{8'd230,8'd151} : s = 471;
	{8'd230,8'd152} : s = 463;
	{8'd230,8'd153} : s = 509;
	{8'd230,8'd154} : s = 3;
	{8'd230,8'd155} : s = 22;
	{8'd230,8'd156} : s = 21;
	{8'd230,8'd157} : s = 85;
	{8'd230,8'd158} : s = 19;
	{8'd230,8'd159} : s = 83;
	{8'd230,8'd160} : s = 78;
	{8'd230,8'd161} : s = 186;
	{8'd230,8'd162} : s = 14;
	{8'd230,8'd163} : s = 77;
	{8'd230,8'd164} : s = 75;
	{8'd230,8'd165} : s = 185;
	{8'd230,8'd166} : s = 71;
	{8'd230,8'd167} : s = 182;
	{8'd230,8'd168} : s = 181;
	{8'd230,8'd169} : s = 335;
	{8'd230,8'd170} : s = 13;
	{8'd230,8'd171} : s = 60;
	{8'd230,8'd172} : s = 58;
	{8'd230,8'd173} : s = 179;
	{8'd230,8'd174} : s = 57;
	{8'd230,8'd175} : s = 174;
	{8'd230,8'd176} : s = 173;
	{8'd230,8'd177} : s = 318;
	{8'd230,8'd178} : s = 54;
	{8'd230,8'd179} : s = 171;
	{8'd230,8'd180} : s = 167;
	{8'd230,8'd181} : s = 317;
	{8'd230,8'd182} : s = 158;
	{8'd230,8'd183} : s = 315;
	{8'd230,8'd184} : s = 311;
	{8'd230,8'd185} : s = 446;
	{8'd230,8'd186} : s = 11;
	{8'd230,8'd187} : s = 53;
	{8'd230,8'd188} : s = 51;
	{8'd230,8'd189} : s = 157;
	{8'd230,8'd190} : s = 46;
	{8'd230,8'd191} : s = 155;
	{8'd230,8'd192} : s = 151;
	{8'd230,8'd193} : s = 303;
	{8'd230,8'd194} : s = 45;
	{8'd230,8'd195} : s = 143;
	{8'd230,8'd196} : s = 124;
	{8'd230,8'd197} : s = 287;
	{8'd230,8'd198} : s = 122;
	{8'd230,8'd199} : s = 252;
	{8'd230,8'd200} : s = 250;
	{8'd230,8'd201} : s = 445;
	{8'd230,8'd202} : s = 43;
	{8'd230,8'd203} : s = 121;
	{8'd230,8'd204} : s = 118;
	{8'd230,8'd205} : s = 249;
	{8'd230,8'd206} : s = 117;
	{8'd230,8'd207} : s = 246;
	{8'd230,8'd208} : s = 245;
	{8'd230,8'd209} : s = 443;
	{8'd230,8'd210} : s = 115;
	{8'd230,8'd211} : s = 243;
	{8'd230,8'd212} : s = 238;
	{8'd230,8'd213} : s = 439;
	{8'd230,8'd214} : s = 237;
	{8'd230,8'd215} : s = 431;
	{8'd230,8'd216} : s = 415;
	{8'd230,8'd217} : s = 507;
	{8'd230,8'd218} : s = 7;
	{8'd230,8'd219} : s = 39;
	{8'd230,8'd220} : s = 30;
	{8'd230,8'd221} : s = 110;
	{8'd230,8'd222} : s = 29;
	{8'd230,8'd223} : s = 109;
	{8'd230,8'd224} : s = 107;
	{8'd230,8'd225} : s = 235;
	{8'd230,8'd226} : s = 27;
	{8'd230,8'd227} : s = 103;
	{8'd230,8'd228} : s = 94;
	{8'd230,8'd229} : s = 231;
	{8'd230,8'd230} : s = 93;
	{8'd230,8'd231} : s = 222;
	{8'd230,8'd232} : s = 221;
	{8'd230,8'd233} : s = 382;
	{8'd230,8'd234} : s = 23;
	{8'd230,8'd235} : s = 91;
	{8'd230,8'd236} : s = 87;
	{8'd230,8'd237} : s = 219;
	{8'd230,8'd238} : s = 79;
	{8'd230,8'd239} : s = 215;
	{8'd230,8'd240} : s = 207;
	{8'd230,8'd241} : s = 381;
	{8'd230,8'd242} : s = 62;
	{8'd230,8'd243} : s = 190;
	{8'd230,8'd244} : s = 189;
	{8'd230,8'd245} : s = 379;
	{8'd230,8'd246} : s = 187;
	{8'd230,8'd247} : s = 375;
	{8'd230,8'd248} : s = 367;
	{8'd230,8'd249} : s = 503;
	{8'd230,8'd250} : s = 15;
	{8'd230,8'd251} : s = 61;
	{8'd230,8'd252} : s = 59;
	{8'd230,8'd253} : s = 183;
	{8'd230,8'd254} : s = 55;
	{8'd230,8'd255} : s = 175;
	{8'd231,8'd0} : s = 459;
	{8'd231,8'd1} : s = 198;
	{8'd231,8'd2} : s = 341;
	{8'd231,8'd3} : s = 339;
	{8'd231,8'd4} : s = 455;
	{8'd231,8'd5} : s = 334;
	{8'd231,8'd6} : s = 444;
	{8'd231,8'd7} : s = 442;
	{8'd231,8'd8} : s = 502;
	{8'd231,8'd9} : s = 197;
	{8'd231,8'd10} : s = 333;
	{8'd231,8'd11} : s = 331;
	{8'd231,8'd12} : s = 441;
	{8'd231,8'd13} : s = 327;
	{8'd231,8'd14} : s = 438;
	{8'd231,8'd15} : s = 437;
	{8'd231,8'd16} : s = 501;
	{8'd231,8'd17} : s = 316;
	{8'd231,8'd18} : s = 435;
	{8'd231,8'd19} : s = 430;
	{8'd231,8'd20} : s = 499;
	{8'd231,8'd21} : s = 429;
	{8'd231,8'd22} : s = 494;
	{8'd231,8'd23} : s = 493;
	{8'd231,8'd24} : s = 510;
	{8'd231,8'd25} : s = 1;
	{8'd231,8'd26} : s = 18;
	{8'd231,8'd27} : s = 17;
	{8'd231,8'd28} : s = 82;
	{8'd231,8'd29} : s = 12;
	{8'd231,8'd30} : s = 81;
	{8'd231,8'd31} : s = 76;
	{8'd231,8'd32} : s = 195;
	{8'd231,8'd33} : s = 10;
	{8'd231,8'd34} : s = 74;
	{8'd231,8'd35} : s = 73;
	{8'd231,8'd36} : s = 184;
	{8'd231,8'd37} : s = 70;
	{8'd231,8'd38} : s = 180;
	{8'd231,8'd39} : s = 178;
	{8'd231,8'd40} : s = 314;
	{8'd231,8'd41} : s = 9;
	{8'd231,8'd42} : s = 69;
	{8'd231,8'd43} : s = 67;
	{8'd231,8'd44} : s = 177;
	{8'd231,8'd45} : s = 56;
	{8'd231,8'd46} : s = 172;
	{8'd231,8'd47} : s = 170;
	{8'd231,8'd48} : s = 313;
	{8'd231,8'd49} : s = 52;
	{8'd231,8'd50} : s = 169;
	{8'd231,8'd51} : s = 166;
	{8'd231,8'd52} : s = 310;
	{8'd231,8'd53} : s = 165;
	{8'd231,8'd54} : s = 309;
	{8'd231,8'd55} : s = 307;
	{8'd231,8'd56} : s = 427;
	{8'd231,8'd57} : s = 6;
	{8'd231,8'd58} : s = 50;
	{8'd231,8'd59} : s = 49;
	{8'd231,8'd60} : s = 163;
	{8'd231,8'd61} : s = 44;
	{8'd231,8'd62} : s = 156;
	{8'd231,8'd63} : s = 154;
	{8'd231,8'd64} : s = 302;
	{8'd231,8'd65} : s = 42;
	{8'd231,8'd66} : s = 153;
	{8'd231,8'd67} : s = 150;
	{8'd231,8'd68} : s = 301;
	{8'd231,8'd69} : s = 149;
	{8'd231,8'd70} : s = 299;
	{8'd231,8'd71} : s = 295;
	{8'd231,8'd72} : s = 423;
	{8'd231,8'd73} : s = 41;
	{8'd231,8'd74} : s = 147;
	{8'd231,8'd75} : s = 142;
	{8'd231,8'd76} : s = 286;
	{8'd231,8'd77} : s = 141;
	{8'd231,8'd78} : s = 285;
	{8'd231,8'd79} : s = 283;
	{8'd231,8'd80} : s = 414;
	{8'd231,8'd81} : s = 139;
	{8'd231,8'd82} : s = 279;
	{8'd231,8'd83} : s = 271;
	{8'd231,8'd84} : s = 413;
	{8'd231,8'd85} : s = 248;
	{8'd231,8'd86} : s = 411;
	{8'd231,8'd87} : s = 407;
	{8'd231,8'd88} : s = 491;
	{8'd231,8'd89} : s = 5;
	{8'd231,8'd90} : s = 38;
	{8'd231,8'd91} : s = 37;
	{8'd231,8'd92} : s = 135;
	{8'd231,8'd93} : s = 35;
	{8'd231,8'd94} : s = 120;
	{8'd231,8'd95} : s = 116;
	{8'd231,8'd96} : s = 244;
	{8'd231,8'd97} : s = 28;
	{8'd231,8'd98} : s = 114;
	{8'd231,8'd99} : s = 113;
	{8'd231,8'd100} : s = 242;
	{8'd231,8'd101} : s = 108;
	{8'd231,8'd102} : s = 241;
	{8'd231,8'd103} : s = 236;
	{8'd231,8'd104} : s = 399;
	{8'd231,8'd105} : s = 26;
	{8'd231,8'd106} : s = 106;
	{8'd231,8'd107} : s = 105;
	{8'd231,8'd108} : s = 234;
	{8'd231,8'd109} : s = 102;
	{8'd231,8'd110} : s = 233;
	{8'd231,8'd111} : s = 230;
	{8'd231,8'd112} : s = 380;
	{8'd231,8'd113} : s = 101;
	{8'd231,8'd114} : s = 229;
	{8'd231,8'd115} : s = 227;
	{8'd231,8'd116} : s = 378;
	{8'd231,8'd117} : s = 220;
	{8'd231,8'd118} : s = 377;
	{8'd231,8'd119} : s = 374;
	{8'd231,8'd120} : s = 487;
	{8'd231,8'd121} : s = 25;
	{8'd231,8'd122} : s = 99;
	{8'd231,8'd123} : s = 92;
	{8'd231,8'd124} : s = 218;
	{8'd231,8'd125} : s = 90;
	{8'd231,8'd126} : s = 217;
	{8'd231,8'd127} : s = 214;
	{8'd231,8'd128} : s = 373;
	{8'd231,8'd129} : s = 89;
	{8'd231,8'd130} : s = 213;
	{8'd231,8'd131} : s = 211;
	{8'd231,8'd132} : s = 371;
	{8'd231,8'd133} : s = 206;
	{8'd231,8'd134} : s = 366;
	{8'd231,8'd135} : s = 365;
	{8'd231,8'd136} : s = 478;
	{8'd231,8'd137} : s = 86;
	{8'd231,8'd138} : s = 205;
	{8'd231,8'd139} : s = 203;
	{8'd231,8'd140} : s = 363;
	{8'd231,8'd141} : s = 199;
	{8'd231,8'd142} : s = 359;
	{8'd231,8'd143} : s = 350;
	{8'd231,8'd144} : s = 477;
	{8'd231,8'd145} : s = 188;
	{8'd231,8'd146} : s = 349;
	{8'd231,8'd147} : s = 347;
	{8'd231,8'd148} : s = 475;
	{8'd231,8'd149} : s = 343;
	{8'd231,8'd150} : s = 471;
	{8'd231,8'd151} : s = 463;
	{8'd231,8'd152} : s = 509;
	{8'd231,8'd153} : s = 3;
	{8'd231,8'd154} : s = 22;
	{8'd231,8'd155} : s = 21;
	{8'd231,8'd156} : s = 85;
	{8'd231,8'd157} : s = 19;
	{8'd231,8'd158} : s = 83;
	{8'd231,8'd159} : s = 78;
	{8'd231,8'd160} : s = 186;
	{8'd231,8'd161} : s = 14;
	{8'd231,8'd162} : s = 77;
	{8'd231,8'd163} : s = 75;
	{8'd231,8'd164} : s = 185;
	{8'd231,8'd165} : s = 71;
	{8'd231,8'd166} : s = 182;
	{8'd231,8'd167} : s = 181;
	{8'd231,8'd168} : s = 335;
	{8'd231,8'd169} : s = 13;
	{8'd231,8'd170} : s = 60;
	{8'd231,8'd171} : s = 58;
	{8'd231,8'd172} : s = 179;
	{8'd231,8'd173} : s = 57;
	{8'd231,8'd174} : s = 174;
	{8'd231,8'd175} : s = 173;
	{8'd231,8'd176} : s = 318;
	{8'd231,8'd177} : s = 54;
	{8'd231,8'd178} : s = 171;
	{8'd231,8'd179} : s = 167;
	{8'd231,8'd180} : s = 317;
	{8'd231,8'd181} : s = 158;
	{8'd231,8'd182} : s = 315;
	{8'd231,8'd183} : s = 311;
	{8'd231,8'd184} : s = 446;
	{8'd231,8'd185} : s = 11;
	{8'd231,8'd186} : s = 53;
	{8'd231,8'd187} : s = 51;
	{8'd231,8'd188} : s = 157;
	{8'd231,8'd189} : s = 46;
	{8'd231,8'd190} : s = 155;
	{8'd231,8'd191} : s = 151;
	{8'd231,8'd192} : s = 303;
	{8'd231,8'd193} : s = 45;
	{8'd231,8'd194} : s = 143;
	{8'd231,8'd195} : s = 124;
	{8'd231,8'd196} : s = 287;
	{8'd231,8'd197} : s = 122;
	{8'd231,8'd198} : s = 252;
	{8'd231,8'd199} : s = 250;
	{8'd231,8'd200} : s = 445;
	{8'd231,8'd201} : s = 43;
	{8'd231,8'd202} : s = 121;
	{8'd231,8'd203} : s = 118;
	{8'd231,8'd204} : s = 249;
	{8'd231,8'd205} : s = 117;
	{8'd231,8'd206} : s = 246;
	{8'd231,8'd207} : s = 245;
	{8'd231,8'd208} : s = 443;
	{8'd231,8'd209} : s = 115;
	{8'd231,8'd210} : s = 243;
	{8'd231,8'd211} : s = 238;
	{8'd231,8'd212} : s = 439;
	{8'd231,8'd213} : s = 237;
	{8'd231,8'd214} : s = 431;
	{8'd231,8'd215} : s = 415;
	{8'd231,8'd216} : s = 507;
	{8'd231,8'd217} : s = 7;
	{8'd231,8'd218} : s = 39;
	{8'd231,8'd219} : s = 30;
	{8'd231,8'd220} : s = 110;
	{8'd231,8'd221} : s = 29;
	{8'd231,8'd222} : s = 109;
	{8'd231,8'd223} : s = 107;
	{8'd231,8'd224} : s = 235;
	{8'd231,8'd225} : s = 27;
	{8'd231,8'd226} : s = 103;
	{8'd231,8'd227} : s = 94;
	{8'd231,8'd228} : s = 231;
	{8'd231,8'd229} : s = 93;
	{8'd231,8'd230} : s = 222;
	{8'd231,8'd231} : s = 221;
	{8'd231,8'd232} : s = 382;
	{8'd231,8'd233} : s = 23;
	{8'd231,8'd234} : s = 91;
	{8'd231,8'd235} : s = 87;
	{8'd231,8'd236} : s = 219;
	{8'd231,8'd237} : s = 79;
	{8'd231,8'd238} : s = 215;
	{8'd231,8'd239} : s = 207;
	{8'd231,8'd240} : s = 381;
	{8'd231,8'd241} : s = 62;
	{8'd231,8'd242} : s = 190;
	{8'd231,8'd243} : s = 189;
	{8'd231,8'd244} : s = 379;
	{8'd231,8'd245} : s = 187;
	{8'd231,8'd246} : s = 375;
	{8'd231,8'd247} : s = 367;
	{8'd231,8'd248} : s = 503;
	{8'd231,8'd249} : s = 15;
	{8'd231,8'd250} : s = 61;
	{8'd231,8'd251} : s = 59;
	{8'd231,8'd252} : s = 183;
	{8'd231,8'd253} : s = 55;
	{8'd231,8'd254} : s = 175;
	{8'd231,8'd255} : s = 159;
	{8'd232,8'd0} : s = 198;
	{8'd232,8'd1} : s = 341;
	{8'd232,8'd2} : s = 339;
	{8'd232,8'd3} : s = 455;
	{8'd232,8'd4} : s = 334;
	{8'd232,8'd5} : s = 444;
	{8'd232,8'd6} : s = 442;
	{8'd232,8'd7} : s = 502;
	{8'd232,8'd8} : s = 197;
	{8'd232,8'd9} : s = 333;
	{8'd232,8'd10} : s = 331;
	{8'd232,8'd11} : s = 441;
	{8'd232,8'd12} : s = 327;
	{8'd232,8'd13} : s = 438;
	{8'd232,8'd14} : s = 437;
	{8'd232,8'd15} : s = 501;
	{8'd232,8'd16} : s = 316;
	{8'd232,8'd17} : s = 435;
	{8'd232,8'd18} : s = 430;
	{8'd232,8'd19} : s = 499;
	{8'd232,8'd20} : s = 429;
	{8'd232,8'd21} : s = 494;
	{8'd232,8'd22} : s = 493;
	{8'd232,8'd23} : s = 510;
	{8'd232,8'd24} : s = 1;
	{8'd232,8'd25} : s = 18;
	{8'd232,8'd26} : s = 17;
	{8'd232,8'd27} : s = 82;
	{8'd232,8'd28} : s = 12;
	{8'd232,8'd29} : s = 81;
	{8'd232,8'd30} : s = 76;
	{8'd232,8'd31} : s = 195;
	{8'd232,8'd32} : s = 10;
	{8'd232,8'd33} : s = 74;
	{8'd232,8'd34} : s = 73;
	{8'd232,8'd35} : s = 184;
	{8'd232,8'd36} : s = 70;
	{8'd232,8'd37} : s = 180;
	{8'd232,8'd38} : s = 178;
	{8'd232,8'd39} : s = 314;
	{8'd232,8'd40} : s = 9;
	{8'd232,8'd41} : s = 69;
	{8'd232,8'd42} : s = 67;
	{8'd232,8'd43} : s = 177;
	{8'd232,8'd44} : s = 56;
	{8'd232,8'd45} : s = 172;
	{8'd232,8'd46} : s = 170;
	{8'd232,8'd47} : s = 313;
	{8'd232,8'd48} : s = 52;
	{8'd232,8'd49} : s = 169;
	{8'd232,8'd50} : s = 166;
	{8'd232,8'd51} : s = 310;
	{8'd232,8'd52} : s = 165;
	{8'd232,8'd53} : s = 309;
	{8'd232,8'd54} : s = 307;
	{8'd232,8'd55} : s = 427;
	{8'd232,8'd56} : s = 6;
	{8'd232,8'd57} : s = 50;
	{8'd232,8'd58} : s = 49;
	{8'd232,8'd59} : s = 163;
	{8'd232,8'd60} : s = 44;
	{8'd232,8'd61} : s = 156;
	{8'd232,8'd62} : s = 154;
	{8'd232,8'd63} : s = 302;
	{8'd232,8'd64} : s = 42;
	{8'd232,8'd65} : s = 153;
	{8'd232,8'd66} : s = 150;
	{8'd232,8'd67} : s = 301;
	{8'd232,8'd68} : s = 149;
	{8'd232,8'd69} : s = 299;
	{8'd232,8'd70} : s = 295;
	{8'd232,8'd71} : s = 423;
	{8'd232,8'd72} : s = 41;
	{8'd232,8'd73} : s = 147;
	{8'd232,8'd74} : s = 142;
	{8'd232,8'd75} : s = 286;
	{8'd232,8'd76} : s = 141;
	{8'd232,8'd77} : s = 285;
	{8'd232,8'd78} : s = 283;
	{8'd232,8'd79} : s = 414;
	{8'd232,8'd80} : s = 139;
	{8'd232,8'd81} : s = 279;
	{8'd232,8'd82} : s = 271;
	{8'd232,8'd83} : s = 413;
	{8'd232,8'd84} : s = 248;
	{8'd232,8'd85} : s = 411;
	{8'd232,8'd86} : s = 407;
	{8'd232,8'd87} : s = 491;
	{8'd232,8'd88} : s = 5;
	{8'd232,8'd89} : s = 38;
	{8'd232,8'd90} : s = 37;
	{8'd232,8'd91} : s = 135;
	{8'd232,8'd92} : s = 35;
	{8'd232,8'd93} : s = 120;
	{8'd232,8'd94} : s = 116;
	{8'd232,8'd95} : s = 244;
	{8'd232,8'd96} : s = 28;
	{8'd232,8'd97} : s = 114;
	{8'd232,8'd98} : s = 113;
	{8'd232,8'd99} : s = 242;
	{8'd232,8'd100} : s = 108;
	{8'd232,8'd101} : s = 241;
	{8'd232,8'd102} : s = 236;
	{8'd232,8'd103} : s = 399;
	{8'd232,8'd104} : s = 26;
	{8'd232,8'd105} : s = 106;
	{8'd232,8'd106} : s = 105;
	{8'd232,8'd107} : s = 234;
	{8'd232,8'd108} : s = 102;
	{8'd232,8'd109} : s = 233;
	{8'd232,8'd110} : s = 230;
	{8'd232,8'd111} : s = 380;
	{8'd232,8'd112} : s = 101;
	{8'd232,8'd113} : s = 229;
	{8'd232,8'd114} : s = 227;
	{8'd232,8'd115} : s = 378;
	{8'd232,8'd116} : s = 220;
	{8'd232,8'd117} : s = 377;
	{8'd232,8'd118} : s = 374;
	{8'd232,8'd119} : s = 487;
	{8'd232,8'd120} : s = 25;
	{8'd232,8'd121} : s = 99;
	{8'd232,8'd122} : s = 92;
	{8'd232,8'd123} : s = 218;
	{8'd232,8'd124} : s = 90;
	{8'd232,8'd125} : s = 217;
	{8'd232,8'd126} : s = 214;
	{8'd232,8'd127} : s = 373;
	{8'd232,8'd128} : s = 89;
	{8'd232,8'd129} : s = 213;
	{8'd232,8'd130} : s = 211;
	{8'd232,8'd131} : s = 371;
	{8'd232,8'd132} : s = 206;
	{8'd232,8'd133} : s = 366;
	{8'd232,8'd134} : s = 365;
	{8'd232,8'd135} : s = 478;
	{8'd232,8'd136} : s = 86;
	{8'd232,8'd137} : s = 205;
	{8'd232,8'd138} : s = 203;
	{8'd232,8'd139} : s = 363;
	{8'd232,8'd140} : s = 199;
	{8'd232,8'd141} : s = 359;
	{8'd232,8'd142} : s = 350;
	{8'd232,8'd143} : s = 477;
	{8'd232,8'd144} : s = 188;
	{8'd232,8'd145} : s = 349;
	{8'd232,8'd146} : s = 347;
	{8'd232,8'd147} : s = 475;
	{8'd232,8'd148} : s = 343;
	{8'd232,8'd149} : s = 471;
	{8'd232,8'd150} : s = 463;
	{8'd232,8'd151} : s = 509;
	{8'd232,8'd152} : s = 3;
	{8'd232,8'd153} : s = 22;
	{8'd232,8'd154} : s = 21;
	{8'd232,8'd155} : s = 85;
	{8'd232,8'd156} : s = 19;
	{8'd232,8'd157} : s = 83;
	{8'd232,8'd158} : s = 78;
	{8'd232,8'd159} : s = 186;
	{8'd232,8'd160} : s = 14;
	{8'd232,8'd161} : s = 77;
	{8'd232,8'd162} : s = 75;
	{8'd232,8'd163} : s = 185;
	{8'd232,8'd164} : s = 71;
	{8'd232,8'd165} : s = 182;
	{8'd232,8'd166} : s = 181;
	{8'd232,8'd167} : s = 335;
	{8'd232,8'd168} : s = 13;
	{8'd232,8'd169} : s = 60;
	{8'd232,8'd170} : s = 58;
	{8'd232,8'd171} : s = 179;
	{8'd232,8'd172} : s = 57;
	{8'd232,8'd173} : s = 174;
	{8'd232,8'd174} : s = 173;
	{8'd232,8'd175} : s = 318;
	{8'd232,8'd176} : s = 54;
	{8'd232,8'd177} : s = 171;
	{8'd232,8'd178} : s = 167;
	{8'd232,8'd179} : s = 317;
	{8'd232,8'd180} : s = 158;
	{8'd232,8'd181} : s = 315;
	{8'd232,8'd182} : s = 311;
	{8'd232,8'd183} : s = 446;
	{8'd232,8'd184} : s = 11;
	{8'd232,8'd185} : s = 53;
	{8'd232,8'd186} : s = 51;
	{8'd232,8'd187} : s = 157;
	{8'd232,8'd188} : s = 46;
	{8'd232,8'd189} : s = 155;
	{8'd232,8'd190} : s = 151;
	{8'd232,8'd191} : s = 303;
	{8'd232,8'd192} : s = 45;
	{8'd232,8'd193} : s = 143;
	{8'd232,8'd194} : s = 124;
	{8'd232,8'd195} : s = 287;
	{8'd232,8'd196} : s = 122;
	{8'd232,8'd197} : s = 252;
	{8'd232,8'd198} : s = 250;
	{8'd232,8'd199} : s = 445;
	{8'd232,8'd200} : s = 43;
	{8'd232,8'd201} : s = 121;
	{8'd232,8'd202} : s = 118;
	{8'd232,8'd203} : s = 249;
	{8'd232,8'd204} : s = 117;
	{8'd232,8'd205} : s = 246;
	{8'd232,8'd206} : s = 245;
	{8'd232,8'd207} : s = 443;
	{8'd232,8'd208} : s = 115;
	{8'd232,8'd209} : s = 243;
	{8'd232,8'd210} : s = 238;
	{8'd232,8'd211} : s = 439;
	{8'd232,8'd212} : s = 237;
	{8'd232,8'd213} : s = 431;
	{8'd232,8'd214} : s = 415;
	{8'd232,8'd215} : s = 507;
	{8'd232,8'd216} : s = 7;
	{8'd232,8'd217} : s = 39;
	{8'd232,8'd218} : s = 30;
	{8'd232,8'd219} : s = 110;
	{8'd232,8'd220} : s = 29;
	{8'd232,8'd221} : s = 109;
	{8'd232,8'd222} : s = 107;
	{8'd232,8'd223} : s = 235;
	{8'd232,8'd224} : s = 27;
	{8'd232,8'd225} : s = 103;
	{8'd232,8'd226} : s = 94;
	{8'd232,8'd227} : s = 231;
	{8'd232,8'd228} : s = 93;
	{8'd232,8'd229} : s = 222;
	{8'd232,8'd230} : s = 221;
	{8'd232,8'd231} : s = 382;
	{8'd232,8'd232} : s = 23;
	{8'd232,8'd233} : s = 91;
	{8'd232,8'd234} : s = 87;
	{8'd232,8'd235} : s = 219;
	{8'd232,8'd236} : s = 79;
	{8'd232,8'd237} : s = 215;
	{8'd232,8'd238} : s = 207;
	{8'd232,8'd239} : s = 381;
	{8'd232,8'd240} : s = 62;
	{8'd232,8'd241} : s = 190;
	{8'd232,8'd242} : s = 189;
	{8'd232,8'd243} : s = 379;
	{8'd232,8'd244} : s = 187;
	{8'd232,8'd245} : s = 375;
	{8'd232,8'd246} : s = 367;
	{8'd232,8'd247} : s = 503;
	{8'd232,8'd248} : s = 15;
	{8'd232,8'd249} : s = 61;
	{8'd232,8'd250} : s = 59;
	{8'd232,8'd251} : s = 183;
	{8'd232,8'd252} : s = 55;
	{8'd232,8'd253} : s = 175;
	{8'd232,8'd254} : s = 159;
	{8'd232,8'd255} : s = 351;
	{8'd233,8'd0} : s = 341;
	{8'd233,8'd1} : s = 339;
	{8'd233,8'd2} : s = 455;
	{8'd233,8'd3} : s = 334;
	{8'd233,8'd4} : s = 444;
	{8'd233,8'd5} : s = 442;
	{8'd233,8'd6} : s = 502;
	{8'd233,8'd7} : s = 197;
	{8'd233,8'd8} : s = 333;
	{8'd233,8'd9} : s = 331;
	{8'd233,8'd10} : s = 441;
	{8'd233,8'd11} : s = 327;
	{8'd233,8'd12} : s = 438;
	{8'd233,8'd13} : s = 437;
	{8'd233,8'd14} : s = 501;
	{8'd233,8'd15} : s = 316;
	{8'd233,8'd16} : s = 435;
	{8'd233,8'd17} : s = 430;
	{8'd233,8'd18} : s = 499;
	{8'd233,8'd19} : s = 429;
	{8'd233,8'd20} : s = 494;
	{8'd233,8'd21} : s = 493;
	{8'd233,8'd22} : s = 510;
	{8'd233,8'd23} : s = 1;
	{8'd233,8'd24} : s = 18;
	{8'd233,8'd25} : s = 17;
	{8'd233,8'd26} : s = 82;
	{8'd233,8'd27} : s = 12;
	{8'd233,8'd28} : s = 81;
	{8'd233,8'd29} : s = 76;
	{8'd233,8'd30} : s = 195;
	{8'd233,8'd31} : s = 10;
	{8'd233,8'd32} : s = 74;
	{8'd233,8'd33} : s = 73;
	{8'd233,8'd34} : s = 184;
	{8'd233,8'd35} : s = 70;
	{8'd233,8'd36} : s = 180;
	{8'd233,8'd37} : s = 178;
	{8'd233,8'd38} : s = 314;
	{8'd233,8'd39} : s = 9;
	{8'd233,8'd40} : s = 69;
	{8'd233,8'd41} : s = 67;
	{8'd233,8'd42} : s = 177;
	{8'd233,8'd43} : s = 56;
	{8'd233,8'd44} : s = 172;
	{8'd233,8'd45} : s = 170;
	{8'd233,8'd46} : s = 313;
	{8'd233,8'd47} : s = 52;
	{8'd233,8'd48} : s = 169;
	{8'd233,8'd49} : s = 166;
	{8'd233,8'd50} : s = 310;
	{8'd233,8'd51} : s = 165;
	{8'd233,8'd52} : s = 309;
	{8'd233,8'd53} : s = 307;
	{8'd233,8'd54} : s = 427;
	{8'd233,8'd55} : s = 6;
	{8'd233,8'd56} : s = 50;
	{8'd233,8'd57} : s = 49;
	{8'd233,8'd58} : s = 163;
	{8'd233,8'd59} : s = 44;
	{8'd233,8'd60} : s = 156;
	{8'd233,8'd61} : s = 154;
	{8'd233,8'd62} : s = 302;
	{8'd233,8'd63} : s = 42;
	{8'd233,8'd64} : s = 153;
	{8'd233,8'd65} : s = 150;
	{8'd233,8'd66} : s = 301;
	{8'd233,8'd67} : s = 149;
	{8'd233,8'd68} : s = 299;
	{8'd233,8'd69} : s = 295;
	{8'd233,8'd70} : s = 423;
	{8'd233,8'd71} : s = 41;
	{8'd233,8'd72} : s = 147;
	{8'd233,8'd73} : s = 142;
	{8'd233,8'd74} : s = 286;
	{8'd233,8'd75} : s = 141;
	{8'd233,8'd76} : s = 285;
	{8'd233,8'd77} : s = 283;
	{8'd233,8'd78} : s = 414;
	{8'd233,8'd79} : s = 139;
	{8'd233,8'd80} : s = 279;
	{8'd233,8'd81} : s = 271;
	{8'd233,8'd82} : s = 413;
	{8'd233,8'd83} : s = 248;
	{8'd233,8'd84} : s = 411;
	{8'd233,8'd85} : s = 407;
	{8'd233,8'd86} : s = 491;
	{8'd233,8'd87} : s = 5;
	{8'd233,8'd88} : s = 38;
	{8'd233,8'd89} : s = 37;
	{8'd233,8'd90} : s = 135;
	{8'd233,8'd91} : s = 35;
	{8'd233,8'd92} : s = 120;
	{8'd233,8'd93} : s = 116;
	{8'd233,8'd94} : s = 244;
	{8'd233,8'd95} : s = 28;
	{8'd233,8'd96} : s = 114;
	{8'd233,8'd97} : s = 113;
	{8'd233,8'd98} : s = 242;
	{8'd233,8'd99} : s = 108;
	{8'd233,8'd100} : s = 241;
	{8'd233,8'd101} : s = 236;
	{8'd233,8'd102} : s = 399;
	{8'd233,8'd103} : s = 26;
	{8'd233,8'd104} : s = 106;
	{8'd233,8'd105} : s = 105;
	{8'd233,8'd106} : s = 234;
	{8'd233,8'd107} : s = 102;
	{8'd233,8'd108} : s = 233;
	{8'd233,8'd109} : s = 230;
	{8'd233,8'd110} : s = 380;
	{8'd233,8'd111} : s = 101;
	{8'd233,8'd112} : s = 229;
	{8'd233,8'd113} : s = 227;
	{8'd233,8'd114} : s = 378;
	{8'd233,8'd115} : s = 220;
	{8'd233,8'd116} : s = 377;
	{8'd233,8'd117} : s = 374;
	{8'd233,8'd118} : s = 487;
	{8'd233,8'd119} : s = 25;
	{8'd233,8'd120} : s = 99;
	{8'd233,8'd121} : s = 92;
	{8'd233,8'd122} : s = 218;
	{8'd233,8'd123} : s = 90;
	{8'd233,8'd124} : s = 217;
	{8'd233,8'd125} : s = 214;
	{8'd233,8'd126} : s = 373;
	{8'd233,8'd127} : s = 89;
	{8'd233,8'd128} : s = 213;
	{8'd233,8'd129} : s = 211;
	{8'd233,8'd130} : s = 371;
	{8'd233,8'd131} : s = 206;
	{8'd233,8'd132} : s = 366;
	{8'd233,8'd133} : s = 365;
	{8'd233,8'd134} : s = 478;
	{8'd233,8'd135} : s = 86;
	{8'd233,8'd136} : s = 205;
	{8'd233,8'd137} : s = 203;
	{8'd233,8'd138} : s = 363;
	{8'd233,8'd139} : s = 199;
	{8'd233,8'd140} : s = 359;
	{8'd233,8'd141} : s = 350;
	{8'd233,8'd142} : s = 477;
	{8'd233,8'd143} : s = 188;
	{8'd233,8'd144} : s = 349;
	{8'd233,8'd145} : s = 347;
	{8'd233,8'd146} : s = 475;
	{8'd233,8'd147} : s = 343;
	{8'd233,8'd148} : s = 471;
	{8'd233,8'd149} : s = 463;
	{8'd233,8'd150} : s = 509;
	{8'd233,8'd151} : s = 3;
	{8'd233,8'd152} : s = 22;
	{8'd233,8'd153} : s = 21;
	{8'd233,8'd154} : s = 85;
	{8'd233,8'd155} : s = 19;
	{8'd233,8'd156} : s = 83;
	{8'd233,8'd157} : s = 78;
	{8'd233,8'd158} : s = 186;
	{8'd233,8'd159} : s = 14;
	{8'd233,8'd160} : s = 77;
	{8'd233,8'd161} : s = 75;
	{8'd233,8'd162} : s = 185;
	{8'd233,8'd163} : s = 71;
	{8'd233,8'd164} : s = 182;
	{8'd233,8'd165} : s = 181;
	{8'd233,8'd166} : s = 335;
	{8'd233,8'd167} : s = 13;
	{8'd233,8'd168} : s = 60;
	{8'd233,8'd169} : s = 58;
	{8'd233,8'd170} : s = 179;
	{8'd233,8'd171} : s = 57;
	{8'd233,8'd172} : s = 174;
	{8'd233,8'd173} : s = 173;
	{8'd233,8'd174} : s = 318;
	{8'd233,8'd175} : s = 54;
	{8'd233,8'd176} : s = 171;
	{8'd233,8'd177} : s = 167;
	{8'd233,8'd178} : s = 317;
	{8'd233,8'd179} : s = 158;
	{8'd233,8'd180} : s = 315;
	{8'd233,8'd181} : s = 311;
	{8'd233,8'd182} : s = 446;
	{8'd233,8'd183} : s = 11;
	{8'd233,8'd184} : s = 53;
	{8'd233,8'd185} : s = 51;
	{8'd233,8'd186} : s = 157;
	{8'd233,8'd187} : s = 46;
	{8'd233,8'd188} : s = 155;
	{8'd233,8'd189} : s = 151;
	{8'd233,8'd190} : s = 303;
	{8'd233,8'd191} : s = 45;
	{8'd233,8'd192} : s = 143;
	{8'd233,8'd193} : s = 124;
	{8'd233,8'd194} : s = 287;
	{8'd233,8'd195} : s = 122;
	{8'd233,8'd196} : s = 252;
	{8'd233,8'd197} : s = 250;
	{8'd233,8'd198} : s = 445;
	{8'd233,8'd199} : s = 43;
	{8'd233,8'd200} : s = 121;
	{8'd233,8'd201} : s = 118;
	{8'd233,8'd202} : s = 249;
	{8'd233,8'd203} : s = 117;
	{8'd233,8'd204} : s = 246;
	{8'd233,8'd205} : s = 245;
	{8'd233,8'd206} : s = 443;
	{8'd233,8'd207} : s = 115;
	{8'd233,8'd208} : s = 243;
	{8'd233,8'd209} : s = 238;
	{8'd233,8'd210} : s = 439;
	{8'd233,8'd211} : s = 237;
	{8'd233,8'd212} : s = 431;
	{8'd233,8'd213} : s = 415;
	{8'd233,8'd214} : s = 507;
	{8'd233,8'd215} : s = 7;
	{8'd233,8'd216} : s = 39;
	{8'd233,8'd217} : s = 30;
	{8'd233,8'd218} : s = 110;
	{8'd233,8'd219} : s = 29;
	{8'd233,8'd220} : s = 109;
	{8'd233,8'd221} : s = 107;
	{8'd233,8'd222} : s = 235;
	{8'd233,8'd223} : s = 27;
	{8'd233,8'd224} : s = 103;
	{8'd233,8'd225} : s = 94;
	{8'd233,8'd226} : s = 231;
	{8'd233,8'd227} : s = 93;
	{8'd233,8'd228} : s = 222;
	{8'd233,8'd229} : s = 221;
	{8'd233,8'd230} : s = 382;
	{8'd233,8'd231} : s = 23;
	{8'd233,8'd232} : s = 91;
	{8'd233,8'd233} : s = 87;
	{8'd233,8'd234} : s = 219;
	{8'd233,8'd235} : s = 79;
	{8'd233,8'd236} : s = 215;
	{8'd233,8'd237} : s = 207;
	{8'd233,8'd238} : s = 381;
	{8'd233,8'd239} : s = 62;
	{8'd233,8'd240} : s = 190;
	{8'd233,8'd241} : s = 189;
	{8'd233,8'd242} : s = 379;
	{8'd233,8'd243} : s = 187;
	{8'd233,8'd244} : s = 375;
	{8'd233,8'd245} : s = 367;
	{8'd233,8'd246} : s = 503;
	{8'd233,8'd247} : s = 15;
	{8'd233,8'd248} : s = 61;
	{8'd233,8'd249} : s = 59;
	{8'd233,8'd250} : s = 183;
	{8'd233,8'd251} : s = 55;
	{8'd233,8'd252} : s = 175;
	{8'd233,8'd253} : s = 159;
	{8'd233,8'd254} : s = 351;
	{8'd233,8'd255} : s = 47;
	{8'd234,8'd0} : s = 339;
	{8'd234,8'd1} : s = 455;
	{8'd234,8'd2} : s = 334;
	{8'd234,8'd3} : s = 444;
	{8'd234,8'd4} : s = 442;
	{8'd234,8'd5} : s = 502;
	{8'd234,8'd6} : s = 197;
	{8'd234,8'd7} : s = 333;
	{8'd234,8'd8} : s = 331;
	{8'd234,8'd9} : s = 441;
	{8'd234,8'd10} : s = 327;
	{8'd234,8'd11} : s = 438;
	{8'd234,8'd12} : s = 437;
	{8'd234,8'd13} : s = 501;
	{8'd234,8'd14} : s = 316;
	{8'd234,8'd15} : s = 435;
	{8'd234,8'd16} : s = 430;
	{8'd234,8'd17} : s = 499;
	{8'd234,8'd18} : s = 429;
	{8'd234,8'd19} : s = 494;
	{8'd234,8'd20} : s = 493;
	{8'd234,8'd21} : s = 510;
	{8'd234,8'd22} : s = 1;
	{8'd234,8'd23} : s = 18;
	{8'd234,8'd24} : s = 17;
	{8'd234,8'd25} : s = 82;
	{8'd234,8'd26} : s = 12;
	{8'd234,8'd27} : s = 81;
	{8'd234,8'd28} : s = 76;
	{8'd234,8'd29} : s = 195;
	{8'd234,8'd30} : s = 10;
	{8'd234,8'd31} : s = 74;
	{8'd234,8'd32} : s = 73;
	{8'd234,8'd33} : s = 184;
	{8'd234,8'd34} : s = 70;
	{8'd234,8'd35} : s = 180;
	{8'd234,8'd36} : s = 178;
	{8'd234,8'd37} : s = 314;
	{8'd234,8'd38} : s = 9;
	{8'd234,8'd39} : s = 69;
	{8'd234,8'd40} : s = 67;
	{8'd234,8'd41} : s = 177;
	{8'd234,8'd42} : s = 56;
	{8'd234,8'd43} : s = 172;
	{8'd234,8'd44} : s = 170;
	{8'd234,8'd45} : s = 313;
	{8'd234,8'd46} : s = 52;
	{8'd234,8'd47} : s = 169;
	{8'd234,8'd48} : s = 166;
	{8'd234,8'd49} : s = 310;
	{8'd234,8'd50} : s = 165;
	{8'd234,8'd51} : s = 309;
	{8'd234,8'd52} : s = 307;
	{8'd234,8'd53} : s = 427;
	{8'd234,8'd54} : s = 6;
	{8'd234,8'd55} : s = 50;
	{8'd234,8'd56} : s = 49;
	{8'd234,8'd57} : s = 163;
	{8'd234,8'd58} : s = 44;
	{8'd234,8'd59} : s = 156;
	{8'd234,8'd60} : s = 154;
	{8'd234,8'd61} : s = 302;
	{8'd234,8'd62} : s = 42;
	{8'd234,8'd63} : s = 153;
	{8'd234,8'd64} : s = 150;
	{8'd234,8'd65} : s = 301;
	{8'd234,8'd66} : s = 149;
	{8'd234,8'd67} : s = 299;
	{8'd234,8'd68} : s = 295;
	{8'd234,8'd69} : s = 423;
	{8'd234,8'd70} : s = 41;
	{8'd234,8'd71} : s = 147;
	{8'd234,8'd72} : s = 142;
	{8'd234,8'd73} : s = 286;
	{8'd234,8'd74} : s = 141;
	{8'd234,8'd75} : s = 285;
	{8'd234,8'd76} : s = 283;
	{8'd234,8'd77} : s = 414;
	{8'd234,8'd78} : s = 139;
	{8'd234,8'd79} : s = 279;
	{8'd234,8'd80} : s = 271;
	{8'd234,8'd81} : s = 413;
	{8'd234,8'd82} : s = 248;
	{8'd234,8'd83} : s = 411;
	{8'd234,8'd84} : s = 407;
	{8'd234,8'd85} : s = 491;
	{8'd234,8'd86} : s = 5;
	{8'd234,8'd87} : s = 38;
	{8'd234,8'd88} : s = 37;
	{8'd234,8'd89} : s = 135;
	{8'd234,8'd90} : s = 35;
	{8'd234,8'd91} : s = 120;
	{8'd234,8'd92} : s = 116;
	{8'd234,8'd93} : s = 244;
	{8'd234,8'd94} : s = 28;
	{8'd234,8'd95} : s = 114;
	{8'd234,8'd96} : s = 113;
	{8'd234,8'd97} : s = 242;
	{8'd234,8'd98} : s = 108;
	{8'd234,8'd99} : s = 241;
	{8'd234,8'd100} : s = 236;
	{8'd234,8'd101} : s = 399;
	{8'd234,8'd102} : s = 26;
	{8'd234,8'd103} : s = 106;
	{8'd234,8'd104} : s = 105;
	{8'd234,8'd105} : s = 234;
	{8'd234,8'd106} : s = 102;
	{8'd234,8'd107} : s = 233;
	{8'd234,8'd108} : s = 230;
	{8'd234,8'd109} : s = 380;
	{8'd234,8'd110} : s = 101;
	{8'd234,8'd111} : s = 229;
	{8'd234,8'd112} : s = 227;
	{8'd234,8'd113} : s = 378;
	{8'd234,8'd114} : s = 220;
	{8'd234,8'd115} : s = 377;
	{8'd234,8'd116} : s = 374;
	{8'd234,8'd117} : s = 487;
	{8'd234,8'd118} : s = 25;
	{8'd234,8'd119} : s = 99;
	{8'd234,8'd120} : s = 92;
	{8'd234,8'd121} : s = 218;
	{8'd234,8'd122} : s = 90;
	{8'd234,8'd123} : s = 217;
	{8'd234,8'd124} : s = 214;
	{8'd234,8'd125} : s = 373;
	{8'd234,8'd126} : s = 89;
	{8'd234,8'd127} : s = 213;
	{8'd234,8'd128} : s = 211;
	{8'd234,8'd129} : s = 371;
	{8'd234,8'd130} : s = 206;
	{8'd234,8'd131} : s = 366;
	{8'd234,8'd132} : s = 365;
	{8'd234,8'd133} : s = 478;
	{8'd234,8'd134} : s = 86;
	{8'd234,8'd135} : s = 205;
	{8'd234,8'd136} : s = 203;
	{8'd234,8'd137} : s = 363;
	{8'd234,8'd138} : s = 199;
	{8'd234,8'd139} : s = 359;
	{8'd234,8'd140} : s = 350;
	{8'd234,8'd141} : s = 477;
	{8'd234,8'd142} : s = 188;
	{8'd234,8'd143} : s = 349;
	{8'd234,8'd144} : s = 347;
	{8'd234,8'd145} : s = 475;
	{8'd234,8'd146} : s = 343;
	{8'd234,8'd147} : s = 471;
	{8'd234,8'd148} : s = 463;
	{8'd234,8'd149} : s = 509;
	{8'd234,8'd150} : s = 3;
	{8'd234,8'd151} : s = 22;
	{8'd234,8'd152} : s = 21;
	{8'd234,8'd153} : s = 85;
	{8'd234,8'd154} : s = 19;
	{8'd234,8'd155} : s = 83;
	{8'd234,8'd156} : s = 78;
	{8'd234,8'd157} : s = 186;
	{8'd234,8'd158} : s = 14;
	{8'd234,8'd159} : s = 77;
	{8'd234,8'd160} : s = 75;
	{8'd234,8'd161} : s = 185;
	{8'd234,8'd162} : s = 71;
	{8'd234,8'd163} : s = 182;
	{8'd234,8'd164} : s = 181;
	{8'd234,8'd165} : s = 335;
	{8'd234,8'd166} : s = 13;
	{8'd234,8'd167} : s = 60;
	{8'd234,8'd168} : s = 58;
	{8'd234,8'd169} : s = 179;
	{8'd234,8'd170} : s = 57;
	{8'd234,8'd171} : s = 174;
	{8'd234,8'd172} : s = 173;
	{8'd234,8'd173} : s = 318;
	{8'd234,8'd174} : s = 54;
	{8'd234,8'd175} : s = 171;
	{8'd234,8'd176} : s = 167;
	{8'd234,8'd177} : s = 317;
	{8'd234,8'd178} : s = 158;
	{8'd234,8'd179} : s = 315;
	{8'd234,8'd180} : s = 311;
	{8'd234,8'd181} : s = 446;
	{8'd234,8'd182} : s = 11;
	{8'd234,8'd183} : s = 53;
	{8'd234,8'd184} : s = 51;
	{8'd234,8'd185} : s = 157;
	{8'd234,8'd186} : s = 46;
	{8'd234,8'd187} : s = 155;
	{8'd234,8'd188} : s = 151;
	{8'd234,8'd189} : s = 303;
	{8'd234,8'd190} : s = 45;
	{8'd234,8'd191} : s = 143;
	{8'd234,8'd192} : s = 124;
	{8'd234,8'd193} : s = 287;
	{8'd234,8'd194} : s = 122;
	{8'd234,8'd195} : s = 252;
	{8'd234,8'd196} : s = 250;
	{8'd234,8'd197} : s = 445;
	{8'd234,8'd198} : s = 43;
	{8'd234,8'd199} : s = 121;
	{8'd234,8'd200} : s = 118;
	{8'd234,8'd201} : s = 249;
	{8'd234,8'd202} : s = 117;
	{8'd234,8'd203} : s = 246;
	{8'd234,8'd204} : s = 245;
	{8'd234,8'd205} : s = 443;
	{8'd234,8'd206} : s = 115;
	{8'd234,8'd207} : s = 243;
	{8'd234,8'd208} : s = 238;
	{8'd234,8'd209} : s = 439;
	{8'd234,8'd210} : s = 237;
	{8'd234,8'd211} : s = 431;
	{8'd234,8'd212} : s = 415;
	{8'd234,8'd213} : s = 507;
	{8'd234,8'd214} : s = 7;
	{8'd234,8'd215} : s = 39;
	{8'd234,8'd216} : s = 30;
	{8'd234,8'd217} : s = 110;
	{8'd234,8'd218} : s = 29;
	{8'd234,8'd219} : s = 109;
	{8'd234,8'd220} : s = 107;
	{8'd234,8'd221} : s = 235;
	{8'd234,8'd222} : s = 27;
	{8'd234,8'd223} : s = 103;
	{8'd234,8'd224} : s = 94;
	{8'd234,8'd225} : s = 231;
	{8'd234,8'd226} : s = 93;
	{8'd234,8'd227} : s = 222;
	{8'd234,8'd228} : s = 221;
	{8'd234,8'd229} : s = 382;
	{8'd234,8'd230} : s = 23;
	{8'd234,8'd231} : s = 91;
	{8'd234,8'd232} : s = 87;
	{8'd234,8'd233} : s = 219;
	{8'd234,8'd234} : s = 79;
	{8'd234,8'd235} : s = 215;
	{8'd234,8'd236} : s = 207;
	{8'd234,8'd237} : s = 381;
	{8'd234,8'd238} : s = 62;
	{8'd234,8'd239} : s = 190;
	{8'd234,8'd240} : s = 189;
	{8'd234,8'd241} : s = 379;
	{8'd234,8'd242} : s = 187;
	{8'd234,8'd243} : s = 375;
	{8'd234,8'd244} : s = 367;
	{8'd234,8'd245} : s = 503;
	{8'd234,8'd246} : s = 15;
	{8'd234,8'd247} : s = 61;
	{8'd234,8'd248} : s = 59;
	{8'd234,8'd249} : s = 183;
	{8'd234,8'd250} : s = 55;
	{8'd234,8'd251} : s = 175;
	{8'd234,8'd252} : s = 159;
	{8'd234,8'd253} : s = 351;
	{8'd234,8'd254} : s = 47;
	{8'd234,8'd255} : s = 126;
	{8'd235,8'd0} : s = 455;
	{8'd235,8'd1} : s = 334;
	{8'd235,8'd2} : s = 444;
	{8'd235,8'd3} : s = 442;
	{8'd235,8'd4} : s = 502;
	{8'd235,8'd5} : s = 197;
	{8'd235,8'd6} : s = 333;
	{8'd235,8'd7} : s = 331;
	{8'd235,8'd8} : s = 441;
	{8'd235,8'd9} : s = 327;
	{8'd235,8'd10} : s = 438;
	{8'd235,8'd11} : s = 437;
	{8'd235,8'd12} : s = 501;
	{8'd235,8'd13} : s = 316;
	{8'd235,8'd14} : s = 435;
	{8'd235,8'd15} : s = 430;
	{8'd235,8'd16} : s = 499;
	{8'd235,8'd17} : s = 429;
	{8'd235,8'd18} : s = 494;
	{8'd235,8'd19} : s = 493;
	{8'd235,8'd20} : s = 510;
	{8'd235,8'd21} : s = 1;
	{8'd235,8'd22} : s = 18;
	{8'd235,8'd23} : s = 17;
	{8'd235,8'd24} : s = 82;
	{8'd235,8'd25} : s = 12;
	{8'd235,8'd26} : s = 81;
	{8'd235,8'd27} : s = 76;
	{8'd235,8'd28} : s = 195;
	{8'd235,8'd29} : s = 10;
	{8'd235,8'd30} : s = 74;
	{8'd235,8'd31} : s = 73;
	{8'd235,8'd32} : s = 184;
	{8'd235,8'd33} : s = 70;
	{8'd235,8'd34} : s = 180;
	{8'd235,8'd35} : s = 178;
	{8'd235,8'd36} : s = 314;
	{8'd235,8'd37} : s = 9;
	{8'd235,8'd38} : s = 69;
	{8'd235,8'd39} : s = 67;
	{8'd235,8'd40} : s = 177;
	{8'd235,8'd41} : s = 56;
	{8'd235,8'd42} : s = 172;
	{8'd235,8'd43} : s = 170;
	{8'd235,8'd44} : s = 313;
	{8'd235,8'd45} : s = 52;
	{8'd235,8'd46} : s = 169;
	{8'd235,8'd47} : s = 166;
	{8'd235,8'd48} : s = 310;
	{8'd235,8'd49} : s = 165;
	{8'd235,8'd50} : s = 309;
	{8'd235,8'd51} : s = 307;
	{8'd235,8'd52} : s = 427;
	{8'd235,8'd53} : s = 6;
	{8'd235,8'd54} : s = 50;
	{8'd235,8'd55} : s = 49;
	{8'd235,8'd56} : s = 163;
	{8'd235,8'd57} : s = 44;
	{8'd235,8'd58} : s = 156;
	{8'd235,8'd59} : s = 154;
	{8'd235,8'd60} : s = 302;
	{8'd235,8'd61} : s = 42;
	{8'd235,8'd62} : s = 153;
	{8'd235,8'd63} : s = 150;
	{8'd235,8'd64} : s = 301;
	{8'd235,8'd65} : s = 149;
	{8'd235,8'd66} : s = 299;
	{8'd235,8'd67} : s = 295;
	{8'd235,8'd68} : s = 423;
	{8'd235,8'd69} : s = 41;
	{8'd235,8'd70} : s = 147;
	{8'd235,8'd71} : s = 142;
	{8'd235,8'd72} : s = 286;
	{8'd235,8'd73} : s = 141;
	{8'd235,8'd74} : s = 285;
	{8'd235,8'd75} : s = 283;
	{8'd235,8'd76} : s = 414;
	{8'd235,8'd77} : s = 139;
	{8'd235,8'd78} : s = 279;
	{8'd235,8'd79} : s = 271;
	{8'd235,8'd80} : s = 413;
	{8'd235,8'd81} : s = 248;
	{8'd235,8'd82} : s = 411;
	{8'd235,8'd83} : s = 407;
	{8'd235,8'd84} : s = 491;
	{8'd235,8'd85} : s = 5;
	{8'd235,8'd86} : s = 38;
	{8'd235,8'd87} : s = 37;
	{8'd235,8'd88} : s = 135;
	{8'd235,8'd89} : s = 35;
	{8'd235,8'd90} : s = 120;
	{8'd235,8'd91} : s = 116;
	{8'd235,8'd92} : s = 244;
	{8'd235,8'd93} : s = 28;
	{8'd235,8'd94} : s = 114;
	{8'd235,8'd95} : s = 113;
	{8'd235,8'd96} : s = 242;
	{8'd235,8'd97} : s = 108;
	{8'd235,8'd98} : s = 241;
	{8'd235,8'd99} : s = 236;
	{8'd235,8'd100} : s = 399;
	{8'd235,8'd101} : s = 26;
	{8'd235,8'd102} : s = 106;
	{8'd235,8'd103} : s = 105;
	{8'd235,8'd104} : s = 234;
	{8'd235,8'd105} : s = 102;
	{8'd235,8'd106} : s = 233;
	{8'd235,8'd107} : s = 230;
	{8'd235,8'd108} : s = 380;
	{8'd235,8'd109} : s = 101;
	{8'd235,8'd110} : s = 229;
	{8'd235,8'd111} : s = 227;
	{8'd235,8'd112} : s = 378;
	{8'd235,8'd113} : s = 220;
	{8'd235,8'd114} : s = 377;
	{8'd235,8'd115} : s = 374;
	{8'd235,8'd116} : s = 487;
	{8'd235,8'd117} : s = 25;
	{8'd235,8'd118} : s = 99;
	{8'd235,8'd119} : s = 92;
	{8'd235,8'd120} : s = 218;
	{8'd235,8'd121} : s = 90;
	{8'd235,8'd122} : s = 217;
	{8'd235,8'd123} : s = 214;
	{8'd235,8'd124} : s = 373;
	{8'd235,8'd125} : s = 89;
	{8'd235,8'd126} : s = 213;
	{8'd235,8'd127} : s = 211;
	{8'd235,8'd128} : s = 371;
	{8'd235,8'd129} : s = 206;
	{8'd235,8'd130} : s = 366;
	{8'd235,8'd131} : s = 365;
	{8'd235,8'd132} : s = 478;
	{8'd235,8'd133} : s = 86;
	{8'd235,8'd134} : s = 205;
	{8'd235,8'd135} : s = 203;
	{8'd235,8'd136} : s = 363;
	{8'd235,8'd137} : s = 199;
	{8'd235,8'd138} : s = 359;
	{8'd235,8'd139} : s = 350;
	{8'd235,8'd140} : s = 477;
	{8'd235,8'd141} : s = 188;
	{8'd235,8'd142} : s = 349;
	{8'd235,8'd143} : s = 347;
	{8'd235,8'd144} : s = 475;
	{8'd235,8'd145} : s = 343;
	{8'd235,8'd146} : s = 471;
	{8'd235,8'd147} : s = 463;
	{8'd235,8'd148} : s = 509;
	{8'd235,8'd149} : s = 3;
	{8'd235,8'd150} : s = 22;
	{8'd235,8'd151} : s = 21;
	{8'd235,8'd152} : s = 85;
	{8'd235,8'd153} : s = 19;
	{8'd235,8'd154} : s = 83;
	{8'd235,8'd155} : s = 78;
	{8'd235,8'd156} : s = 186;
	{8'd235,8'd157} : s = 14;
	{8'd235,8'd158} : s = 77;
	{8'd235,8'd159} : s = 75;
	{8'd235,8'd160} : s = 185;
	{8'd235,8'd161} : s = 71;
	{8'd235,8'd162} : s = 182;
	{8'd235,8'd163} : s = 181;
	{8'd235,8'd164} : s = 335;
	{8'd235,8'd165} : s = 13;
	{8'd235,8'd166} : s = 60;
	{8'd235,8'd167} : s = 58;
	{8'd235,8'd168} : s = 179;
	{8'd235,8'd169} : s = 57;
	{8'd235,8'd170} : s = 174;
	{8'd235,8'd171} : s = 173;
	{8'd235,8'd172} : s = 318;
	{8'd235,8'd173} : s = 54;
	{8'd235,8'd174} : s = 171;
	{8'd235,8'd175} : s = 167;
	{8'd235,8'd176} : s = 317;
	{8'd235,8'd177} : s = 158;
	{8'd235,8'd178} : s = 315;
	{8'd235,8'd179} : s = 311;
	{8'd235,8'd180} : s = 446;
	{8'd235,8'd181} : s = 11;
	{8'd235,8'd182} : s = 53;
	{8'd235,8'd183} : s = 51;
	{8'd235,8'd184} : s = 157;
	{8'd235,8'd185} : s = 46;
	{8'd235,8'd186} : s = 155;
	{8'd235,8'd187} : s = 151;
	{8'd235,8'd188} : s = 303;
	{8'd235,8'd189} : s = 45;
	{8'd235,8'd190} : s = 143;
	{8'd235,8'd191} : s = 124;
	{8'd235,8'd192} : s = 287;
	{8'd235,8'd193} : s = 122;
	{8'd235,8'd194} : s = 252;
	{8'd235,8'd195} : s = 250;
	{8'd235,8'd196} : s = 445;
	{8'd235,8'd197} : s = 43;
	{8'd235,8'd198} : s = 121;
	{8'd235,8'd199} : s = 118;
	{8'd235,8'd200} : s = 249;
	{8'd235,8'd201} : s = 117;
	{8'd235,8'd202} : s = 246;
	{8'd235,8'd203} : s = 245;
	{8'd235,8'd204} : s = 443;
	{8'd235,8'd205} : s = 115;
	{8'd235,8'd206} : s = 243;
	{8'd235,8'd207} : s = 238;
	{8'd235,8'd208} : s = 439;
	{8'd235,8'd209} : s = 237;
	{8'd235,8'd210} : s = 431;
	{8'd235,8'd211} : s = 415;
	{8'd235,8'd212} : s = 507;
	{8'd235,8'd213} : s = 7;
	{8'd235,8'd214} : s = 39;
	{8'd235,8'd215} : s = 30;
	{8'd235,8'd216} : s = 110;
	{8'd235,8'd217} : s = 29;
	{8'd235,8'd218} : s = 109;
	{8'd235,8'd219} : s = 107;
	{8'd235,8'd220} : s = 235;
	{8'd235,8'd221} : s = 27;
	{8'd235,8'd222} : s = 103;
	{8'd235,8'd223} : s = 94;
	{8'd235,8'd224} : s = 231;
	{8'd235,8'd225} : s = 93;
	{8'd235,8'd226} : s = 222;
	{8'd235,8'd227} : s = 221;
	{8'd235,8'd228} : s = 382;
	{8'd235,8'd229} : s = 23;
	{8'd235,8'd230} : s = 91;
	{8'd235,8'd231} : s = 87;
	{8'd235,8'd232} : s = 219;
	{8'd235,8'd233} : s = 79;
	{8'd235,8'd234} : s = 215;
	{8'd235,8'd235} : s = 207;
	{8'd235,8'd236} : s = 381;
	{8'd235,8'd237} : s = 62;
	{8'd235,8'd238} : s = 190;
	{8'd235,8'd239} : s = 189;
	{8'd235,8'd240} : s = 379;
	{8'd235,8'd241} : s = 187;
	{8'd235,8'd242} : s = 375;
	{8'd235,8'd243} : s = 367;
	{8'd235,8'd244} : s = 503;
	{8'd235,8'd245} : s = 15;
	{8'd235,8'd246} : s = 61;
	{8'd235,8'd247} : s = 59;
	{8'd235,8'd248} : s = 183;
	{8'd235,8'd249} : s = 55;
	{8'd235,8'd250} : s = 175;
	{8'd235,8'd251} : s = 159;
	{8'd235,8'd252} : s = 351;
	{8'd235,8'd253} : s = 47;
	{8'd235,8'd254} : s = 126;
	{8'd235,8'd255} : s = 125;
	{8'd236,8'd0} : s = 334;
	{8'd236,8'd1} : s = 444;
	{8'd236,8'd2} : s = 442;
	{8'd236,8'd3} : s = 502;
	{8'd236,8'd4} : s = 197;
	{8'd236,8'd5} : s = 333;
	{8'd236,8'd6} : s = 331;
	{8'd236,8'd7} : s = 441;
	{8'd236,8'd8} : s = 327;
	{8'd236,8'd9} : s = 438;
	{8'd236,8'd10} : s = 437;
	{8'd236,8'd11} : s = 501;
	{8'd236,8'd12} : s = 316;
	{8'd236,8'd13} : s = 435;
	{8'd236,8'd14} : s = 430;
	{8'd236,8'd15} : s = 499;
	{8'd236,8'd16} : s = 429;
	{8'd236,8'd17} : s = 494;
	{8'd236,8'd18} : s = 493;
	{8'd236,8'd19} : s = 510;
	{8'd236,8'd20} : s = 1;
	{8'd236,8'd21} : s = 18;
	{8'd236,8'd22} : s = 17;
	{8'd236,8'd23} : s = 82;
	{8'd236,8'd24} : s = 12;
	{8'd236,8'd25} : s = 81;
	{8'd236,8'd26} : s = 76;
	{8'd236,8'd27} : s = 195;
	{8'd236,8'd28} : s = 10;
	{8'd236,8'd29} : s = 74;
	{8'd236,8'd30} : s = 73;
	{8'd236,8'd31} : s = 184;
	{8'd236,8'd32} : s = 70;
	{8'd236,8'd33} : s = 180;
	{8'd236,8'd34} : s = 178;
	{8'd236,8'd35} : s = 314;
	{8'd236,8'd36} : s = 9;
	{8'd236,8'd37} : s = 69;
	{8'd236,8'd38} : s = 67;
	{8'd236,8'd39} : s = 177;
	{8'd236,8'd40} : s = 56;
	{8'd236,8'd41} : s = 172;
	{8'd236,8'd42} : s = 170;
	{8'd236,8'd43} : s = 313;
	{8'd236,8'd44} : s = 52;
	{8'd236,8'd45} : s = 169;
	{8'd236,8'd46} : s = 166;
	{8'd236,8'd47} : s = 310;
	{8'd236,8'd48} : s = 165;
	{8'd236,8'd49} : s = 309;
	{8'd236,8'd50} : s = 307;
	{8'd236,8'd51} : s = 427;
	{8'd236,8'd52} : s = 6;
	{8'd236,8'd53} : s = 50;
	{8'd236,8'd54} : s = 49;
	{8'd236,8'd55} : s = 163;
	{8'd236,8'd56} : s = 44;
	{8'd236,8'd57} : s = 156;
	{8'd236,8'd58} : s = 154;
	{8'd236,8'd59} : s = 302;
	{8'd236,8'd60} : s = 42;
	{8'd236,8'd61} : s = 153;
	{8'd236,8'd62} : s = 150;
	{8'd236,8'd63} : s = 301;
	{8'd236,8'd64} : s = 149;
	{8'd236,8'd65} : s = 299;
	{8'd236,8'd66} : s = 295;
	{8'd236,8'd67} : s = 423;
	{8'd236,8'd68} : s = 41;
	{8'd236,8'd69} : s = 147;
	{8'd236,8'd70} : s = 142;
	{8'd236,8'd71} : s = 286;
	{8'd236,8'd72} : s = 141;
	{8'd236,8'd73} : s = 285;
	{8'd236,8'd74} : s = 283;
	{8'd236,8'd75} : s = 414;
	{8'd236,8'd76} : s = 139;
	{8'd236,8'd77} : s = 279;
	{8'd236,8'd78} : s = 271;
	{8'd236,8'd79} : s = 413;
	{8'd236,8'd80} : s = 248;
	{8'd236,8'd81} : s = 411;
	{8'd236,8'd82} : s = 407;
	{8'd236,8'd83} : s = 491;
	{8'd236,8'd84} : s = 5;
	{8'd236,8'd85} : s = 38;
	{8'd236,8'd86} : s = 37;
	{8'd236,8'd87} : s = 135;
	{8'd236,8'd88} : s = 35;
	{8'd236,8'd89} : s = 120;
	{8'd236,8'd90} : s = 116;
	{8'd236,8'd91} : s = 244;
	{8'd236,8'd92} : s = 28;
	{8'd236,8'd93} : s = 114;
	{8'd236,8'd94} : s = 113;
	{8'd236,8'd95} : s = 242;
	{8'd236,8'd96} : s = 108;
	{8'd236,8'd97} : s = 241;
	{8'd236,8'd98} : s = 236;
	{8'd236,8'd99} : s = 399;
	{8'd236,8'd100} : s = 26;
	{8'd236,8'd101} : s = 106;
	{8'd236,8'd102} : s = 105;
	{8'd236,8'd103} : s = 234;
	{8'd236,8'd104} : s = 102;
	{8'd236,8'd105} : s = 233;
	{8'd236,8'd106} : s = 230;
	{8'd236,8'd107} : s = 380;
	{8'd236,8'd108} : s = 101;
	{8'd236,8'd109} : s = 229;
	{8'd236,8'd110} : s = 227;
	{8'd236,8'd111} : s = 378;
	{8'd236,8'd112} : s = 220;
	{8'd236,8'd113} : s = 377;
	{8'd236,8'd114} : s = 374;
	{8'd236,8'd115} : s = 487;
	{8'd236,8'd116} : s = 25;
	{8'd236,8'd117} : s = 99;
	{8'd236,8'd118} : s = 92;
	{8'd236,8'd119} : s = 218;
	{8'd236,8'd120} : s = 90;
	{8'd236,8'd121} : s = 217;
	{8'd236,8'd122} : s = 214;
	{8'd236,8'd123} : s = 373;
	{8'd236,8'd124} : s = 89;
	{8'd236,8'd125} : s = 213;
	{8'd236,8'd126} : s = 211;
	{8'd236,8'd127} : s = 371;
	{8'd236,8'd128} : s = 206;
	{8'd236,8'd129} : s = 366;
	{8'd236,8'd130} : s = 365;
	{8'd236,8'd131} : s = 478;
	{8'd236,8'd132} : s = 86;
	{8'd236,8'd133} : s = 205;
	{8'd236,8'd134} : s = 203;
	{8'd236,8'd135} : s = 363;
	{8'd236,8'd136} : s = 199;
	{8'd236,8'd137} : s = 359;
	{8'd236,8'd138} : s = 350;
	{8'd236,8'd139} : s = 477;
	{8'd236,8'd140} : s = 188;
	{8'd236,8'd141} : s = 349;
	{8'd236,8'd142} : s = 347;
	{8'd236,8'd143} : s = 475;
	{8'd236,8'd144} : s = 343;
	{8'd236,8'd145} : s = 471;
	{8'd236,8'd146} : s = 463;
	{8'd236,8'd147} : s = 509;
	{8'd236,8'd148} : s = 3;
	{8'd236,8'd149} : s = 22;
	{8'd236,8'd150} : s = 21;
	{8'd236,8'd151} : s = 85;
	{8'd236,8'd152} : s = 19;
	{8'd236,8'd153} : s = 83;
	{8'd236,8'd154} : s = 78;
	{8'd236,8'd155} : s = 186;
	{8'd236,8'd156} : s = 14;
	{8'd236,8'd157} : s = 77;
	{8'd236,8'd158} : s = 75;
	{8'd236,8'd159} : s = 185;
	{8'd236,8'd160} : s = 71;
	{8'd236,8'd161} : s = 182;
	{8'd236,8'd162} : s = 181;
	{8'd236,8'd163} : s = 335;
	{8'd236,8'd164} : s = 13;
	{8'd236,8'd165} : s = 60;
	{8'd236,8'd166} : s = 58;
	{8'd236,8'd167} : s = 179;
	{8'd236,8'd168} : s = 57;
	{8'd236,8'd169} : s = 174;
	{8'd236,8'd170} : s = 173;
	{8'd236,8'd171} : s = 318;
	{8'd236,8'd172} : s = 54;
	{8'd236,8'd173} : s = 171;
	{8'd236,8'd174} : s = 167;
	{8'd236,8'd175} : s = 317;
	{8'd236,8'd176} : s = 158;
	{8'd236,8'd177} : s = 315;
	{8'd236,8'd178} : s = 311;
	{8'd236,8'd179} : s = 446;
	{8'd236,8'd180} : s = 11;
	{8'd236,8'd181} : s = 53;
	{8'd236,8'd182} : s = 51;
	{8'd236,8'd183} : s = 157;
	{8'd236,8'd184} : s = 46;
	{8'd236,8'd185} : s = 155;
	{8'd236,8'd186} : s = 151;
	{8'd236,8'd187} : s = 303;
	{8'd236,8'd188} : s = 45;
	{8'd236,8'd189} : s = 143;
	{8'd236,8'd190} : s = 124;
	{8'd236,8'd191} : s = 287;
	{8'd236,8'd192} : s = 122;
	{8'd236,8'd193} : s = 252;
	{8'd236,8'd194} : s = 250;
	{8'd236,8'd195} : s = 445;
	{8'd236,8'd196} : s = 43;
	{8'd236,8'd197} : s = 121;
	{8'd236,8'd198} : s = 118;
	{8'd236,8'd199} : s = 249;
	{8'd236,8'd200} : s = 117;
	{8'd236,8'd201} : s = 246;
	{8'd236,8'd202} : s = 245;
	{8'd236,8'd203} : s = 443;
	{8'd236,8'd204} : s = 115;
	{8'd236,8'd205} : s = 243;
	{8'd236,8'd206} : s = 238;
	{8'd236,8'd207} : s = 439;
	{8'd236,8'd208} : s = 237;
	{8'd236,8'd209} : s = 431;
	{8'd236,8'd210} : s = 415;
	{8'd236,8'd211} : s = 507;
	{8'd236,8'd212} : s = 7;
	{8'd236,8'd213} : s = 39;
	{8'd236,8'd214} : s = 30;
	{8'd236,8'd215} : s = 110;
	{8'd236,8'd216} : s = 29;
	{8'd236,8'd217} : s = 109;
	{8'd236,8'd218} : s = 107;
	{8'd236,8'd219} : s = 235;
	{8'd236,8'd220} : s = 27;
	{8'd236,8'd221} : s = 103;
	{8'd236,8'd222} : s = 94;
	{8'd236,8'd223} : s = 231;
	{8'd236,8'd224} : s = 93;
	{8'd236,8'd225} : s = 222;
	{8'd236,8'd226} : s = 221;
	{8'd236,8'd227} : s = 382;
	{8'd236,8'd228} : s = 23;
	{8'd236,8'd229} : s = 91;
	{8'd236,8'd230} : s = 87;
	{8'd236,8'd231} : s = 219;
	{8'd236,8'd232} : s = 79;
	{8'd236,8'd233} : s = 215;
	{8'd236,8'd234} : s = 207;
	{8'd236,8'd235} : s = 381;
	{8'd236,8'd236} : s = 62;
	{8'd236,8'd237} : s = 190;
	{8'd236,8'd238} : s = 189;
	{8'd236,8'd239} : s = 379;
	{8'd236,8'd240} : s = 187;
	{8'd236,8'd241} : s = 375;
	{8'd236,8'd242} : s = 367;
	{8'd236,8'd243} : s = 503;
	{8'd236,8'd244} : s = 15;
	{8'd236,8'd245} : s = 61;
	{8'd236,8'd246} : s = 59;
	{8'd236,8'd247} : s = 183;
	{8'd236,8'd248} : s = 55;
	{8'd236,8'd249} : s = 175;
	{8'd236,8'd250} : s = 159;
	{8'd236,8'd251} : s = 351;
	{8'd236,8'd252} : s = 47;
	{8'd236,8'd253} : s = 126;
	{8'd236,8'd254} : s = 125;
	{8'd236,8'd255} : s = 319;
	{8'd237,8'd0} : s = 444;
	{8'd237,8'd1} : s = 442;
	{8'd237,8'd2} : s = 502;
	{8'd237,8'd3} : s = 197;
	{8'd237,8'd4} : s = 333;
	{8'd237,8'd5} : s = 331;
	{8'd237,8'd6} : s = 441;
	{8'd237,8'd7} : s = 327;
	{8'd237,8'd8} : s = 438;
	{8'd237,8'd9} : s = 437;
	{8'd237,8'd10} : s = 501;
	{8'd237,8'd11} : s = 316;
	{8'd237,8'd12} : s = 435;
	{8'd237,8'd13} : s = 430;
	{8'd237,8'd14} : s = 499;
	{8'd237,8'd15} : s = 429;
	{8'd237,8'd16} : s = 494;
	{8'd237,8'd17} : s = 493;
	{8'd237,8'd18} : s = 510;
	{8'd237,8'd19} : s = 1;
	{8'd237,8'd20} : s = 18;
	{8'd237,8'd21} : s = 17;
	{8'd237,8'd22} : s = 82;
	{8'd237,8'd23} : s = 12;
	{8'd237,8'd24} : s = 81;
	{8'd237,8'd25} : s = 76;
	{8'd237,8'd26} : s = 195;
	{8'd237,8'd27} : s = 10;
	{8'd237,8'd28} : s = 74;
	{8'd237,8'd29} : s = 73;
	{8'd237,8'd30} : s = 184;
	{8'd237,8'd31} : s = 70;
	{8'd237,8'd32} : s = 180;
	{8'd237,8'd33} : s = 178;
	{8'd237,8'd34} : s = 314;
	{8'd237,8'd35} : s = 9;
	{8'd237,8'd36} : s = 69;
	{8'd237,8'd37} : s = 67;
	{8'd237,8'd38} : s = 177;
	{8'd237,8'd39} : s = 56;
	{8'd237,8'd40} : s = 172;
	{8'd237,8'd41} : s = 170;
	{8'd237,8'd42} : s = 313;
	{8'd237,8'd43} : s = 52;
	{8'd237,8'd44} : s = 169;
	{8'd237,8'd45} : s = 166;
	{8'd237,8'd46} : s = 310;
	{8'd237,8'd47} : s = 165;
	{8'd237,8'd48} : s = 309;
	{8'd237,8'd49} : s = 307;
	{8'd237,8'd50} : s = 427;
	{8'd237,8'd51} : s = 6;
	{8'd237,8'd52} : s = 50;
	{8'd237,8'd53} : s = 49;
	{8'd237,8'd54} : s = 163;
	{8'd237,8'd55} : s = 44;
	{8'd237,8'd56} : s = 156;
	{8'd237,8'd57} : s = 154;
	{8'd237,8'd58} : s = 302;
	{8'd237,8'd59} : s = 42;
	{8'd237,8'd60} : s = 153;
	{8'd237,8'd61} : s = 150;
	{8'd237,8'd62} : s = 301;
	{8'd237,8'd63} : s = 149;
	{8'd237,8'd64} : s = 299;
	{8'd237,8'd65} : s = 295;
	{8'd237,8'd66} : s = 423;
	{8'd237,8'd67} : s = 41;
	{8'd237,8'd68} : s = 147;
	{8'd237,8'd69} : s = 142;
	{8'd237,8'd70} : s = 286;
	{8'd237,8'd71} : s = 141;
	{8'd237,8'd72} : s = 285;
	{8'd237,8'd73} : s = 283;
	{8'd237,8'd74} : s = 414;
	{8'd237,8'd75} : s = 139;
	{8'd237,8'd76} : s = 279;
	{8'd237,8'd77} : s = 271;
	{8'd237,8'd78} : s = 413;
	{8'd237,8'd79} : s = 248;
	{8'd237,8'd80} : s = 411;
	{8'd237,8'd81} : s = 407;
	{8'd237,8'd82} : s = 491;
	{8'd237,8'd83} : s = 5;
	{8'd237,8'd84} : s = 38;
	{8'd237,8'd85} : s = 37;
	{8'd237,8'd86} : s = 135;
	{8'd237,8'd87} : s = 35;
	{8'd237,8'd88} : s = 120;
	{8'd237,8'd89} : s = 116;
	{8'd237,8'd90} : s = 244;
	{8'd237,8'd91} : s = 28;
	{8'd237,8'd92} : s = 114;
	{8'd237,8'd93} : s = 113;
	{8'd237,8'd94} : s = 242;
	{8'd237,8'd95} : s = 108;
	{8'd237,8'd96} : s = 241;
	{8'd237,8'd97} : s = 236;
	{8'd237,8'd98} : s = 399;
	{8'd237,8'd99} : s = 26;
	{8'd237,8'd100} : s = 106;
	{8'd237,8'd101} : s = 105;
	{8'd237,8'd102} : s = 234;
	{8'd237,8'd103} : s = 102;
	{8'd237,8'd104} : s = 233;
	{8'd237,8'd105} : s = 230;
	{8'd237,8'd106} : s = 380;
	{8'd237,8'd107} : s = 101;
	{8'd237,8'd108} : s = 229;
	{8'd237,8'd109} : s = 227;
	{8'd237,8'd110} : s = 378;
	{8'd237,8'd111} : s = 220;
	{8'd237,8'd112} : s = 377;
	{8'd237,8'd113} : s = 374;
	{8'd237,8'd114} : s = 487;
	{8'd237,8'd115} : s = 25;
	{8'd237,8'd116} : s = 99;
	{8'd237,8'd117} : s = 92;
	{8'd237,8'd118} : s = 218;
	{8'd237,8'd119} : s = 90;
	{8'd237,8'd120} : s = 217;
	{8'd237,8'd121} : s = 214;
	{8'd237,8'd122} : s = 373;
	{8'd237,8'd123} : s = 89;
	{8'd237,8'd124} : s = 213;
	{8'd237,8'd125} : s = 211;
	{8'd237,8'd126} : s = 371;
	{8'd237,8'd127} : s = 206;
	{8'd237,8'd128} : s = 366;
	{8'd237,8'd129} : s = 365;
	{8'd237,8'd130} : s = 478;
	{8'd237,8'd131} : s = 86;
	{8'd237,8'd132} : s = 205;
	{8'd237,8'd133} : s = 203;
	{8'd237,8'd134} : s = 363;
	{8'd237,8'd135} : s = 199;
	{8'd237,8'd136} : s = 359;
	{8'd237,8'd137} : s = 350;
	{8'd237,8'd138} : s = 477;
	{8'd237,8'd139} : s = 188;
	{8'd237,8'd140} : s = 349;
	{8'd237,8'd141} : s = 347;
	{8'd237,8'd142} : s = 475;
	{8'd237,8'd143} : s = 343;
	{8'd237,8'd144} : s = 471;
	{8'd237,8'd145} : s = 463;
	{8'd237,8'd146} : s = 509;
	{8'd237,8'd147} : s = 3;
	{8'd237,8'd148} : s = 22;
	{8'd237,8'd149} : s = 21;
	{8'd237,8'd150} : s = 85;
	{8'd237,8'd151} : s = 19;
	{8'd237,8'd152} : s = 83;
	{8'd237,8'd153} : s = 78;
	{8'd237,8'd154} : s = 186;
	{8'd237,8'd155} : s = 14;
	{8'd237,8'd156} : s = 77;
	{8'd237,8'd157} : s = 75;
	{8'd237,8'd158} : s = 185;
	{8'd237,8'd159} : s = 71;
	{8'd237,8'd160} : s = 182;
	{8'd237,8'd161} : s = 181;
	{8'd237,8'd162} : s = 335;
	{8'd237,8'd163} : s = 13;
	{8'd237,8'd164} : s = 60;
	{8'd237,8'd165} : s = 58;
	{8'd237,8'd166} : s = 179;
	{8'd237,8'd167} : s = 57;
	{8'd237,8'd168} : s = 174;
	{8'd237,8'd169} : s = 173;
	{8'd237,8'd170} : s = 318;
	{8'd237,8'd171} : s = 54;
	{8'd237,8'd172} : s = 171;
	{8'd237,8'd173} : s = 167;
	{8'd237,8'd174} : s = 317;
	{8'd237,8'd175} : s = 158;
	{8'd237,8'd176} : s = 315;
	{8'd237,8'd177} : s = 311;
	{8'd237,8'd178} : s = 446;
	{8'd237,8'd179} : s = 11;
	{8'd237,8'd180} : s = 53;
	{8'd237,8'd181} : s = 51;
	{8'd237,8'd182} : s = 157;
	{8'd237,8'd183} : s = 46;
	{8'd237,8'd184} : s = 155;
	{8'd237,8'd185} : s = 151;
	{8'd237,8'd186} : s = 303;
	{8'd237,8'd187} : s = 45;
	{8'd237,8'd188} : s = 143;
	{8'd237,8'd189} : s = 124;
	{8'd237,8'd190} : s = 287;
	{8'd237,8'd191} : s = 122;
	{8'd237,8'd192} : s = 252;
	{8'd237,8'd193} : s = 250;
	{8'd237,8'd194} : s = 445;
	{8'd237,8'd195} : s = 43;
	{8'd237,8'd196} : s = 121;
	{8'd237,8'd197} : s = 118;
	{8'd237,8'd198} : s = 249;
	{8'd237,8'd199} : s = 117;
	{8'd237,8'd200} : s = 246;
	{8'd237,8'd201} : s = 245;
	{8'd237,8'd202} : s = 443;
	{8'd237,8'd203} : s = 115;
	{8'd237,8'd204} : s = 243;
	{8'd237,8'd205} : s = 238;
	{8'd237,8'd206} : s = 439;
	{8'd237,8'd207} : s = 237;
	{8'd237,8'd208} : s = 431;
	{8'd237,8'd209} : s = 415;
	{8'd237,8'd210} : s = 507;
	{8'd237,8'd211} : s = 7;
	{8'd237,8'd212} : s = 39;
	{8'd237,8'd213} : s = 30;
	{8'd237,8'd214} : s = 110;
	{8'd237,8'd215} : s = 29;
	{8'd237,8'd216} : s = 109;
	{8'd237,8'd217} : s = 107;
	{8'd237,8'd218} : s = 235;
	{8'd237,8'd219} : s = 27;
	{8'd237,8'd220} : s = 103;
	{8'd237,8'd221} : s = 94;
	{8'd237,8'd222} : s = 231;
	{8'd237,8'd223} : s = 93;
	{8'd237,8'd224} : s = 222;
	{8'd237,8'd225} : s = 221;
	{8'd237,8'd226} : s = 382;
	{8'd237,8'd227} : s = 23;
	{8'd237,8'd228} : s = 91;
	{8'd237,8'd229} : s = 87;
	{8'd237,8'd230} : s = 219;
	{8'd237,8'd231} : s = 79;
	{8'd237,8'd232} : s = 215;
	{8'd237,8'd233} : s = 207;
	{8'd237,8'd234} : s = 381;
	{8'd237,8'd235} : s = 62;
	{8'd237,8'd236} : s = 190;
	{8'd237,8'd237} : s = 189;
	{8'd237,8'd238} : s = 379;
	{8'd237,8'd239} : s = 187;
	{8'd237,8'd240} : s = 375;
	{8'd237,8'd241} : s = 367;
	{8'd237,8'd242} : s = 503;
	{8'd237,8'd243} : s = 15;
	{8'd237,8'd244} : s = 61;
	{8'd237,8'd245} : s = 59;
	{8'd237,8'd246} : s = 183;
	{8'd237,8'd247} : s = 55;
	{8'd237,8'd248} : s = 175;
	{8'd237,8'd249} : s = 159;
	{8'd237,8'd250} : s = 351;
	{8'd237,8'd251} : s = 47;
	{8'd237,8'd252} : s = 126;
	{8'd237,8'd253} : s = 125;
	{8'd237,8'd254} : s = 319;
	{8'd237,8'd255} : s = 123;
	{8'd238,8'd0} : s = 442;
	{8'd238,8'd1} : s = 502;
	{8'd238,8'd2} : s = 197;
	{8'd238,8'd3} : s = 333;
	{8'd238,8'd4} : s = 331;
	{8'd238,8'd5} : s = 441;
	{8'd238,8'd6} : s = 327;
	{8'd238,8'd7} : s = 438;
	{8'd238,8'd8} : s = 437;
	{8'd238,8'd9} : s = 501;
	{8'd238,8'd10} : s = 316;
	{8'd238,8'd11} : s = 435;
	{8'd238,8'd12} : s = 430;
	{8'd238,8'd13} : s = 499;
	{8'd238,8'd14} : s = 429;
	{8'd238,8'd15} : s = 494;
	{8'd238,8'd16} : s = 493;
	{8'd238,8'd17} : s = 510;
	{8'd238,8'd18} : s = 1;
	{8'd238,8'd19} : s = 18;
	{8'd238,8'd20} : s = 17;
	{8'd238,8'd21} : s = 82;
	{8'd238,8'd22} : s = 12;
	{8'd238,8'd23} : s = 81;
	{8'd238,8'd24} : s = 76;
	{8'd238,8'd25} : s = 195;
	{8'd238,8'd26} : s = 10;
	{8'd238,8'd27} : s = 74;
	{8'd238,8'd28} : s = 73;
	{8'd238,8'd29} : s = 184;
	{8'd238,8'd30} : s = 70;
	{8'd238,8'd31} : s = 180;
	{8'd238,8'd32} : s = 178;
	{8'd238,8'd33} : s = 314;
	{8'd238,8'd34} : s = 9;
	{8'd238,8'd35} : s = 69;
	{8'd238,8'd36} : s = 67;
	{8'd238,8'd37} : s = 177;
	{8'd238,8'd38} : s = 56;
	{8'd238,8'd39} : s = 172;
	{8'd238,8'd40} : s = 170;
	{8'd238,8'd41} : s = 313;
	{8'd238,8'd42} : s = 52;
	{8'd238,8'd43} : s = 169;
	{8'd238,8'd44} : s = 166;
	{8'd238,8'd45} : s = 310;
	{8'd238,8'd46} : s = 165;
	{8'd238,8'd47} : s = 309;
	{8'd238,8'd48} : s = 307;
	{8'd238,8'd49} : s = 427;
	{8'd238,8'd50} : s = 6;
	{8'd238,8'd51} : s = 50;
	{8'd238,8'd52} : s = 49;
	{8'd238,8'd53} : s = 163;
	{8'd238,8'd54} : s = 44;
	{8'd238,8'd55} : s = 156;
	{8'd238,8'd56} : s = 154;
	{8'd238,8'd57} : s = 302;
	{8'd238,8'd58} : s = 42;
	{8'd238,8'd59} : s = 153;
	{8'd238,8'd60} : s = 150;
	{8'd238,8'd61} : s = 301;
	{8'd238,8'd62} : s = 149;
	{8'd238,8'd63} : s = 299;
	{8'd238,8'd64} : s = 295;
	{8'd238,8'd65} : s = 423;
	{8'd238,8'd66} : s = 41;
	{8'd238,8'd67} : s = 147;
	{8'd238,8'd68} : s = 142;
	{8'd238,8'd69} : s = 286;
	{8'd238,8'd70} : s = 141;
	{8'd238,8'd71} : s = 285;
	{8'd238,8'd72} : s = 283;
	{8'd238,8'd73} : s = 414;
	{8'd238,8'd74} : s = 139;
	{8'd238,8'd75} : s = 279;
	{8'd238,8'd76} : s = 271;
	{8'd238,8'd77} : s = 413;
	{8'd238,8'd78} : s = 248;
	{8'd238,8'd79} : s = 411;
	{8'd238,8'd80} : s = 407;
	{8'd238,8'd81} : s = 491;
	{8'd238,8'd82} : s = 5;
	{8'd238,8'd83} : s = 38;
	{8'd238,8'd84} : s = 37;
	{8'd238,8'd85} : s = 135;
	{8'd238,8'd86} : s = 35;
	{8'd238,8'd87} : s = 120;
	{8'd238,8'd88} : s = 116;
	{8'd238,8'd89} : s = 244;
	{8'd238,8'd90} : s = 28;
	{8'd238,8'd91} : s = 114;
	{8'd238,8'd92} : s = 113;
	{8'd238,8'd93} : s = 242;
	{8'd238,8'd94} : s = 108;
	{8'd238,8'd95} : s = 241;
	{8'd238,8'd96} : s = 236;
	{8'd238,8'd97} : s = 399;
	{8'd238,8'd98} : s = 26;
	{8'd238,8'd99} : s = 106;
	{8'd238,8'd100} : s = 105;
	{8'd238,8'd101} : s = 234;
	{8'd238,8'd102} : s = 102;
	{8'd238,8'd103} : s = 233;
	{8'd238,8'd104} : s = 230;
	{8'd238,8'd105} : s = 380;
	{8'd238,8'd106} : s = 101;
	{8'd238,8'd107} : s = 229;
	{8'd238,8'd108} : s = 227;
	{8'd238,8'd109} : s = 378;
	{8'd238,8'd110} : s = 220;
	{8'd238,8'd111} : s = 377;
	{8'd238,8'd112} : s = 374;
	{8'd238,8'd113} : s = 487;
	{8'd238,8'd114} : s = 25;
	{8'd238,8'd115} : s = 99;
	{8'd238,8'd116} : s = 92;
	{8'd238,8'd117} : s = 218;
	{8'd238,8'd118} : s = 90;
	{8'd238,8'd119} : s = 217;
	{8'd238,8'd120} : s = 214;
	{8'd238,8'd121} : s = 373;
	{8'd238,8'd122} : s = 89;
	{8'd238,8'd123} : s = 213;
	{8'd238,8'd124} : s = 211;
	{8'd238,8'd125} : s = 371;
	{8'd238,8'd126} : s = 206;
	{8'd238,8'd127} : s = 366;
	{8'd238,8'd128} : s = 365;
	{8'd238,8'd129} : s = 478;
	{8'd238,8'd130} : s = 86;
	{8'd238,8'd131} : s = 205;
	{8'd238,8'd132} : s = 203;
	{8'd238,8'd133} : s = 363;
	{8'd238,8'd134} : s = 199;
	{8'd238,8'd135} : s = 359;
	{8'd238,8'd136} : s = 350;
	{8'd238,8'd137} : s = 477;
	{8'd238,8'd138} : s = 188;
	{8'd238,8'd139} : s = 349;
	{8'd238,8'd140} : s = 347;
	{8'd238,8'd141} : s = 475;
	{8'd238,8'd142} : s = 343;
	{8'd238,8'd143} : s = 471;
	{8'd238,8'd144} : s = 463;
	{8'd238,8'd145} : s = 509;
	{8'd238,8'd146} : s = 3;
	{8'd238,8'd147} : s = 22;
	{8'd238,8'd148} : s = 21;
	{8'd238,8'd149} : s = 85;
	{8'd238,8'd150} : s = 19;
	{8'd238,8'd151} : s = 83;
	{8'd238,8'd152} : s = 78;
	{8'd238,8'd153} : s = 186;
	{8'd238,8'd154} : s = 14;
	{8'd238,8'd155} : s = 77;
	{8'd238,8'd156} : s = 75;
	{8'd238,8'd157} : s = 185;
	{8'd238,8'd158} : s = 71;
	{8'd238,8'd159} : s = 182;
	{8'd238,8'd160} : s = 181;
	{8'd238,8'd161} : s = 335;
	{8'd238,8'd162} : s = 13;
	{8'd238,8'd163} : s = 60;
	{8'd238,8'd164} : s = 58;
	{8'd238,8'd165} : s = 179;
	{8'd238,8'd166} : s = 57;
	{8'd238,8'd167} : s = 174;
	{8'd238,8'd168} : s = 173;
	{8'd238,8'd169} : s = 318;
	{8'd238,8'd170} : s = 54;
	{8'd238,8'd171} : s = 171;
	{8'd238,8'd172} : s = 167;
	{8'd238,8'd173} : s = 317;
	{8'd238,8'd174} : s = 158;
	{8'd238,8'd175} : s = 315;
	{8'd238,8'd176} : s = 311;
	{8'd238,8'd177} : s = 446;
	{8'd238,8'd178} : s = 11;
	{8'd238,8'd179} : s = 53;
	{8'd238,8'd180} : s = 51;
	{8'd238,8'd181} : s = 157;
	{8'd238,8'd182} : s = 46;
	{8'd238,8'd183} : s = 155;
	{8'd238,8'd184} : s = 151;
	{8'd238,8'd185} : s = 303;
	{8'd238,8'd186} : s = 45;
	{8'd238,8'd187} : s = 143;
	{8'd238,8'd188} : s = 124;
	{8'd238,8'd189} : s = 287;
	{8'd238,8'd190} : s = 122;
	{8'd238,8'd191} : s = 252;
	{8'd238,8'd192} : s = 250;
	{8'd238,8'd193} : s = 445;
	{8'd238,8'd194} : s = 43;
	{8'd238,8'd195} : s = 121;
	{8'd238,8'd196} : s = 118;
	{8'd238,8'd197} : s = 249;
	{8'd238,8'd198} : s = 117;
	{8'd238,8'd199} : s = 246;
	{8'd238,8'd200} : s = 245;
	{8'd238,8'd201} : s = 443;
	{8'd238,8'd202} : s = 115;
	{8'd238,8'd203} : s = 243;
	{8'd238,8'd204} : s = 238;
	{8'd238,8'd205} : s = 439;
	{8'd238,8'd206} : s = 237;
	{8'd238,8'd207} : s = 431;
	{8'd238,8'd208} : s = 415;
	{8'd238,8'd209} : s = 507;
	{8'd238,8'd210} : s = 7;
	{8'd238,8'd211} : s = 39;
	{8'd238,8'd212} : s = 30;
	{8'd238,8'd213} : s = 110;
	{8'd238,8'd214} : s = 29;
	{8'd238,8'd215} : s = 109;
	{8'd238,8'd216} : s = 107;
	{8'd238,8'd217} : s = 235;
	{8'd238,8'd218} : s = 27;
	{8'd238,8'd219} : s = 103;
	{8'd238,8'd220} : s = 94;
	{8'd238,8'd221} : s = 231;
	{8'd238,8'd222} : s = 93;
	{8'd238,8'd223} : s = 222;
	{8'd238,8'd224} : s = 221;
	{8'd238,8'd225} : s = 382;
	{8'd238,8'd226} : s = 23;
	{8'd238,8'd227} : s = 91;
	{8'd238,8'd228} : s = 87;
	{8'd238,8'd229} : s = 219;
	{8'd238,8'd230} : s = 79;
	{8'd238,8'd231} : s = 215;
	{8'd238,8'd232} : s = 207;
	{8'd238,8'd233} : s = 381;
	{8'd238,8'd234} : s = 62;
	{8'd238,8'd235} : s = 190;
	{8'd238,8'd236} : s = 189;
	{8'd238,8'd237} : s = 379;
	{8'd238,8'd238} : s = 187;
	{8'd238,8'd239} : s = 375;
	{8'd238,8'd240} : s = 367;
	{8'd238,8'd241} : s = 503;
	{8'd238,8'd242} : s = 15;
	{8'd238,8'd243} : s = 61;
	{8'd238,8'd244} : s = 59;
	{8'd238,8'd245} : s = 183;
	{8'd238,8'd246} : s = 55;
	{8'd238,8'd247} : s = 175;
	{8'd238,8'd248} : s = 159;
	{8'd238,8'd249} : s = 351;
	{8'd238,8'd250} : s = 47;
	{8'd238,8'd251} : s = 126;
	{8'd238,8'd252} : s = 125;
	{8'd238,8'd253} : s = 319;
	{8'd238,8'd254} : s = 123;
	{8'd238,8'd255} : s = 254;
	{8'd239,8'd0} : s = 502;
	{8'd239,8'd1} : s = 197;
	{8'd239,8'd2} : s = 333;
	{8'd239,8'd3} : s = 331;
	{8'd239,8'd4} : s = 441;
	{8'd239,8'd5} : s = 327;
	{8'd239,8'd6} : s = 438;
	{8'd239,8'd7} : s = 437;
	{8'd239,8'd8} : s = 501;
	{8'd239,8'd9} : s = 316;
	{8'd239,8'd10} : s = 435;
	{8'd239,8'd11} : s = 430;
	{8'd239,8'd12} : s = 499;
	{8'd239,8'd13} : s = 429;
	{8'd239,8'd14} : s = 494;
	{8'd239,8'd15} : s = 493;
	{8'd239,8'd16} : s = 510;
	{8'd239,8'd17} : s = 1;
	{8'd239,8'd18} : s = 18;
	{8'd239,8'd19} : s = 17;
	{8'd239,8'd20} : s = 82;
	{8'd239,8'd21} : s = 12;
	{8'd239,8'd22} : s = 81;
	{8'd239,8'd23} : s = 76;
	{8'd239,8'd24} : s = 195;
	{8'd239,8'd25} : s = 10;
	{8'd239,8'd26} : s = 74;
	{8'd239,8'd27} : s = 73;
	{8'd239,8'd28} : s = 184;
	{8'd239,8'd29} : s = 70;
	{8'd239,8'd30} : s = 180;
	{8'd239,8'd31} : s = 178;
	{8'd239,8'd32} : s = 314;
	{8'd239,8'd33} : s = 9;
	{8'd239,8'd34} : s = 69;
	{8'd239,8'd35} : s = 67;
	{8'd239,8'd36} : s = 177;
	{8'd239,8'd37} : s = 56;
	{8'd239,8'd38} : s = 172;
	{8'd239,8'd39} : s = 170;
	{8'd239,8'd40} : s = 313;
	{8'd239,8'd41} : s = 52;
	{8'd239,8'd42} : s = 169;
	{8'd239,8'd43} : s = 166;
	{8'd239,8'd44} : s = 310;
	{8'd239,8'd45} : s = 165;
	{8'd239,8'd46} : s = 309;
	{8'd239,8'd47} : s = 307;
	{8'd239,8'd48} : s = 427;
	{8'd239,8'd49} : s = 6;
	{8'd239,8'd50} : s = 50;
	{8'd239,8'd51} : s = 49;
	{8'd239,8'd52} : s = 163;
	{8'd239,8'd53} : s = 44;
	{8'd239,8'd54} : s = 156;
	{8'd239,8'd55} : s = 154;
	{8'd239,8'd56} : s = 302;
	{8'd239,8'd57} : s = 42;
	{8'd239,8'd58} : s = 153;
	{8'd239,8'd59} : s = 150;
	{8'd239,8'd60} : s = 301;
	{8'd239,8'd61} : s = 149;
	{8'd239,8'd62} : s = 299;
	{8'd239,8'd63} : s = 295;
	{8'd239,8'd64} : s = 423;
	{8'd239,8'd65} : s = 41;
	{8'd239,8'd66} : s = 147;
	{8'd239,8'd67} : s = 142;
	{8'd239,8'd68} : s = 286;
	{8'd239,8'd69} : s = 141;
	{8'd239,8'd70} : s = 285;
	{8'd239,8'd71} : s = 283;
	{8'd239,8'd72} : s = 414;
	{8'd239,8'd73} : s = 139;
	{8'd239,8'd74} : s = 279;
	{8'd239,8'd75} : s = 271;
	{8'd239,8'd76} : s = 413;
	{8'd239,8'd77} : s = 248;
	{8'd239,8'd78} : s = 411;
	{8'd239,8'd79} : s = 407;
	{8'd239,8'd80} : s = 491;
	{8'd239,8'd81} : s = 5;
	{8'd239,8'd82} : s = 38;
	{8'd239,8'd83} : s = 37;
	{8'd239,8'd84} : s = 135;
	{8'd239,8'd85} : s = 35;
	{8'd239,8'd86} : s = 120;
	{8'd239,8'd87} : s = 116;
	{8'd239,8'd88} : s = 244;
	{8'd239,8'd89} : s = 28;
	{8'd239,8'd90} : s = 114;
	{8'd239,8'd91} : s = 113;
	{8'd239,8'd92} : s = 242;
	{8'd239,8'd93} : s = 108;
	{8'd239,8'd94} : s = 241;
	{8'd239,8'd95} : s = 236;
	{8'd239,8'd96} : s = 399;
	{8'd239,8'd97} : s = 26;
	{8'd239,8'd98} : s = 106;
	{8'd239,8'd99} : s = 105;
	{8'd239,8'd100} : s = 234;
	{8'd239,8'd101} : s = 102;
	{8'd239,8'd102} : s = 233;
	{8'd239,8'd103} : s = 230;
	{8'd239,8'd104} : s = 380;
	{8'd239,8'd105} : s = 101;
	{8'd239,8'd106} : s = 229;
	{8'd239,8'd107} : s = 227;
	{8'd239,8'd108} : s = 378;
	{8'd239,8'd109} : s = 220;
	{8'd239,8'd110} : s = 377;
	{8'd239,8'd111} : s = 374;
	{8'd239,8'd112} : s = 487;
	{8'd239,8'd113} : s = 25;
	{8'd239,8'd114} : s = 99;
	{8'd239,8'd115} : s = 92;
	{8'd239,8'd116} : s = 218;
	{8'd239,8'd117} : s = 90;
	{8'd239,8'd118} : s = 217;
	{8'd239,8'd119} : s = 214;
	{8'd239,8'd120} : s = 373;
	{8'd239,8'd121} : s = 89;
	{8'd239,8'd122} : s = 213;
	{8'd239,8'd123} : s = 211;
	{8'd239,8'd124} : s = 371;
	{8'd239,8'd125} : s = 206;
	{8'd239,8'd126} : s = 366;
	{8'd239,8'd127} : s = 365;
	{8'd239,8'd128} : s = 478;
	{8'd239,8'd129} : s = 86;
	{8'd239,8'd130} : s = 205;
	{8'd239,8'd131} : s = 203;
	{8'd239,8'd132} : s = 363;
	{8'd239,8'd133} : s = 199;
	{8'd239,8'd134} : s = 359;
	{8'd239,8'd135} : s = 350;
	{8'd239,8'd136} : s = 477;
	{8'd239,8'd137} : s = 188;
	{8'd239,8'd138} : s = 349;
	{8'd239,8'd139} : s = 347;
	{8'd239,8'd140} : s = 475;
	{8'd239,8'd141} : s = 343;
	{8'd239,8'd142} : s = 471;
	{8'd239,8'd143} : s = 463;
	{8'd239,8'd144} : s = 509;
	{8'd239,8'd145} : s = 3;
	{8'd239,8'd146} : s = 22;
	{8'd239,8'd147} : s = 21;
	{8'd239,8'd148} : s = 85;
	{8'd239,8'd149} : s = 19;
	{8'd239,8'd150} : s = 83;
	{8'd239,8'd151} : s = 78;
	{8'd239,8'd152} : s = 186;
	{8'd239,8'd153} : s = 14;
	{8'd239,8'd154} : s = 77;
	{8'd239,8'd155} : s = 75;
	{8'd239,8'd156} : s = 185;
	{8'd239,8'd157} : s = 71;
	{8'd239,8'd158} : s = 182;
	{8'd239,8'd159} : s = 181;
	{8'd239,8'd160} : s = 335;
	{8'd239,8'd161} : s = 13;
	{8'd239,8'd162} : s = 60;
	{8'd239,8'd163} : s = 58;
	{8'd239,8'd164} : s = 179;
	{8'd239,8'd165} : s = 57;
	{8'd239,8'd166} : s = 174;
	{8'd239,8'd167} : s = 173;
	{8'd239,8'd168} : s = 318;
	{8'd239,8'd169} : s = 54;
	{8'd239,8'd170} : s = 171;
	{8'd239,8'd171} : s = 167;
	{8'd239,8'd172} : s = 317;
	{8'd239,8'd173} : s = 158;
	{8'd239,8'd174} : s = 315;
	{8'd239,8'd175} : s = 311;
	{8'd239,8'd176} : s = 446;
	{8'd239,8'd177} : s = 11;
	{8'd239,8'd178} : s = 53;
	{8'd239,8'd179} : s = 51;
	{8'd239,8'd180} : s = 157;
	{8'd239,8'd181} : s = 46;
	{8'd239,8'd182} : s = 155;
	{8'd239,8'd183} : s = 151;
	{8'd239,8'd184} : s = 303;
	{8'd239,8'd185} : s = 45;
	{8'd239,8'd186} : s = 143;
	{8'd239,8'd187} : s = 124;
	{8'd239,8'd188} : s = 287;
	{8'd239,8'd189} : s = 122;
	{8'd239,8'd190} : s = 252;
	{8'd239,8'd191} : s = 250;
	{8'd239,8'd192} : s = 445;
	{8'd239,8'd193} : s = 43;
	{8'd239,8'd194} : s = 121;
	{8'd239,8'd195} : s = 118;
	{8'd239,8'd196} : s = 249;
	{8'd239,8'd197} : s = 117;
	{8'd239,8'd198} : s = 246;
	{8'd239,8'd199} : s = 245;
	{8'd239,8'd200} : s = 443;
	{8'd239,8'd201} : s = 115;
	{8'd239,8'd202} : s = 243;
	{8'd239,8'd203} : s = 238;
	{8'd239,8'd204} : s = 439;
	{8'd239,8'd205} : s = 237;
	{8'd239,8'd206} : s = 431;
	{8'd239,8'd207} : s = 415;
	{8'd239,8'd208} : s = 507;
	{8'd239,8'd209} : s = 7;
	{8'd239,8'd210} : s = 39;
	{8'd239,8'd211} : s = 30;
	{8'd239,8'd212} : s = 110;
	{8'd239,8'd213} : s = 29;
	{8'd239,8'd214} : s = 109;
	{8'd239,8'd215} : s = 107;
	{8'd239,8'd216} : s = 235;
	{8'd239,8'd217} : s = 27;
	{8'd239,8'd218} : s = 103;
	{8'd239,8'd219} : s = 94;
	{8'd239,8'd220} : s = 231;
	{8'd239,8'd221} : s = 93;
	{8'd239,8'd222} : s = 222;
	{8'd239,8'd223} : s = 221;
	{8'd239,8'd224} : s = 382;
	{8'd239,8'd225} : s = 23;
	{8'd239,8'd226} : s = 91;
	{8'd239,8'd227} : s = 87;
	{8'd239,8'd228} : s = 219;
	{8'd239,8'd229} : s = 79;
	{8'd239,8'd230} : s = 215;
	{8'd239,8'd231} : s = 207;
	{8'd239,8'd232} : s = 381;
	{8'd239,8'd233} : s = 62;
	{8'd239,8'd234} : s = 190;
	{8'd239,8'd235} : s = 189;
	{8'd239,8'd236} : s = 379;
	{8'd239,8'd237} : s = 187;
	{8'd239,8'd238} : s = 375;
	{8'd239,8'd239} : s = 367;
	{8'd239,8'd240} : s = 503;
	{8'd239,8'd241} : s = 15;
	{8'd239,8'd242} : s = 61;
	{8'd239,8'd243} : s = 59;
	{8'd239,8'd244} : s = 183;
	{8'd239,8'd245} : s = 55;
	{8'd239,8'd246} : s = 175;
	{8'd239,8'd247} : s = 159;
	{8'd239,8'd248} : s = 351;
	{8'd239,8'd249} : s = 47;
	{8'd239,8'd250} : s = 126;
	{8'd239,8'd251} : s = 125;
	{8'd239,8'd252} : s = 319;
	{8'd239,8'd253} : s = 123;
	{8'd239,8'd254} : s = 254;
	{8'd239,8'd255} : s = 253;
	{8'd240,8'd0} : s = 197;
	{8'd240,8'd1} : s = 333;
	{8'd240,8'd2} : s = 331;
	{8'd240,8'd3} : s = 441;
	{8'd240,8'd4} : s = 327;
	{8'd240,8'd5} : s = 438;
	{8'd240,8'd6} : s = 437;
	{8'd240,8'd7} : s = 501;
	{8'd240,8'd8} : s = 316;
	{8'd240,8'd9} : s = 435;
	{8'd240,8'd10} : s = 430;
	{8'd240,8'd11} : s = 499;
	{8'd240,8'd12} : s = 429;
	{8'd240,8'd13} : s = 494;
	{8'd240,8'd14} : s = 493;
	{8'd240,8'd15} : s = 510;
	{8'd240,8'd16} : s = 1;
	{8'd240,8'd17} : s = 18;
	{8'd240,8'd18} : s = 17;
	{8'd240,8'd19} : s = 82;
	{8'd240,8'd20} : s = 12;
	{8'd240,8'd21} : s = 81;
	{8'd240,8'd22} : s = 76;
	{8'd240,8'd23} : s = 195;
	{8'd240,8'd24} : s = 10;
	{8'd240,8'd25} : s = 74;
	{8'd240,8'd26} : s = 73;
	{8'd240,8'd27} : s = 184;
	{8'd240,8'd28} : s = 70;
	{8'd240,8'd29} : s = 180;
	{8'd240,8'd30} : s = 178;
	{8'd240,8'd31} : s = 314;
	{8'd240,8'd32} : s = 9;
	{8'd240,8'd33} : s = 69;
	{8'd240,8'd34} : s = 67;
	{8'd240,8'd35} : s = 177;
	{8'd240,8'd36} : s = 56;
	{8'd240,8'd37} : s = 172;
	{8'd240,8'd38} : s = 170;
	{8'd240,8'd39} : s = 313;
	{8'd240,8'd40} : s = 52;
	{8'd240,8'd41} : s = 169;
	{8'd240,8'd42} : s = 166;
	{8'd240,8'd43} : s = 310;
	{8'd240,8'd44} : s = 165;
	{8'd240,8'd45} : s = 309;
	{8'd240,8'd46} : s = 307;
	{8'd240,8'd47} : s = 427;
	{8'd240,8'd48} : s = 6;
	{8'd240,8'd49} : s = 50;
	{8'd240,8'd50} : s = 49;
	{8'd240,8'd51} : s = 163;
	{8'd240,8'd52} : s = 44;
	{8'd240,8'd53} : s = 156;
	{8'd240,8'd54} : s = 154;
	{8'd240,8'd55} : s = 302;
	{8'd240,8'd56} : s = 42;
	{8'd240,8'd57} : s = 153;
	{8'd240,8'd58} : s = 150;
	{8'd240,8'd59} : s = 301;
	{8'd240,8'd60} : s = 149;
	{8'd240,8'd61} : s = 299;
	{8'd240,8'd62} : s = 295;
	{8'd240,8'd63} : s = 423;
	{8'd240,8'd64} : s = 41;
	{8'd240,8'd65} : s = 147;
	{8'd240,8'd66} : s = 142;
	{8'd240,8'd67} : s = 286;
	{8'd240,8'd68} : s = 141;
	{8'd240,8'd69} : s = 285;
	{8'd240,8'd70} : s = 283;
	{8'd240,8'd71} : s = 414;
	{8'd240,8'd72} : s = 139;
	{8'd240,8'd73} : s = 279;
	{8'd240,8'd74} : s = 271;
	{8'd240,8'd75} : s = 413;
	{8'd240,8'd76} : s = 248;
	{8'd240,8'd77} : s = 411;
	{8'd240,8'd78} : s = 407;
	{8'd240,8'd79} : s = 491;
	{8'd240,8'd80} : s = 5;
	{8'd240,8'd81} : s = 38;
	{8'd240,8'd82} : s = 37;
	{8'd240,8'd83} : s = 135;
	{8'd240,8'd84} : s = 35;
	{8'd240,8'd85} : s = 120;
	{8'd240,8'd86} : s = 116;
	{8'd240,8'd87} : s = 244;
	{8'd240,8'd88} : s = 28;
	{8'd240,8'd89} : s = 114;
	{8'd240,8'd90} : s = 113;
	{8'd240,8'd91} : s = 242;
	{8'd240,8'd92} : s = 108;
	{8'd240,8'd93} : s = 241;
	{8'd240,8'd94} : s = 236;
	{8'd240,8'd95} : s = 399;
	{8'd240,8'd96} : s = 26;
	{8'd240,8'd97} : s = 106;
	{8'd240,8'd98} : s = 105;
	{8'd240,8'd99} : s = 234;
	{8'd240,8'd100} : s = 102;
	{8'd240,8'd101} : s = 233;
	{8'd240,8'd102} : s = 230;
	{8'd240,8'd103} : s = 380;
	{8'd240,8'd104} : s = 101;
	{8'd240,8'd105} : s = 229;
	{8'd240,8'd106} : s = 227;
	{8'd240,8'd107} : s = 378;
	{8'd240,8'd108} : s = 220;
	{8'd240,8'd109} : s = 377;
	{8'd240,8'd110} : s = 374;
	{8'd240,8'd111} : s = 487;
	{8'd240,8'd112} : s = 25;
	{8'd240,8'd113} : s = 99;
	{8'd240,8'd114} : s = 92;
	{8'd240,8'd115} : s = 218;
	{8'd240,8'd116} : s = 90;
	{8'd240,8'd117} : s = 217;
	{8'd240,8'd118} : s = 214;
	{8'd240,8'd119} : s = 373;
	{8'd240,8'd120} : s = 89;
	{8'd240,8'd121} : s = 213;
	{8'd240,8'd122} : s = 211;
	{8'd240,8'd123} : s = 371;
	{8'd240,8'd124} : s = 206;
	{8'd240,8'd125} : s = 366;
	{8'd240,8'd126} : s = 365;
	{8'd240,8'd127} : s = 478;
	{8'd240,8'd128} : s = 86;
	{8'd240,8'd129} : s = 205;
	{8'd240,8'd130} : s = 203;
	{8'd240,8'd131} : s = 363;
	{8'd240,8'd132} : s = 199;
	{8'd240,8'd133} : s = 359;
	{8'd240,8'd134} : s = 350;
	{8'd240,8'd135} : s = 477;
	{8'd240,8'd136} : s = 188;
	{8'd240,8'd137} : s = 349;
	{8'd240,8'd138} : s = 347;
	{8'd240,8'd139} : s = 475;
	{8'd240,8'd140} : s = 343;
	{8'd240,8'd141} : s = 471;
	{8'd240,8'd142} : s = 463;
	{8'd240,8'd143} : s = 509;
	{8'd240,8'd144} : s = 3;
	{8'd240,8'd145} : s = 22;
	{8'd240,8'd146} : s = 21;
	{8'd240,8'd147} : s = 85;
	{8'd240,8'd148} : s = 19;
	{8'd240,8'd149} : s = 83;
	{8'd240,8'd150} : s = 78;
	{8'd240,8'd151} : s = 186;
	{8'd240,8'd152} : s = 14;
	{8'd240,8'd153} : s = 77;
	{8'd240,8'd154} : s = 75;
	{8'd240,8'd155} : s = 185;
	{8'd240,8'd156} : s = 71;
	{8'd240,8'd157} : s = 182;
	{8'd240,8'd158} : s = 181;
	{8'd240,8'd159} : s = 335;
	{8'd240,8'd160} : s = 13;
	{8'd240,8'd161} : s = 60;
	{8'd240,8'd162} : s = 58;
	{8'd240,8'd163} : s = 179;
	{8'd240,8'd164} : s = 57;
	{8'd240,8'd165} : s = 174;
	{8'd240,8'd166} : s = 173;
	{8'd240,8'd167} : s = 318;
	{8'd240,8'd168} : s = 54;
	{8'd240,8'd169} : s = 171;
	{8'd240,8'd170} : s = 167;
	{8'd240,8'd171} : s = 317;
	{8'd240,8'd172} : s = 158;
	{8'd240,8'd173} : s = 315;
	{8'd240,8'd174} : s = 311;
	{8'd240,8'd175} : s = 446;
	{8'd240,8'd176} : s = 11;
	{8'd240,8'd177} : s = 53;
	{8'd240,8'd178} : s = 51;
	{8'd240,8'd179} : s = 157;
	{8'd240,8'd180} : s = 46;
	{8'd240,8'd181} : s = 155;
	{8'd240,8'd182} : s = 151;
	{8'd240,8'd183} : s = 303;
	{8'd240,8'd184} : s = 45;
	{8'd240,8'd185} : s = 143;
	{8'd240,8'd186} : s = 124;
	{8'd240,8'd187} : s = 287;
	{8'd240,8'd188} : s = 122;
	{8'd240,8'd189} : s = 252;
	{8'd240,8'd190} : s = 250;
	{8'd240,8'd191} : s = 445;
	{8'd240,8'd192} : s = 43;
	{8'd240,8'd193} : s = 121;
	{8'd240,8'd194} : s = 118;
	{8'd240,8'd195} : s = 249;
	{8'd240,8'd196} : s = 117;
	{8'd240,8'd197} : s = 246;
	{8'd240,8'd198} : s = 245;
	{8'd240,8'd199} : s = 443;
	{8'd240,8'd200} : s = 115;
	{8'd240,8'd201} : s = 243;
	{8'd240,8'd202} : s = 238;
	{8'd240,8'd203} : s = 439;
	{8'd240,8'd204} : s = 237;
	{8'd240,8'd205} : s = 431;
	{8'd240,8'd206} : s = 415;
	{8'd240,8'd207} : s = 507;
	{8'd240,8'd208} : s = 7;
	{8'd240,8'd209} : s = 39;
	{8'd240,8'd210} : s = 30;
	{8'd240,8'd211} : s = 110;
	{8'd240,8'd212} : s = 29;
	{8'd240,8'd213} : s = 109;
	{8'd240,8'd214} : s = 107;
	{8'd240,8'd215} : s = 235;
	{8'd240,8'd216} : s = 27;
	{8'd240,8'd217} : s = 103;
	{8'd240,8'd218} : s = 94;
	{8'd240,8'd219} : s = 231;
	{8'd240,8'd220} : s = 93;
	{8'd240,8'd221} : s = 222;
	{8'd240,8'd222} : s = 221;
	{8'd240,8'd223} : s = 382;
	{8'd240,8'd224} : s = 23;
	{8'd240,8'd225} : s = 91;
	{8'd240,8'd226} : s = 87;
	{8'd240,8'd227} : s = 219;
	{8'd240,8'd228} : s = 79;
	{8'd240,8'd229} : s = 215;
	{8'd240,8'd230} : s = 207;
	{8'd240,8'd231} : s = 381;
	{8'd240,8'd232} : s = 62;
	{8'd240,8'd233} : s = 190;
	{8'd240,8'd234} : s = 189;
	{8'd240,8'd235} : s = 379;
	{8'd240,8'd236} : s = 187;
	{8'd240,8'd237} : s = 375;
	{8'd240,8'd238} : s = 367;
	{8'd240,8'd239} : s = 503;
	{8'd240,8'd240} : s = 15;
	{8'd240,8'd241} : s = 61;
	{8'd240,8'd242} : s = 59;
	{8'd240,8'd243} : s = 183;
	{8'd240,8'd244} : s = 55;
	{8'd240,8'd245} : s = 175;
	{8'd240,8'd246} : s = 159;
	{8'd240,8'd247} : s = 351;
	{8'd240,8'd248} : s = 47;
	{8'd240,8'd249} : s = 126;
	{8'd240,8'd250} : s = 125;
	{8'd240,8'd251} : s = 319;
	{8'd240,8'd252} : s = 123;
	{8'd240,8'd253} : s = 254;
	{8'd240,8'd254} : s = 253;
	{8'd240,8'd255} : s = 479;
	{8'd241,8'd0} : s = 333;
	{8'd241,8'd1} : s = 331;
	{8'd241,8'd2} : s = 441;
	{8'd241,8'd3} : s = 327;
	{8'd241,8'd4} : s = 438;
	{8'd241,8'd5} : s = 437;
	{8'd241,8'd6} : s = 501;
	{8'd241,8'd7} : s = 316;
	{8'd241,8'd8} : s = 435;
	{8'd241,8'd9} : s = 430;
	{8'd241,8'd10} : s = 499;
	{8'd241,8'd11} : s = 429;
	{8'd241,8'd12} : s = 494;
	{8'd241,8'd13} : s = 493;
	{8'd241,8'd14} : s = 510;
	{8'd241,8'd15} : s = 1;
	{8'd241,8'd16} : s = 18;
	{8'd241,8'd17} : s = 17;
	{8'd241,8'd18} : s = 82;
	{8'd241,8'd19} : s = 12;
	{8'd241,8'd20} : s = 81;
	{8'd241,8'd21} : s = 76;
	{8'd241,8'd22} : s = 195;
	{8'd241,8'd23} : s = 10;
	{8'd241,8'd24} : s = 74;
	{8'd241,8'd25} : s = 73;
	{8'd241,8'd26} : s = 184;
	{8'd241,8'd27} : s = 70;
	{8'd241,8'd28} : s = 180;
	{8'd241,8'd29} : s = 178;
	{8'd241,8'd30} : s = 314;
	{8'd241,8'd31} : s = 9;
	{8'd241,8'd32} : s = 69;
	{8'd241,8'd33} : s = 67;
	{8'd241,8'd34} : s = 177;
	{8'd241,8'd35} : s = 56;
	{8'd241,8'd36} : s = 172;
	{8'd241,8'd37} : s = 170;
	{8'd241,8'd38} : s = 313;
	{8'd241,8'd39} : s = 52;
	{8'd241,8'd40} : s = 169;
	{8'd241,8'd41} : s = 166;
	{8'd241,8'd42} : s = 310;
	{8'd241,8'd43} : s = 165;
	{8'd241,8'd44} : s = 309;
	{8'd241,8'd45} : s = 307;
	{8'd241,8'd46} : s = 427;
	{8'd241,8'd47} : s = 6;
	{8'd241,8'd48} : s = 50;
	{8'd241,8'd49} : s = 49;
	{8'd241,8'd50} : s = 163;
	{8'd241,8'd51} : s = 44;
	{8'd241,8'd52} : s = 156;
	{8'd241,8'd53} : s = 154;
	{8'd241,8'd54} : s = 302;
	{8'd241,8'd55} : s = 42;
	{8'd241,8'd56} : s = 153;
	{8'd241,8'd57} : s = 150;
	{8'd241,8'd58} : s = 301;
	{8'd241,8'd59} : s = 149;
	{8'd241,8'd60} : s = 299;
	{8'd241,8'd61} : s = 295;
	{8'd241,8'd62} : s = 423;
	{8'd241,8'd63} : s = 41;
	{8'd241,8'd64} : s = 147;
	{8'd241,8'd65} : s = 142;
	{8'd241,8'd66} : s = 286;
	{8'd241,8'd67} : s = 141;
	{8'd241,8'd68} : s = 285;
	{8'd241,8'd69} : s = 283;
	{8'd241,8'd70} : s = 414;
	{8'd241,8'd71} : s = 139;
	{8'd241,8'd72} : s = 279;
	{8'd241,8'd73} : s = 271;
	{8'd241,8'd74} : s = 413;
	{8'd241,8'd75} : s = 248;
	{8'd241,8'd76} : s = 411;
	{8'd241,8'd77} : s = 407;
	{8'd241,8'd78} : s = 491;
	{8'd241,8'd79} : s = 5;
	{8'd241,8'd80} : s = 38;
	{8'd241,8'd81} : s = 37;
	{8'd241,8'd82} : s = 135;
	{8'd241,8'd83} : s = 35;
	{8'd241,8'd84} : s = 120;
	{8'd241,8'd85} : s = 116;
	{8'd241,8'd86} : s = 244;
	{8'd241,8'd87} : s = 28;
	{8'd241,8'd88} : s = 114;
	{8'd241,8'd89} : s = 113;
	{8'd241,8'd90} : s = 242;
	{8'd241,8'd91} : s = 108;
	{8'd241,8'd92} : s = 241;
	{8'd241,8'd93} : s = 236;
	{8'd241,8'd94} : s = 399;
	{8'd241,8'd95} : s = 26;
	{8'd241,8'd96} : s = 106;
	{8'd241,8'd97} : s = 105;
	{8'd241,8'd98} : s = 234;
	{8'd241,8'd99} : s = 102;
	{8'd241,8'd100} : s = 233;
	{8'd241,8'd101} : s = 230;
	{8'd241,8'd102} : s = 380;
	{8'd241,8'd103} : s = 101;
	{8'd241,8'd104} : s = 229;
	{8'd241,8'd105} : s = 227;
	{8'd241,8'd106} : s = 378;
	{8'd241,8'd107} : s = 220;
	{8'd241,8'd108} : s = 377;
	{8'd241,8'd109} : s = 374;
	{8'd241,8'd110} : s = 487;
	{8'd241,8'd111} : s = 25;
	{8'd241,8'd112} : s = 99;
	{8'd241,8'd113} : s = 92;
	{8'd241,8'd114} : s = 218;
	{8'd241,8'd115} : s = 90;
	{8'd241,8'd116} : s = 217;
	{8'd241,8'd117} : s = 214;
	{8'd241,8'd118} : s = 373;
	{8'd241,8'd119} : s = 89;
	{8'd241,8'd120} : s = 213;
	{8'd241,8'd121} : s = 211;
	{8'd241,8'd122} : s = 371;
	{8'd241,8'd123} : s = 206;
	{8'd241,8'd124} : s = 366;
	{8'd241,8'd125} : s = 365;
	{8'd241,8'd126} : s = 478;
	{8'd241,8'd127} : s = 86;
	{8'd241,8'd128} : s = 205;
	{8'd241,8'd129} : s = 203;
	{8'd241,8'd130} : s = 363;
	{8'd241,8'd131} : s = 199;
	{8'd241,8'd132} : s = 359;
	{8'd241,8'd133} : s = 350;
	{8'd241,8'd134} : s = 477;
	{8'd241,8'd135} : s = 188;
	{8'd241,8'd136} : s = 349;
	{8'd241,8'd137} : s = 347;
	{8'd241,8'd138} : s = 475;
	{8'd241,8'd139} : s = 343;
	{8'd241,8'd140} : s = 471;
	{8'd241,8'd141} : s = 463;
	{8'd241,8'd142} : s = 509;
	{8'd241,8'd143} : s = 3;
	{8'd241,8'd144} : s = 22;
	{8'd241,8'd145} : s = 21;
	{8'd241,8'd146} : s = 85;
	{8'd241,8'd147} : s = 19;
	{8'd241,8'd148} : s = 83;
	{8'd241,8'd149} : s = 78;
	{8'd241,8'd150} : s = 186;
	{8'd241,8'd151} : s = 14;
	{8'd241,8'd152} : s = 77;
	{8'd241,8'd153} : s = 75;
	{8'd241,8'd154} : s = 185;
	{8'd241,8'd155} : s = 71;
	{8'd241,8'd156} : s = 182;
	{8'd241,8'd157} : s = 181;
	{8'd241,8'd158} : s = 335;
	{8'd241,8'd159} : s = 13;
	{8'd241,8'd160} : s = 60;
	{8'd241,8'd161} : s = 58;
	{8'd241,8'd162} : s = 179;
	{8'd241,8'd163} : s = 57;
	{8'd241,8'd164} : s = 174;
	{8'd241,8'd165} : s = 173;
	{8'd241,8'd166} : s = 318;
	{8'd241,8'd167} : s = 54;
	{8'd241,8'd168} : s = 171;
	{8'd241,8'd169} : s = 167;
	{8'd241,8'd170} : s = 317;
	{8'd241,8'd171} : s = 158;
	{8'd241,8'd172} : s = 315;
	{8'd241,8'd173} : s = 311;
	{8'd241,8'd174} : s = 446;
	{8'd241,8'd175} : s = 11;
	{8'd241,8'd176} : s = 53;
	{8'd241,8'd177} : s = 51;
	{8'd241,8'd178} : s = 157;
	{8'd241,8'd179} : s = 46;
	{8'd241,8'd180} : s = 155;
	{8'd241,8'd181} : s = 151;
	{8'd241,8'd182} : s = 303;
	{8'd241,8'd183} : s = 45;
	{8'd241,8'd184} : s = 143;
	{8'd241,8'd185} : s = 124;
	{8'd241,8'd186} : s = 287;
	{8'd241,8'd187} : s = 122;
	{8'd241,8'd188} : s = 252;
	{8'd241,8'd189} : s = 250;
	{8'd241,8'd190} : s = 445;
	{8'd241,8'd191} : s = 43;
	{8'd241,8'd192} : s = 121;
	{8'd241,8'd193} : s = 118;
	{8'd241,8'd194} : s = 249;
	{8'd241,8'd195} : s = 117;
	{8'd241,8'd196} : s = 246;
	{8'd241,8'd197} : s = 245;
	{8'd241,8'd198} : s = 443;
	{8'd241,8'd199} : s = 115;
	{8'd241,8'd200} : s = 243;
	{8'd241,8'd201} : s = 238;
	{8'd241,8'd202} : s = 439;
	{8'd241,8'd203} : s = 237;
	{8'd241,8'd204} : s = 431;
	{8'd241,8'd205} : s = 415;
	{8'd241,8'd206} : s = 507;
	{8'd241,8'd207} : s = 7;
	{8'd241,8'd208} : s = 39;
	{8'd241,8'd209} : s = 30;
	{8'd241,8'd210} : s = 110;
	{8'd241,8'd211} : s = 29;
	{8'd241,8'd212} : s = 109;
	{8'd241,8'd213} : s = 107;
	{8'd241,8'd214} : s = 235;
	{8'd241,8'd215} : s = 27;
	{8'd241,8'd216} : s = 103;
	{8'd241,8'd217} : s = 94;
	{8'd241,8'd218} : s = 231;
	{8'd241,8'd219} : s = 93;
	{8'd241,8'd220} : s = 222;
	{8'd241,8'd221} : s = 221;
	{8'd241,8'd222} : s = 382;
	{8'd241,8'd223} : s = 23;
	{8'd241,8'd224} : s = 91;
	{8'd241,8'd225} : s = 87;
	{8'd241,8'd226} : s = 219;
	{8'd241,8'd227} : s = 79;
	{8'd241,8'd228} : s = 215;
	{8'd241,8'd229} : s = 207;
	{8'd241,8'd230} : s = 381;
	{8'd241,8'd231} : s = 62;
	{8'd241,8'd232} : s = 190;
	{8'd241,8'd233} : s = 189;
	{8'd241,8'd234} : s = 379;
	{8'd241,8'd235} : s = 187;
	{8'd241,8'd236} : s = 375;
	{8'd241,8'd237} : s = 367;
	{8'd241,8'd238} : s = 503;
	{8'd241,8'd239} : s = 15;
	{8'd241,8'd240} : s = 61;
	{8'd241,8'd241} : s = 59;
	{8'd241,8'd242} : s = 183;
	{8'd241,8'd243} : s = 55;
	{8'd241,8'd244} : s = 175;
	{8'd241,8'd245} : s = 159;
	{8'd241,8'd246} : s = 351;
	{8'd241,8'd247} : s = 47;
	{8'd241,8'd248} : s = 126;
	{8'd241,8'd249} : s = 125;
	{8'd241,8'd250} : s = 319;
	{8'd241,8'd251} : s = 123;
	{8'd241,8'd252} : s = 254;
	{8'd241,8'd253} : s = 253;
	{8'd241,8'd254} : s = 479;
	{8'd241,8'd255} : s = 31;
	{8'd242,8'd0} : s = 331;
	{8'd242,8'd1} : s = 441;
	{8'd242,8'd2} : s = 327;
	{8'd242,8'd3} : s = 438;
	{8'd242,8'd4} : s = 437;
	{8'd242,8'd5} : s = 501;
	{8'd242,8'd6} : s = 316;
	{8'd242,8'd7} : s = 435;
	{8'd242,8'd8} : s = 430;
	{8'd242,8'd9} : s = 499;
	{8'd242,8'd10} : s = 429;
	{8'd242,8'd11} : s = 494;
	{8'd242,8'd12} : s = 493;
	{8'd242,8'd13} : s = 510;
	{8'd242,8'd14} : s = 1;
	{8'd242,8'd15} : s = 18;
	{8'd242,8'd16} : s = 17;
	{8'd242,8'd17} : s = 82;
	{8'd242,8'd18} : s = 12;
	{8'd242,8'd19} : s = 81;
	{8'd242,8'd20} : s = 76;
	{8'd242,8'd21} : s = 195;
	{8'd242,8'd22} : s = 10;
	{8'd242,8'd23} : s = 74;
	{8'd242,8'd24} : s = 73;
	{8'd242,8'd25} : s = 184;
	{8'd242,8'd26} : s = 70;
	{8'd242,8'd27} : s = 180;
	{8'd242,8'd28} : s = 178;
	{8'd242,8'd29} : s = 314;
	{8'd242,8'd30} : s = 9;
	{8'd242,8'd31} : s = 69;
	{8'd242,8'd32} : s = 67;
	{8'd242,8'd33} : s = 177;
	{8'd242,8'd34} : s = 56;
	{8'd242,8'd35} : s = 172;
	{8'd242,8'd36} : s = 170;
	{8'd242,8'd37} : s = 313;
	{8'd242,8'd38} : s = 52;
	{8'd242,8'd39} : s = 169;
	{8'd242,8'd40} : s = 166;
	{8'd242,8'd41} : s = 310;
	{8'd242,8'd42} : s = 165;
	{8'd242,8'd43} : s = 309;
	{8'd242,8'd44} : s = 307;
	{8'd242,8'd45} : s = 427;
	{8'd242,8'd46} : s = 6;
	{8'd242,8'd47} : s = 50;
	{8'd242,8'd48} : s = 49;
	{8'd242,8'd49} : s = 163;
	{8'd242,8'd50} : s = 44;
	{8'd242,8'd51} : s = 156;
	{8'd242,8'd52} : s = 154;
	{8'd242,8'd53} : s = 302;
	{8'd242,8'd54} : s = 42;
	{8'd242,8'd55} : s = 153;
	{8'd242,8'd56} : s = 150;
	{8'd242,8'd57} : s = 301;
	{8'd242,8'd58} : s = 149;
	{8'd242,8'd59} : s = 299;
	{8'd242,8'd60} : s = 295;
	{8'd242,8'd61} : s = 423;
	{8'd242,8'd62} : s = 41;
	{8'd242,8'd63} : s = 147;
	{8'd242,8'd64} : s = 142;
	{8'd242,8'd65} : s = 286;
	{8'd242,8'd66} : s = 141;
	{8'd242,8'd67} : s = 285;
	{8'd242,8'd68} : s = 283;
	{8'd242,8'd69} : s = 414;
	{8'd242,8'd70} : s = 139;
	{8'd242,8'd71} : s = 279;
	{8'd242,8'd72} : s = 271;
	{8'd242,8'd73} : s = 413;
	{8'd242,8'd74} : s = 248;
	{8'd242,8'd75} : s = 411;
	{8'd242,8'd76} : s = 407;
	{8'd242,8'd77} : s = 491;
	{8'd242,8'd78} : s = 5;
	{8'd242,8'd79} : s = 38;
	{8'd242,8'd80} : s = 37;
	{8'd242,8'd81} : s = 135;
	{8'd242,8'd82} : s = 35;
	{8'd242,8'd83} : s = 120;
	{8'd242,8'd84} : s = 116;
	{8'd242,8'd85} : s = 244;
	{8'd242,8'd86} : s = 28;
	{8'd242,8'd87} : s = 114;
	{8'd242,8'd88} : s = 113;
	{8'd242,8'd89} : s = 242;
	{8'd242,8'd90} : s = 108;
	{8'd242,8'd91} : s = 241;
	{8'd242,8'd92} : s = 236;
	{8'd242,8'd93} : s = 399;
	{8'd242,8'd94} : s = 26;
	{8'd242,8'd95} : s = 106;
	{8'd242,8'd96} : s = 105;
	{8'd242,8'd97} : s = 234;
	{8'd242,8'd98} : s = 102;
	{8'd242,8'd99} : s = 233;
	{8'd242,8'd100} : s = 230;
	{8'd242,8'd101} : s = 380;
	{8'd242,8'd102} : s = 101;
	{8'd242,8'd103} : s = 229;
	{8'd242,8'd104} : s = 227;
	{8'd242,8'd105} : s = 378;
	{8'd242,8'd106} : s = 220;
	{8'd242,8'd107} : s = 377;
	{8'd242,8'd108} : s = 374;
	{8'd242,8'd109} : s = 487;
	{8'd242,8'd110} : s = 25;
	{8'd242,8'd111} : s = 99;
	{8'd242,8'd112} : s = 92;
	{8'd242,8'd113} : s = 218;
	{8'd242,8'd114} : s = 90;
	{8'd242,8'd115} : s = 217;
	{8'd242,8'd116} : s = 214;
	{8'd242,8'd117} : s = 373;
	{8'd242,8'd118} : s = 89;
	{8'd242,8'd119} : s = 213;
	{8'd242,8'd120} : s = 211;
	{8'd242,8'd121} : s = 371;
	{8'd242,8'd122} : s = 206;
	{8'd242,8'd123} : s = 366;
	{8'd242,8'd124} : s = 365;
	{8'd242,8'd125} : s = 478;
	{8'd242,8'd126} : s = 86;
	{8'd242,8'd127} : s = 205;
	{8'd242,8'd128} : s = 203;
	{8'd242,8'd129} : s = 363;
	{8'd242,8'd130} : s = 199;
	{8'd242,8'd131} : s = 359;
	{8'd242,8'd132} : s = 350;
	{8'd242,8'd133} : s = 477;
	{8'd242,8'd134} : s = 188;
	{8'd242,8'd135} : s = 349;
	{8'd242,8'd136} : s = 347;
	{8'd242,8'd137} : s = 475;
	{8'd242,8'd138} : s = 343;
	{8'd242,8'd139} : s = 471;
	{8'd242,8'd140} : s = 463;
	{8'd242,8'd141} : s = 509;
	{8'd242,8'd142} : s = 3;
	{8'd242,8'd143} : s = 22;
	{8'd242,8'd144} : s = 21;
	{8'd242,8'd145} : s = 85;
	{8'd242,8'd146} : s = 19;
	{8'd242,8'd147} : s = 83;
	{8'd242,8'd148} : s = 78;
	{8'd242,8'd149} : s = 186;
	{8'd242,8'd150} : s = 14;
	{8'd242,8'd151} : s = 77;
	{8'd242,8'd152} : s = 75;
	{8'd242,8'd153} : s = 185;
	{8'd242,8'd154} : s = 71;
	{8'd242,8'd155} : s = 182;
	{8'd242,8'd156} : s = 181;
	{8'd242,8'd157} : s = 335;
	{8'd242,8'd158} : s = 13;
	{8'd242,8'd159} : s = 60;
	{8'd242,8'd160} : s = 58;
	{8'd242,8'd161} : s = 179;
	{8'd242,8'd162} : s = 57;
	{8'd242,8'd163} : s = 174;
	{8'd242,8'd164} : s = 173;
	{8'd242,8'd165} : s = 318;
	{8'd242,8'd166} : s = 54;
	{8'd242,8'd167} : s = 171;
	{8'd242,8'd168} : s = 167;
	{8'd242,8'd169} : s = 317;
	{8'd242,8'd170} : s = 158;
	{8'd242,8'd171} : s = 315;
	{8'd242,8'd172} : s = 311;
	{8'd242,8'd173} : s = 446;
	{8'd242,8'd174} : s = 11;
	{8'd242,8'd175} : s = 53;
	{8'd242,8'd176} : s = 51;
	{8'd242,8'd177} : s = 157;
	{8'd242,8'd178} : s = 46;
	{8'd242,8'd179} : s = 155;
	{8'd242,8'd180} : s = 151;
	{8'd242,8'd181} : s = 303;
	{8'd242,8'd182} : s = 45;
	{8'd242,8'd183} : s = 143;
	{8'd242,8'd184} : s = 124;
	{8'd242,8'd185} : s = 287;
	{8'd242,8'd186} : s = 122;
	{8'd242,8'd187} : s = 252;
	{8'd242,8'd188} : s = 250;
	{8'd242,8'd189} : s = 445;
	{8'd242,8'd190} : s = 43;
	{8'd242,8'd191} : s = 121;
	{8'd242,8'd192} : s = 118;
	{8'd242,8'd193} : s = 249;
	{8'd242,8'd194} : s = 117;
	{8'd242,8'd195} : s = 246;
	{8'd242,8'd196} : s = 245;
	{8'd242,8'd197} : s = 443;
	{8'd242,8'd198} : s = 115;
	{8'd242,8'd199} : s = 243;
	{8'd242,8'd200} : s = 238;
	{8'd242,8'd201} : s = 439;
	{8'd242,8'd202} : s = 237;
	{8'd242,8'd203} : s = 431;
	{8'd242,8'd204} : s = 415;
	{8'd242,8'd205} : s = 507;
	{8'd242,8'd206} : s = 7;
	{8'd242,8'd207} : s = 39;
	{8'd242,8'd208} : s = 30;
	{8'd242,8'd209} : s = 110;
	{8'd242,8'd210} : s = 29;
	{8'd242,8'd211} : s = 109;
	{8'd242,8'd212} : s = 107;
	{8'd242,8'd213} : s = 235;
	{8'd242,8'd214} : s = 27;
	{8'd242,8'd215} : s = 103;
	{8'd242,8'd216} : s = 94;
	{8'd242,8'd217} : s = 231;
	{8'd242,8'd218} : s = 93;
	{8'd242,8'd219} : s = 222;
	{8'd242,8'd220} : s = 221;
	{8'd242,8'd221} : s = 382;
	{8'd242,8'd222} : s = 23;
	{8'd242,8'd223} : s = 91;
	{8'd242,8'd224} : s = 87;
	{8'd242,8'd225} : s = 219;
	{8'd242,8'd226} : s = 79;
	{8'd242,8'd227} : s = 215;
	{8'd242,8'd228} : s = 207;
	{8'd242,8'd229} : s = 381;
	{8'd242,8'd230} : s = 62;
	{8'd242,8'd231} : s = 190;
	{8'd242,8'd232} : s = 189;
	{8'd242,8'd233} : s = 379;
	{8'd242,8'd234} : s = 187;
	{8'd242,8'd235} : s = 375;
	{8'd242,8'd236} : s = 367;
	{8'd242,8'd237} : s = 503;
	{8'd242,8'd238} : s = 15;
	{8'd242,8'd239} : s = 61;
	{8'd242,8'd240} : s = 59;
	{8'd242,8'd241} : s = 183;
	{8'd242,8'd242} : s = 55;
	{8'd242,8'd243} : s = 175;
	{8'd242,8'd244} : s = 159;
	{8'd242,8'd245} : s = 351;
	{8'd242,8'd246} : s = 47;
	{8'd242,8'd247} : s = 126;
	{8'd242,8'd248} : s = 125;
	{8'd242,8'd249} : s = 319;
	{8'd242,8'd250} : s = 123;
	{8'd242,8'd251} : s = 254;
	{8'd242,8'd252} : s = 253;
	{8'd242,8'd253} : s = 479;
	{8'd242,8'd254} : s = 31;
	{8'd242,8'd255} : s = 119;
	{8'd243,8'd0} : s = 441;
	{8'd243,8'd1} : s = 327;
	{8'd243,8'd2} : s = 438;
	{8'd243,8'd3} : s = 437;
	{8'd243,8'd4} : s = 501;
	{8'd243,8'd5} : s = 316;
	{8'd243,8'd6} : s = 435;
	{8'd243,8'd7} : s = 430;
	{8'd243,8'd8} : s = 499;
	{8'd243,8'd9} : s = 429;
	{8'd243,8'd10} : s = 494;
	{8'd243,8'd11} : s = 493;
	{8'd243,8'd12} : s = 510;
	{8'd243,8'd13} : s = 1;
	{8'd243,8'd14} : s = 18;
	{8'd243,8'd15} : s = 17;
	{8'd243,8'd16} : s = 82;
	{8'd243,8'd17} : s = 12;
	{8'd243,8'd18} : s = 81;
	{8'd243,8'd19} : s = 76;
	{8'd243,8'd20} : s = 195;
	{8'd243,8'd21} : s = 10;
	{8'd243,8'd22} : s = 74;
	{8'd243,8'd23} : s = 73;
	{8'd243,8'd24} : s = 184;
	{8'd243,8'd25} : s = 70;
	{8'd243,8'd26} : s = 180;
	{8'd243,8'd27} : s = 178;
	{8'd243,8'd28} : s = 314;
	{8'd243,8'd29} : s = 9;
	{8'd243,8'd30} : s = 69;
	{8'd243,8'd31} : s = 67;
	{8'd243,8'd32} : s = 177;
	{8'd243,8'd33} : s = 56;
	{8'd243,8'd34} : s = 172;
	{8'd243,8'd35} : s = 170;
	{8'd243,8'd36} : s = 313;
	{8'd243,8'd37} : s = 52;
	{8'd243,8'd38} : s = 169;
	{8'd243,8'd39} : s = 166;
	{8'd243,8'd40} : s = 310;
	{8'd243,8'd41} : s = 165;
	{8'd243,8'd42} : s = 309;
	{8'd243,8'd43} : s = 307;
	{8'd243,8'd44} : s = 427;
	{8'd243,8'd45} : s = 6;
	{8'd243,8'd46} : s = 50;
	{8'd243,8'd47} : s = 49;
	{8'd243,8'd48} : s = 163;
	{8'd243,8'd49} : s = 44;
	{8'd243,8'd50} : s = 156;
	{8'd243,8'd51} : s = 154;
	{8'd243,8'd52} : s = 302;
	{8'd243,8'd53} : s = 42;
	{8'd243,8'd54} : s = 153;
	{8'd243,8'd55} : s = 150;
	{8'd243,8'd56} : s = 301;
	{8'd243,8'd57} : s = 149;
	{8'd243,8'd58} : s = 299;
	{8'd243,8'd59} : s = 295;
	{8'd243,8'd60} : s = 423;
	{8'd243,8'd61} : s = 41;
	{8'd243,8'd62} : s = 147;
	{8'd243,8'd63} : s = 142;
	{8'd243,8'd64} : s = 286;
	{8'd243,8'd65} : s = 141;
	{8'd243,8'd66} : s = 285;
	{8'd243,8'd67} : s = 283;
	{8'd243,8'd68} : s = 414;
	{8'd243,8'd69} : s = 139;
	{8'd243,8'd70} : s = 279;
	{8'd243,8'd71} : s = 271;
	{8'd243,8'd72} : s = 413;
	{8'd243,8'd73} : s = 248;
	{8'd243,8'd74} : s = 411;
	{8'd243,8'd75} : s = 407;
	{8'd243,8'd76} : s = 491;
	{8'd243,8'd77} : s = 5;
	{8'd243,8'd78} : s = 38;
	{8'd243,8'd79} : s = 37;
	{8'd243,8'd80} : s = 135;
	{8'd243,8'd81} : s = 35;
	{8'd243,8'd82} : s = 120;
	{8'd243,8'd83} : s = 116;
	{8'd243,8'd84} : s = 244;
	{8'd243,8'd85} : s = 28;
	{8'd243,8'd86} : s = 114;
	{8'd243,8'd87} : s = 113;
	{8'd243,8'd88} : s = 242;
	{8'd243,8'd89} : s = 108;
	{8'd243,8'd90} : s = 241;
	{8'd243,8'd91} : s = 236;
	{8'd243,8'd92} : s = 399;
	{8'd243,8'd93} : s = 26;
	{8'd243,8'd94} : s = 106;
	{8'd243,8'd95} : s = 105;
	{8'd243,8'd96} : s = 234;
	{8'd243,8'd97} : s = 102;
	{8'd243,8'd98} : s = 233;
	{8'd243,8'd99} : s = 230;
	{8'd243,8'd100} : s = 380;
	{8'd243,8'd101} : s = 101;
	{8'd243,8'd102} : s = 229;
	{8'd243,8'd103} : s = 227;
	{8'd243,8'd104} : s = 378;
	{8'd243,8'd105} : s = 220;
	{8'd243,8'd106} : s = 377;
	{8'd243,8'd107} : s = 374;
	{8'd243,8'd108} : s = 487;
	{8'd243,8'd109} : s = 25;
	{8'd243,8'd110} : s = 99;
	{8'd243,8'd111} : s = 92;
	{8'd243,8'd112} : s = 218;
	{8'd243,8'd113} : s = 90;
	{8'd243,8'd114} : s = 217;
	{8'd243,8'd115} : s = 214;
	{8'd243,8'd116} : s = 373;
	{8'd243,8'd117} : s = 89;
	{8'd243,8'd118} : s = 213;
	{8'd243,8'd119} : s = 211;
	{8'd243,8'd120} : s = 371;
	{8'd243,8'd121} : s = 206;
	{8'd243,8'd122} : s = 366;
	{8'd243,8'd123} : s = 365;
	{8'd243,8'd124} : s = 478;
	{8'd243,8'd125} : s = 86;
	{8'd243,8'd126} : s = 205;
	{8'd243,8'd127} : s = 203;
	{8'd243,8'd128} : s = 363;
	{8'd243,8'd129} : s = 199;
	{8'd243,8'd130} : s = 359;
	{8'd243,8'd131} : s = 350;
	{8'd243,8'd132} : s = 477;
	{8'd243,8'd133} : s = 188;
	{8'd243,8'd134} : s = 349;
	{8'd243,8'd135} : s = 347;
	{8'd243,8'd136} : s = 475;
	{8'd243,8'd137} : s = 343;
	{8'd243,8'd138} : s = 471;
	{8'd243,8'd139} : s = 463;
	{8'd243,8'd140} : s = 509;
	{8'd243,8'd141} : s = 3;
	{8'd243,8'd142} : s = 22;
	{8'd243,8'd143} : s = 21;
	{8'd243,8'd144} : s = 85;
	{8'd243,8'd145} : s = 19;
	{8'd243,8'd146} : s = 83;
	{8'd243,8'd147} : s = 78;
	{8'd243,8'd148} : s = 186;
	{8'd243,8'd149} : s = 14;
	{8'd243,8'd150} : s = 77;
	{8'd243,8'd151} : s = 75;
	{8'd243,8'd152} : s = 185;
	{8'd243,8'd153} : s = 71;
	{8'd243,8'd154} : s = 182;
	{8'd243,8'd155} : s = 181;
	{8'd243,8'd156} : s = 335;
	{8'd243,8'd157} : s = 13;
	{8'd243,8'd158} : s = 60;
	{8'd243,8'd159} : s = 58;
	{8'd243,8'd160} : s = 179;
	{8'd243,8'd161} : s = 57;
	{8'd243,8'd162} : s = 174;
	{8'd243,8'd163} : s = 173;
	{8'd243,8'd164} : s = 318;
	{8'd243,8'd165} : s = 54;
	{8'd243,8'd166} : s = 171;
	{8'd243,8'd167} : s = 167;
	{8'd243,8'd168} : s = 317;
	{8'd243,8'd169} : s = 158;
	{8'd243,8'd170} : s = 315;
	{8'd243,8'd171} : s = 311;
	{8'd243,8'd172} : s = 446;
	{8'd243,8'd173} : s = 11;
	{8'd243,8'd174} : s = 53;
	{8'd243,8'd175} : s = 51;
	{8'd243,8'd176} : s = 157;
	{8'd243,8'd177} : s = 46;
	{8'd243,8'd178} : s = 155;
	{8'd243,8'd179} : s = 151;
	{8'd243,8'd180} : s = 303;
	{8'd243,8'd181} : s = 45;
	{8'd243,8'd182} : s = 143;
	{8'd243,8'd183} : s = 124;
	{8'd243,8'd184} : s = 287;
	{8'd243,8'd185} : s = 122;
	{8'd243,8'd186} : s = 252;
	{8'd243,8'd187} : s = 250;
	{8'd243,8'd188} : s = 445;
	{8'd243,8'd189} : s = 43;
	{8'd243,8'd190} : s = 121;
	{8'd243,8'd191} : s = 118;
	{8'd243,8'd192} : s = 249;
	{8'd243,8'd193} : s = 117;
	{8'd243,8'd194} : s = 246;
	{8'd243,8'd195} : s = 245;
	{8'd243,8'd196} : s = 443;
	{8'd243,8'd197} : s = 115;
	{8'd243,8'd198} : s = 243;
	{8'd243,8'd199} : s = 238;
	{8'd243,8'd200} : s = 439;
	{8'd243,8'd201} : s = 237;
	{8'd243,8'd202} : s = 431;
	{8'd243,8'd203} : s = 415;
	{8'd243,8'd204} : s = 507;
	{8'd243,8'd205} : s = 7;
	{8'd243,8'd206} : s = 39;
	{8'd243,8'd207} : s = 30;
	{8'd243,8'd208} : s = 110;
	{8'd243,8'd209} : s = 29;
	{8'd243,8'd210} : s = 109;
	{8'd243,8'd211} : s = 107;
	{8'd243,8'd212} : s = 235;
	{8'd243,8'd213} : s = 27;
	{8'd243,8'd214} : s = 103;
	{8'd243,8'd215} : s = 94;
	{8'd243,8'd216} : s = 231;
	{8'd243,8'd217} : s = 93;
	{8'd243,8'd218} : s = 222;
	{8'd243,8'd219} : s = 221;
	{8'd243,8'd220} : s = 382;
	{8'd243,8'd221} : s = 23;
	{8'd243,8'd222} : s = 91;
	{8'd243,8'd223} : s = 87;
	{8'd243,8'd224} : s = 219;
	{8'd243,8'd225} : s = 79;
	{8'd243,8'd226} : s = 215;
	{8'd243,8'd227} : s = 207;
	{8'd243,8'd228} : s = 381;
	{8'd243,8'd229} : s = 62;
	{8'd243,8'd230} : s = 190;
	{8'd243,8'd231} : s = 189;
	{8'd243,8'd232} : s = 379;
	{8'd243,8'd233} : s = 187;
	{8'd243,8'd234} : s = 375;
	{8'd243,8'd235} : s = 367;
	{8'd243,8'd236} : s = 503;
	{8'd243,8'd237} : s = 15;
	{8'd243,8'd238} : s = 61;
	{8'd243,8'd239} : s = 59;
	{8'd243,8'd240} : s = 183;
	{8'd243,8'd241} : s = 55;
	{8'd243,8'd242} : s = 175;
	{8'd243,8'd243} : s = 159;
	{8'd243,8'd244} : s = 351;
	{8'd243,8'd245} : s = 47;
	{8'd243,8'd246} : s = 126;
	{8'd243,8'd247} : s = 125;
	{8'd243,8'd248} : s = 319;
	{8'd243,8'd249} : s = 123;
	{8'd243,8'd250} : s = 254;
	{8'd243,8'd251} : s = 253;
	{8'd243,8'd252} : s = 479;
	{8'd243,8'd253} : s = 31;
	{8'd243,8'd254} : s = 119;
	{8'd243,8'd255} : s = 111;
	{8'd244,8'd0} : s = 327;
	{8'd244,8'd1} : s = 438;
	{8'd244,8'd2} : s = 437;
	{8'd244,8'd3} : s = 501;
	{8'd244,8'd4} : s = 316;
	{8'd244,8'd5} : s = 435;
	{8'd244,8'd6} : s = 430;
	{8'd244,8'd7} : s = 499;
	{8'd244,8'd8} : s = 429;
	{8'd244,8'd9} : s = 494;
	{8'd244,8'd10} : s = 493;
	{8'd244,8'd11} : s = 510;
	{8'd244,8'd12} : s = 1;
	{8'd244,8'd13} : s = 18;
	{8'd244,8'd14} : s = 17;
	{8'd244,8'd15} : s = 82;
	{8'd244,8'd16} : s = 12;
	{8'd244,8'd17} : s = 81;
	{8'd244,8'd18} : s = 76;
	{8'd244,8'd19} : s = 195;
	{8'd244,8'd20} : s = 10;
	{8'd244,8'd21} : s = 74;
	{8'd244,8'd22} : s = 73;
	{8'd244,8'd23} : s = 184;
	{8'd244,8'd24} : s = 70;
	{8'd244,8'd25} : s = 180;
	{8'd244,8'd26} : s = 178;
	{8'd244,8'd27} : s = 314;
	{8'd244,8'd28} : s = 9;
	{8'd244,8'd29} : s = 69;
	{8'd244,8'd30} : s = 67;
	{8'd244,8'd31} : s = 177;
	{8'd244,8'd32} : s = 56;
	{8'd244,8'd33} : s = 172;
	{8'd244,8'd34} : s = 170;
	{8'd244,8'd35} : s = 313;
	{8'd244,8'd36} : s = 52;
	{8'd244,8'd37} : s = 169;
	{8'd244,8'd38} : s = 166;
	{8'd244,8'd39} : s = 310;
	{8'd244,8'd40} : s = 165;
	{8'd244,8'd41} : s = 309;
	{8'd244,8'd42} : s = 307;
	{8'd244,8'd43} : s = 427;
	{8'd244,8'd44} : s = 6;
	{8'd244,8'd45} : s = 50;
	{8'd244,8'd46} : s = 49;
	{8'd244,8'd47} : s = 163;
	{8'd244,8'd48} : s = 44;
	{8'd244,8'd49} : s = 156;
	{8'd244,8'd50} : s = 154;
	{8'd244,8'd51} : s = 302;
	{8'd244,8'd52} : s = 42;
	{8'd244,8'd53} : s = 153;
	{8'd244,8'd54} : s = 150;
	{8'd244,8'd55} : s = 301;
	{8'd244,8'd56} : s = 149;
	{8'd244,8'd57} : s = 299;
	{8'd244,8'd58} : s = 295;
	{8'd244,8'd59} : s = 423;
	{8'd244,8'd60} : s = 41;
	{8'd244,8'd61} : s = 147;
	{8'd244,8'd62} : s = 142;
	{8'd244,8'd63} : s = 286;
	{8'd244,8'd64} : s = 141;
	{8'd244,8'd65} : s = 285;
	{8'd244,8'd66} : s = 283;
	{8'd244,8'd67} : s = 414;
	{8'd244,8'd68} : s = 139;
	{8'd244,8'd69} : s = 279;
	{8'd244,8'd70} : s = 271;
	{8'd244,8'd71} : s = 413;
	{8'd244,8'd72} : s = 248;
	{8'd244,8'd73} : s = 411;
	{8'd244,8'd74} : s = 407;
	{8'd244,8'd75} : s = 491;
	{8'd244,8'd76} : s = 5;
	{8'd244,8'd77} : s = 38;
	{8'd244,8'd78} : s = 37;
	{8'd244,8'd79} : s = 135;
	{8'd244,8'd80} : s = 35;
	{8'd244,8'd81} : s = 120;
	{8'd244,8'd82} : s = 116;
	{8'd244,8'd83} : s = 244;
	{8'd244,8'd84} : s = 28;
	{8'd244,8'd85} : s = 114;
	{8'd244,8'd86} : s = 113;
	{8'd244,8'd87} : s = 242;
	{8'd244,8'd88} : s = 108;
	{8'd244,8'd89} : s = 241;
	{8'd244,8'd90} : s = 236;
	{8'd244,8'd91} : s = 399;
	{8'd244,8'd92} : s = 26;
	{8'd244,8'd93} : s = 106;
	{8'd244,8'd94} : s = 105;
	{8'd244,8'd95} : s = 234;
	{8'd244,8'd96} : s = 102;
	{8'd244,8'd97} : s = 233;
	{8'd244,8'd98} : s = 230;
	{8'd244,8'd99} : s = 380;
	{8'd244,8'd100} : s = 101;
	{8'd244,8'd101} : s = 229;
	{8'd244,8'd102} : s = 227;
	{8'd244,8'd103} : s = 378;
	{8'd244,8'd104} : s = 220;
	{8'd244,8'd105} : s = 377;
	{8'd244,8'd106} : s = 374;
	{8'd244,8'd107} : s = 487;
	{8'd244,8'd108} : s = 25;
	{8'd244,8'd109} : s = 99;
	{8'd244,8'd110} : s = 92;
	{8'd244,8'd111} : s = 218;
	{8'd244,8'd112} : s = 90;
	{8'd244,8'd113} : s = 217;
	{8'd244,8'd114} : s = 214;
	{8'd244,8'd115} : s = 373;
	{8'd244,8'd116} : s = 89;
	{8'd244,8'd117} : s = 213;
	{8'd244,8'd118} : s = 211;
	{8'd244,8'd119} : s = 371;
	{8'd244,8'd120} : s = 206;
	{8'd244,8'd121} : s = 366;
	{8'd244,8'd122} : s = 365;
	{8'd244,8'd123} : s = 478;
	{8'd244,8'd124} : s = 86;
	{8'd244,8'd125} : s = 205;
	{8'd244,8'd126} : s = 203;
	{8'd244,8'd127} : s = 363;
	{8'd244,8'd128} : s = 199;
	{8'd244,8'd129} : s = 359;
	{8'd244,8'd130} : s = 350;
	{8'd244,8'd131} : s = 477;
	{8'd244,8'd132} : s = 188;
	{8'd244,8'd133} : s = 349;
	{8'd244,8'd134} : s = 347;
	{8'd244,8'd135} : s = 475;
	{8'd244,8'd136} : s = 343;
	{8'd244,8'd137} : s = 471;
	{8'd244,8'd138} : s = 463;
	{8'd244,8'd139} : s = 509;
	{8'd244,8'd140} : s = 3;
	{8'd244,8'd141} : s = 22;
	{8'd244,8'd142} : s = 21;
	{8'd244,8'd143} : s = 85;
	{8'd244,8'd144} : s = 19;
	{8'd244,8'd145} : s = 83;
	{8'd244,8'd146} : s = 78;
	{8'd244,8'd147} : s = 186;
	{8'd244,8'd148} : s = 14;
	{8'd244,8'd149} : s = 77;
	{8'd244,8'd150} : s = 75;
	{8'd244,8'd151} : s = 185;
	{8'd244,8'd152} : s = 71;
	{8'd244,8'd153} : s = 182;
	{8'd244,8'd154} : s = 181;
	{8'd244,8'd155} : s = 335;
	{8'd244,8'd156} : s = 13;
	{8'd244,8'd157} : s = 60;
	{8'd244,8'd158} : s = 58;
	{8'd244,8'd159} : s = 179;
	{8'd244,8'd160} : s = 57;
	{8'd244,8'd161} : s = 174;
	{8'd244,8'd162} : s = 173;
	{8'd244,8'd163} : s = 318;
	{8'd244,8'd164} : s = 54;
	{8'd244,8'd165} : s = 171;
	{8'd244,8'd166} : s = 167;
	{8'd244,8'd167} : s = 317;
	{8'd244,8'd168} : s = 158;
	{8'd244,8'd169} : s = 315;
	{8'd244,8'd170} : s = 311;
	{8'd244,8'd171} : s = 446;
	{8'd244,8'd172} : s = 11;
	{8'd244,8'd173} : s = 53;
	{8'd244,8'd174} : s = 51;
	{8'd244,8'd175} : s = 157;
	{8'd244,8'd176} : s = 46;
	{8'd244,8'd177} : s = 155;
	{8'd244,8'd178} : s = 151;
	{8'd244,8'd179} : s = 303;
	{8'd244,8'd180} : s = 45;
	{8'd244,8'd181} : s = 143;
	{8'd244,8'd182} : s = 124;
	{8'd244,8'd183} : s = 287;
	{8'd244,8'd184} : s = 122;
	{8'd244,8'd185} : s = 252;
	{8'd244,8'd186} : s = 250;
	{8'd244,8'd187} : s = 445;
	{8'd244,8'd188} : s = 43;
	{8'd244,8'd189} : s = 121;
	{8'd244,8'd190} : s = 118;
	{8'd244,8'd191} : s = 249;
	{8'd244,8'd192} : s = 117;
	{8'd244,8'd193} : s = 246;
	{8'd244,8'd194} : s = 245;
	{8'd244,8'd195} : s = 443;
	{8'd244,8'd196} : s = 115;
	{8'd244,8'd197} : s = 243;
	{8'd244,8'd198} : s = 238;
	{8'd244,8'd199} : s = 439;
	{8'd244,8'd200} : s = 237;
	{8'd244,8'd201} : s = 431;
	{8'd244,8'd202} : s = 415;
	{8'd244,8'd203} : s = 507;
	{8'd244,8'd204} : s = 7;
	{8'd244,8'd205} : s = 39;
	{8'd244,8'd206} : s = 30;
	{8'd244,8'd207} : s = 110;
	{8'd244,8'd208} : s = 29;
	{8'd244,8'd209} : s = 109;
	{8'd244,8'd210} : s = 107;
	{8'd244,8'd211} : s = 235;
	{8'd244,8'd212} : s = 27;
	{8'd244,8'd213} : s = 103;
	{8'd244,8'd214} : s = 94;
	{8'd244,8'd215} : s = 231;
	{8'd244,8'd216} : s = 93;
	{8'd244,8'd217} : s = 222;
	{8'd244,8'd218} : s = 221;
	{8'd244,8'd219} : s = 382;
	{8'd244,8'd220} : s = 23;
	{8'd244,8'd221} : s = 91;
	{8'd244,8'd222} : s = 87;
	{8'd244,8'd223} : s = 219;
	{8'd244,8'd224} : s = 79;
	{8'd244,8'd225} : s = 215;
	{8'd244,8'd226} : s = 207;
	{8'd244,8'd227} : s = 381;
	{8'd244,8'd228} : s = 62;
	{8'd244,8'd229} : s = 190;
	{8'd244,8'd230} : s = 189;
	{8'd244,8'd231} : s = 379;
	{8'd244,8'd232} : s = 187;
	{8'd244,8'd233} : s = 375;
	{8'd244,8'd234} : s = 367;
	{8'd244,8'd235} : s = 503;
	{8'd244,8'd236} : s = 15;
	{8'd244,8'd237} : s = 61;
	{8'd244,8'd238} : s = 59;
	{8'd244,8'd239} : s = 183;
	{8'd244,8'd240} : s = 55;
	{8'd244,8'd241} : s = 175;
	{8'd244,8'd242} : s = 159;
	{8'd244,8'd243} : s = 351;
	{8'd244,8'd244} : s = 47;
	{8'd244,8'd245} : s = 126;
	{8'd244,8'd246} : s = 125;
	{8'd244,8'd247} : s = 319;
	{8'd244,8'd248} : s = 123;
	{8'd244,8'd249} : s = 254;
	{8'd244,8'd250} : s = 253;
	{8'd244,8'd251} : s = 479;
	{8'd244,8'd252} : s = 31;
	{8'd244,8'd253} : s = 119;
	{8'd244,8'd254} : s = 111;
	{8'd244,8'd255} : s = 251;
	{8'd245,8'd0} : s = 438;
	{8'd245,8'd1} : s = 437;
	{8'd245,8'd2} : s = 501;
	{8'd245,8'd3} : s = 316;
	{8'd245,8'd4} : s = 435;
	{8'd245,8'd5} : s = 430;
	{8'd245,8'd6} : s = 499;
	{8'd245,8'd7} : s = 429;
	{8'd245,8'd8} : s = 494;
	{8'd245,8'd9} : s = 493;
	{8'd245,8'd10} : s = 510;
	{8'd245,8'd11} : s = 1;
	{8'd245,8'd12} : s = 18;
	{8'd245,8'd13} : s = 17;
	{8'd245,8'd14} : s = 82;
	{8'd245,8'd15} : s = 12;
	{8'd245,8'd16} : s = 81;
	{8'd245,8'd17} : s = 76;
	{8'd245,8'd18} : s = 195;
	{8'd245,8'd19} : s = 10;
	{8'd245,8'd20} : s = 74;
	{8'd245,8'd21} : s = 73;
	{8'd245,8'd22} : s = 184;
	{8'd245,8'd23} : s = 70;
	{8'd245,8'd24} : s = 180;
	{8'd245,8'd25} : s = 178;
	{8'd245,8'd26} : s = 314;
	{8'd245,8'd27} : s = 9;
	{8'd245,8'd28} : s = 69;
	{8'd245,8'd29} : s = 67;
	{8'd245,8'd30} : s = 177;
	{8'd245,8'd31} : s = 56;
	{8'd245,8'd32} : s = 172;
	{8'd245,8'd33} : s = 170;
	{8'd245,8'd34} : s = 313;
	{8'd245,8'd35} : s = 52;
	{8'd245,8'd36} : s = 169;
	{8'd245,8'd37} : s = 166;
	{8'd245,8'd38} : s = 310;
	{8'd245,8'd39} : s = 165;
	{8'd245,8'd40} : s = 309;
	{8'd245,8'd41} : s = 307;
	{8'd245,8'd42} : s = 427;
	{8'd245,8'd43} : s = 6;
	{8'd245,8'd44} : s = 50;
	{8'd245,8'd45} : s = 49;
	{8'd245,8'd46} : s = 163;
	{8'd245,8'd47} : s = 44;
	{8'd245,8'd48} : s = 156;
	{8'd245,8'd49} : s = 154;
	{8'd245,8'd50} : s = 302;
	{8'd245,8'd51} : s = 42;
	{8'd245,8'd52} : s = 153;
	{8'd245,8'd53} : s = 150;
	{8'd245,8'd54} : s = 301;
	{8'd245,8'd55} : s = 149;
	{8'd245,8'd56} : s = 299;
	{8'd245,8'd57} : s = 295;
	{8'd245,8'd58} : s = 423;
	{8'd245,8'd59} : s = 41;
	{8'd245,8'd60} : s = 147;
	{8'd245,8'd61} : s = 142;
	{8'd245,8'd62} : s = 286;
	{8'd245,8'd63} : s = 141;
	{8'd245,8'd64} : s = 285;
	{8'd245,8'd65} : s = 283;
	{8'd245,8'd66} : s = 414;
	{8'd245,8'd67} : s = 139;
	{8'd245,8'd68} : s = 279;
	{8'd245,8'd69} : s = 271;
	{8'd245,8'd70} : s = 413;
	{8'd245,8'd71} : s = 248;
	{8'd245,8'd72} : s = 411;
	{8'd245,8'd73} : s = 407;
	{8'd245,8'd74} : s = 491;
	{8'd245,8'd75} : s = 5;
	{8'd245,8'd76} : s = 38;
	{8'd245,8'd77} : s = 37;
	{8'd245,8'd78} : s = 135;
	{8'd245,8'd79} : s = 35;
	{8'd245,8'd80} : s = 120;
	{8'd245,8'd81} : s = 116;
	{8'd245,8'd82} : s = 244;
	{8'd245,8'd83} : s = 28;
	{8'd245,8'd84} : s = 114;
	{8'd245,8'd85} : s = 113;
	{8'd245,8'd86} : s = 242;
	{8'd245,8'd87} : s = 108;
	{8'd245,8'd88} : s = 241;
	{8'd245,8'd89} : s = 236;
	{8'd245,8'd90} : s = 399;
	{8'd245,8'd91} : s = 26;
	{8'd245,8'd92} : s = 106;
	{8'd245,8'd93} : s = 105;
	{8'd245,8'd94} : s = 234;
	{8'd245,8'd95} : s = 102;
	{8'd245,8'd96} : s = 233;
	{8'd245,8'd97} : s = 230;
	{8'd245,8'd98} : s = 380;
	{8'd245,8'd99} : s = 101;
	{8'd245,8'd100} : s = 229;
	{8'd245,8'd101} : s = 227;
	{8'd245,8'd102} : s = 378;
	{8'd245,8'd103} : s = 220;
	{8'd245,8'd104} : s = 377;
	{8'd245,8'd105} : s = 374;
	{8'd245,8'd106} : s = 487;
	{8'd245,8'd107} : s = 25;
	{8'd245,8'd108} : s = 99;
	{8'd245,8'd109} : s = 92;
	{8'd245,8'd110} : s = 218;
	{8'd245,8'd111} : s = 90;
	{8'd245,8'd112} : s = 217;
	{8'd245,8'd113} : s = 214;
	{8'd245,8'd114} : s = 373;
	{8'd245,8'd115} : s = 89;
	{8'd245,8'd116} : s = 213;
	{8'd245,8'd117} : s = 211;
	{8'd245,8'd118} : s = 371;
	{8'd245,8'd119} : s = 206;
	{8'd245,8'd120} : s = 366;
	{8'd245,8'd121} : s = 365;
	{8'd245,8'd122} : s = 478;
	{8'd245,8'd123} : s = 86;
	{8'd245,8'd124} : s = 205;
	{8'd245,8'd125} : s = 203;
	{8'd245,8'd126} : s = 363;
	{8'd245,8'd127} : s = 199;
	{8'd245,8'd128} : s = 359;
	{8'd245,8'd129} : s = 350;
	{8'd245,8'd130} : s = 477;
	{8'd245,8'd131} : s = 188;
	{8'd245,8'd132} : s = 349;
	{8'd245,8'd133} : s = 347;
	{8'd245,8'd134} : s = 475;
	{8'd245,8'd135} : s = 343;
	{8'd245,8'd136} : s = 471;
	{8'd245,8'd137} : s = 463;
	{8'd245,8'd138} : s = 509;
	{8'd245,8'd139} : s = 3;
	{8'd245,8'd140} : s = 22;
	{8'd245,8'd141} : s = 21;
	{8'd245,8'd142} : s = 85;
	{8'd245,8'd143} : s = 19;
	{8'd245,8'd144} : s = 83;
	{8'd245,8'd145} : s = 78;
	{8'd245,8'd146} : s = 186;
	{8'd245,8'd147} : s = 14;
	{8'd245,8'd148} : s = 77;
	{8'd245,8'd149} : s = 75;
	{8'd245,8'd150} : s = 185;
	{8'd245,8'd151} : s = 71;
	{8'd245,8'd152} : s = 182;
	{8'd245,8'd153} : s = 181;
	{8'd245,8'd154} : s = 335;
	{8'd245,8'd155} : s = 13;
	{8'd245,8'd156} : s = 60;
	{8'd245,8'd157} : s = 58;
	{8'd245,8'd158} : s = 179;
	{8'd245,8'd159} : s = 57;
	{8'd245,8'd160} : s = 174;
	{8'd245,8'd161} : s = 173;
	{8'd245,8'd162} : s = 318;
	{8'd245,8'd163} : s = 54;
	{8'd245,8'd164} : s = 171;
	{8'd245,8'd165} : s = 167;
	{8'd245,8'd166} : s = 317;
	{8'd245,8'd167} : s = 158;
	{8'd245,8'd168} : s = 315;
	{8'd245,8'd169} : s = 311;
	{8'd245,8'd170} : s = 446;
	{8'd245,8'd171} : s = 11;
	{8'd245,8'd172} : s = 53;
	{8'd245,8'd173} : s = 51;
	{8'd245,8'd174} : s = 157;
	{8'd245,8'd175} : s = 46;
	{8'd245,8'd176} : s = 155;
	{8'd245,8'd177} : s = 151;
	{8'd245,8'd178} : s = 303;
	{8'd245,8'd179} : s = 45;
	{8'd245,8'd180} : s = 143;
	{8'd245,8'd181} : s = 124;
	{8'd245,8'd182} : s = 287;
	{8'd245,8'd183} : s = 122;
	{8'd245,8'd184} : s = 252;
	{8'd245,8'd185} : s = 250;
	{8'd245,8'd186} : s = 445;
	{8'd245,8'd187} : s = 43;
	{8'd245,8'd188} : s = 121;
	{8'd245,8'd189} : s = 118;
	{8'd245,8'd190} : s = 249;
	{8'd245,8'd191} : s = 117;
	{8'd245,8'd192} : s = 246;
	{8'd245,8'd193} : s = 245;
	{8'd245,8'd194} : s = 443;
	{8'd245,8'd195} : s = 115;
	{8'd245,8'd196} : s = 243;
	{8'd245,8'd197} : s = 238;
	{8'd245,8'd198} : s = 439;
	{8'd245,8'd199} : s = 237;
	{8'd245,8'd200} : s = 431;
	{8'd245,8'd201} : s = 415;
	{8'd245,8'd202} : s = 507;
	{8'd245,8'd203} : s = 7;
	{8'd245,8'd204} : s = 39;
	{8'd245,8'd205} : s = 30;
	{8'd245,8'd206} : s = 110;
	{8'd245,8'd207} : s = 29;
	{8'd245,8'd208} : s = 109;
	{8'd245,8'd209} : s = 107;
	{8'd245,8'd210} : s = 235;
	{8'd245,8'd211} : s = 27;
	{8'd245,8'd212} : s = 103;
	{8'd245,8'd213} : s = 94;
	{8'd245,8'd214} : s = 231;
	{8'd245,8'd215} : s = 93;
	{8'd245,8'd216} : s = 222;
	{8'd245,8'd217} : s = 221;
	{8'd245,8'd218} : s = 382;
	{8'd245,8'd219} : s = 23;
	{8'd245,8'd220} : s = 91;
	{8'd245,8'd221} : s = 87;
	{8'd245,8'd222} : s = 219;
	{8'd245,8'd223} : s = 79;
	{8'd245,8'd224} : s = 215;
	{8'd245,8'd225} : s = 207;
	{8'd245,8'd226} : s = 381;
	{8'd245,8'd227} : s = 62;
	{8'd245,8'd228} : s = 190;
	{8'd245,8'd229} : s = 189;
	{8'd245,8'd230} : s = 379;
	{8'd245,8'd231} : s = 187;
	{8'd245,8'd232} : s = 375;
	{8'd245,8'd233} : s = 367;
	{8'd245,8'd234} : s = 503;
	{8'd245,8'd235} : s = 15;
	{8'd245,8'd236} : s = 61;
	{8'd245,8'd237} : s = 59;
	{8'd245,8'd238} : s = 183;
	{8'd245,8'd239} : s = 55;
	{8'd245,8'd240} : s = 175;
	{8'd245,8'd241} : s = 159;
	{8'd245,8'd242} : s = 351;
	{8'd245,8'd243} : s = 47;
	{8'd245,8'd244} : s = 126;
	{8'd245,8'd245} : s = 125;
	{8'd245,8'd246} : s = 319;
	{8'd245,8'd247} : s = 123;
	{8'd245,8'd248} : s = 254;
	{8'd245,8'd249} : s = 253;
	{8'd245,8'd250} : s = 479;
	{8'd245,8'd251} : s = 31;
	{8'd245,8'd252} : s = 119;
	{8'd245,8'd253} : s = 111;
	{8'd245,8'd254} : s = 251;
	{8'd245,8'd255} : s = 95;
	{8'd246,8'd0} : s = 437;
	{8'd246,8'd1} : s = 501;
	{8'd246,8'd2} : s = 316;
	{8'd246,8'd3} : s = 435;
	{8'd246,8'd4} : s = 430;
	{8'd246,8'd5} : s = 499;
	{8'd246,8'd6} : s = 429;
	{8'd246,8'd7} : s = 494;
	{8'd246,8'd8} : s = 493;
	{8'd246,8'd9} : s = 510;
	{8'd246,8'd10} : s = 1;
	{8'd246,8'd11} : s = 18;
	{8'd246,8'd12} : s = 17;
	{8'd246,8'd13} : s = 82;
	{8'd246,8'd14} : s = 12;
	{8'd246,8'd15} : s = 81;
	{8'd246,8'd16} : s = 76;
	{8'd246,8'd17} : s = 195;
	{8'd246,8'd18} : s = 10;
	{8'd246,8'd19} : s = 74;
	{8'd246,8'd20} : s = 73;
	{8'd246,8'd21} : s = 184;
	{8'd246,8'd22} : s = 70;
	{8'd246,8'd23} : s = 180;
	{8'd246,8'd24} : s = 178;
	{8'd246,8'd25} : s = 314;
	{8'd246,8'd26} : s = 9;
	{8'd246,8'd27} : s = 69;
	{8'd246,8'd28} : s = 67;
	{8'd246,8'd29} : s = 177;
	{8'd246,8'd30} : s = 56;
	{8'd246,8'd31} : s = 172;
	{8'd246,8'd32} : s = 170;
	{8'd246,8'd33} : s = 313;
	{8'd246,8'd34} : s = 52;
	{8'd246,8'd35} : s = 169;
	{8'd246,8'd36} : s = 166;
	{8'd246,8'd37} : s = 310;
	{8'd246,8'd38} : s = 165;
	{8'd246,8'd39} : s = 309;
	{8'd246,8'd40} : s = 307;
	{8'd246,8'd41} : s = 427;
	{8'd246,8'd42} : s = 6;
	{8'd246,8'd43} : s = 50;
	{8'd246,8'd44} : s = 49;
	{8'd246,8'd45} : s = 163;
	{8'd246,8'd46} : s = 44;
	{8'd246,8'd47} : s = 156;
	{8'd246,8'd48} : s = 154;
	{8'd246,8'd49} : s = 302;
	{8'd246,8'd50} : s = 42;
	{8'd246,8'd51} : s = 153;
	{8'd246,8'd52} : s = 150;
	{8'd246,8'd53} : s = 301;
	{8'd246,8'd54} : s = 149;
	{8'd246,8'd55} : s = 299;
	{8'd246,8'd56} : s = 295;
	{8'd246,8'd57} : s = 423;
	{8'd246,8'd58} : s = 41;
	{8'd246,8'd59} : s = 147;
	{8'd246,8'd60} : s = 142;
	{8'd246,8'd61} : s = 286;
	{8'd246,8'd62} : s = 141;
	{8'd246,8'd63} : s = 285;
	{8'd246,8'd64} : s = 283;
	{8'd246,8'd65} : s = 414;
	{8'd246,8'd66} : s = 139;
	{8'd246,8'd67} : s = 279;
	{8'd246,8'd68} : s = 271;
	{8'd246,8'd69} : s = 413;
	{8'd246,8'd70} : s = 248;
	{8'd246,8'd71} : s = 411;
	{8'd246,8'd72} : s = 407;
	{8'd246,8'd73} : s = 491;
	{8'd246,8'd74} : s = 5;
	{8'd246,8'd75} : s = 38;
	{8'd246,8'd76} : s = 37;
	{8'd246,8'd77} : s = 135;
	{8'd246,8'd78} : s = 35;
	{8'd246,8'd79} : s = 120;
	{8'd246,8'd80} : s = 116;
	{8'd246,8'd81} : s = 244;
	{8'd246,8'd82} : s = 28;
	{8'd246,8'd83} : s = 114;
	{8'd246,8'd84} : s = 113;
	{8'd246,8'd85} : s = 242;
	{8'd246,8'd86} : s = 108;
	{8'd246,8'd87} : s = 241;
	{8'd246,8'd88} : s = 236;
	{8'd246,8'd89} : s = 399;
	{8'd246,8'd90} : s = 26;
	{8'd246,8'd91} : s = 106;
	{8'd246,8'd92} : s = 105;
	{8'd246,8'd93} : s = 234;
	{8'd246,8'd94} : s = 102;
	{8'd246,8'd95} : s = 233;
	{8'd246,8'd96} : s = 230;
	{8'd246,8'd97} : s = 380;
	{8'd246,8'd98} : s = 101;
	{8'd246,8'd99} : s = 229;
	{8'd246,8'd100} : s = 227;
	{8'd246,8'd101} : s = 378;
	{8'd246,8'd102} : s = 220;
	{8'd246,8'd103} : s = 377;
	{8'd246,8'd104} : s = 374;
	{8'd246,8'd105} : s = 487;
	{8'd246,8'd106} : s = 25;
	{8'd246,8'd107} : s = 99;
	{8'd246,8'd108} : s = 92;
	{8'd246,8'd109} : s = 218;
	{8'd246,8'd110} : s = 90;
	{8'd246,8'd111} : s = 217;
	{8'd246,8'd112} : s = 214;
	{8'd246,8'd113} : s = 373;
	{8'd246,8'd114} : s = 89;
	{8'd246,8'd115} : s = 213;
	{8'd246,8'd116} : s = 211;
	{8'd246,8'd117} : s = 371;
	{8'd246,8'd118} : s = 206;
	{8'd246,8'd119} : s = 366;
	{8'd246,8'd120} : s = 365;
	{8'd246,8'd121} : s = 478;
	{8'd246,8'd122} : s = 86;
	{8'd246,8'd123} : s = 205;
	{8'd246,8'd124} : s = 203;
	{8'd246,8'd125} : s = 363;
	{8'd246,8'd126} : s = 199;
	{8'd246,8'd127} : s = 359;
	{8'd246,8'd128} : s = 350;
	{8'd246,8'd129} : s = 477;
	{8'd246,8'd130} : s = 188;
	{8'd246,8'd131} : s = 349;
	{8'd246,8'd132} : s = 347;
	{8'd246,8'd133} : s = 475;
	{8'd246,8'd134} : s = 343;
	{8'd246,8'd135} : s = 471;
	{8'd246,8'd136} : s = 463;
	{8'd246,8'd137} : s = 509;
	{8'd246,8'd138} : s = 3;
	{8'd246,8'd139} : s = 22;
	{8'd246,8'd140} : s = 21;
	{8'd246,8'd141} : s = 85;
	{8'd246,8'd142} : s = 19;
	{8'd246,8'd143} : s = 83;
	{8'd246,8'd144} : s = 78;
	{8'd246,8'd145} : s = 186;
	{8'd246,8'd146} : s = 14;
	{8'd246,8'd147} : s = 77;
	{8'd246,8'd148} : s = 75;
	{8'd246,8'd149} : s = 185;
	{8'd246,8'd150} : s = 71;
	{8'd246,8'd151} : s = 182;
	{8'd246,8'd152} : s = 181;
	{8'd246,8'd153} : s = 335;
	{8'd246,8'd154} : s = 13;
	{8'd246,8'd155} : s = 60;
	{8'd246,8'd156} : s = 58;
	{8'd246,8'd157} : s = 179;
	{8'd246,8'd158} : s = 57;
	{8'd246,8'd159} : s = 174;
	{8'd246,8'd160} : s = 173;
	{8'd246,8'd161} : s = 318;
	{8'd246,8'd162} : s = 54;
	{8'd246,8'd163} : s = 171;
	{8'd246,8'd164} : s = 167;
	{8'd246,8'd165} : s = 317;
	{8'd246,8'd166} : s = 158;
	{8'd246,8'd167} : s = 315;
	{8'd246,8'd168} : s = 311;
	{8'd246,8'd169} : s = 446;
	{8'd246,8'd170} : s = 11;
	{8'd246,8'd171} : s = 53;
	{8'd246,8'd172} : s = 51;
	{8'd246,8'd173} : s = 157;
	{8'd246,8'd174} : s = 46;
	{8'd246,8'd175} : s = 155;
	{8'd246,8'd176} : s = 151;
	{8'd246,8'd177} : s = 303;
	{8'd246,8'd178} : s = 45;
	{8'd246,8'd179} : s = 143;
	{8'd246,8'd180} : s = 124;
	{8'd246,8'd181} : s = 287;
	{8'd246,8'd182} : s = 122;
	{8'd246,8'd183} : s = 252;
	{8'd246,8'd184} : s = 250;
	{8'd246,8'd185} : s = 445;
	{8'd246,8'd186} : s = 43;
	{8'd246,8'd187} : s = 121;
	{8'd246,8'd188} : s = 118;
	{8'd246,8'd189} : s = 249;
	{8'd246,8'd190} : s = 117;
	{8'd246,8'd191} : s = 246;
	{8'd246,8'd192} : s = 245;
	{8'd246,8'd193} : s = 443;
	{8'd246,8'd194} : s = 115;
	{8'd246,8'd195} : s = 243;
	{8'd246,8'd196} : s = 238;
	{8'd246,8'd197} : s = 439;
	{8'd246,8'd198} : s = 237;
	{8'd246,8'd199} : s = 431;
	{8'd246,8'd200} : s = 415;
	{8'd246,8'd201} : s = 507;
	{8'd246,8'd202} : s = 7;
	{8'd246,8'd203} : s = 39;
	{8'd246,8'd204} : s = 30;
	{8'd246,8'd205} : s = 110;
	{8'd246,8'd206} : s = 29;
	{8'd246,8'd207} : s = 109;
	{8'd246,8'd208} : s = 107;
	{8'd246,8'd209} : s = 235;
	{8'd246,8'd210} : s = 27;
	{8'd246,8'd211} : s = 103;
	{8'd246,8'd212} : s = 94;
	{8'd246,8'd213} : s = 231;
	{8'd246,8'd214} : s = 93;
	{8'd246,8'd215} : s = 222;
	{8'd246,8'd216} : s = 221;
	{8'd246,8'd217} : s = 382;
	{8'd246,8'd218} : s = 23;
	{8'd246,8'd219} : s = 91;
	{8'd246,8'd220} : s = 87;
	{8'd246,8'd221} : s = 219;
	{8'd246,8'd222} : s = 79;
	{8'd246,8'd223} : s = 215;
	{8'd246,8'd224} : s = 207;
	{8'd246,8'd225} : s = 381;
	{8'd246,8'd226} : s = 62;
	{8'd246,8'd227} : s = 190;
	{8'd246,8'd228} : s = 189;
	{8'd246,8'd229} : s = 379;
	{8'd246,8'd230} : s = 187;
	{8'd246,8'd231} : s = 375;
	{8'd246,8'd232} : s = 367;
	{8'd246,8'd233} : s = 503;
	{8'd246,8'd234} : s = 15;
	{8'd246,8'd235} : s = 61;
	{8'd246,8'd236} : s = 59;
	{8'd246,8'd237} : s = 183;
	{8'd246,8'd238} : s = 55;
	{8'd246,8'd239} : s = 175;
	{8'd246,8'd240} : s = 159;
	{8'd246,8'd241} : s = 351;
	{8'd246,8'd242} : s = 47;
	{8'd246,8'd243} : s = 126;
	{8'd246,8'd244} : s = 125;
	{8'd246,8'd245} : s = 319;
	{8'd246,8'd246} : s = 123;
	{8'd246,8'd247} : s = 254;
	{8'd246,8'd248} : s = 253;
	{8'd246,8'd249} : s = 479;
	{8'd246,8'd250} : s = 31;
	{8'd246,8'd251} : s = 119;
	{8'd246,8'd252} : s = 111;
	{8'd246,8'd253} : s = 251;
	{8'd246,8'd254} : s = 95;
	{8'd246,8'd255} : s = 247;
	{8'd247,8'd0} : s = 501;
	{8'd247,8'd1} : s = 316;
	{8'd247,8'd2} : s = 435;
	{8'd247,8'd3} : s = 430;
	{8'd247,8'd4} : s = 499;
	{8'd247,8'd5} : s = 429;
	{8'd247,8'd6} : s = 494;
	{8'd247,8'd7} : s = 493;
	{8'd247,8'd8} : s = 510;
	{8'd247,8'd9} : s = 1;
	{8'd247,8'd10} : s = 18;
	{8'd247,8'd11} : s = 17;
	{8'd247,8'd12} : s = 82;
	{8'd247,8'd13} : s = 12;
	{8'd247,8'd14} : s = 81;
	{8'd247,8'd15} : s = 76;
	{8'd247,8'd16} : s = 195;
	{8'd247,8'd17} : s = 10;
	{8'd247,8'd18} : s = 74;
	{8'd247,8'd19} : s = 73;
	{8'd247,8'd20} : s = 184;
	{8'd247,8'd21} : s = 70;
	{8'd247,8'd22} : s = 180;
	{8'd247,8'd23} : s = 178;
	{8'd247,8'd24} : s = 314;
	{8'd247,8'd25} : s = 9;
	{8'd247,8'd26} : s = 69;
	{8'd247,8'd27} : s = 67;
	{8'd247,8'd28} : s = 177;
	{8'd247,8'd29} : s = 56;
	{8'd247,8'd30} : s = 172;
	{8'd247,8'd31} : s = 170;
	{8'd247,8'd32} : s = 313;
	{8'd247,8'd33} : s = 52;
	{8'd247,8'd34} : s = 169;
	{8'd247,8'd35} : s = 166;
	{8'd247,8'd36} : s = 310;
	{8'd247,8'd37} : s = 165;
	{8'd247,8'd38} : s = 309;
	{8'd247,8'd39} : s = 307;
	{8'd247,8'd40} : s = 427;
	{8'd247,8'd41} : s = 6;
	{8'd247,8'd42} : s = 50;
	{8'd247,8'd43} : s = 49;
	{8'd247,8'd44} : s = 163;
	{8'd247,8'd45} : s = 44;
	{8'd247,8'd46} : s = 156;
	{8'd247,8'd47} : s = 154;
	{8'd247,8'd48} : s = 302;
	{8'd247,8'd49} : s = 42;
	{8'd247,8'd50} : s = 153;
	{8'd247,8'd51} : s = 150;
	{8'd247,8'd52} : s = 301;
	{8'd247,8'd53} : s = 149;
	{8'd247,8'd54} : s = 299;
	{8'd247,8'd55} : s = 295;
	{8'd247,8'd56} : s = 423;
	{8'd247,8'd57} : s = 41;
	{8'd247,8'd58} : s = 147;
	{8'd247,8'd59} : s = 142;
	{8'd247,8'd60} : s = 286;
	{8'd247,8'd61} : s = 141;
	{8'd247,8'd62} : s = 285;
	{8'd247,8'd63} : s = 283;
	{8'd247,8'd64} : s = 414;
	{8'd247,8'd65} : s = 139;
	{8'd247,8'd66} : s = 279;
	{8'd247,8'd67} : s = 271;
	{8'd247,8'd68} : s = 413;
	{8'd247,8'd69} : s = 248;
	{8'd247,8'd70} : s = 411;
	{8'd247,8'd71} : s = 407;
	{8'd247,8'd72} : s = 491;
	{8'd247,8'd73} : s = 5;
	{8'd247,8'd74} : s = 38;
	{8'd247,8'd75} : s = 37;
	{8'd247,8'd76} : s = 135;
	{8'd247,8'd77} : s = 35;
	{8'd247,8'd78} : s = 120;
	{8'd247,8'd79} : s = 116;
	{8'd247,8'd80} : s = 244;
	{8'd247,8'd81} : s = 28;
	{8'd247,8'd82} : s = 114;
	{8'd247,8'd83} : s = 113;
	{8'd247,8'd84} : s = 242;
	{8'd247,8'd85} : s = 108;
	{8'd247,8'd86} : s = 241;
	{8'd247,8'd87} : s = 236;
	{8'd247,8'd88} : s = 399;
	{8'd247,8'd89} : s = 26;
	{8'd247,8'd90} : s = 106;
	{8'd247,8'd91} : s = 105;
	{8'd247,8'd92} : s = 234;
	{8'd247,8'd93} : s = 102;
	{8'd247,8'd94} : s = 233;
	{8'd247,8'd95} : s = 230;
	{8'd247,8'd96} : s = 380;
	{8'd247,8'd97} : s = 101;
	{8'd247,8'd98} : s = 229;
	{8'd247,8'd99} : s = 227;
	{8'd247,8'd100} : s = 378;
	{8'd247,8'd101} : s = 220;
	{8'd247,8'd102} : s = 377;
	{8'd247,8'd103} : s = 374;
	{8'd247,8'd104} : s = 487;
	{8'd247,8'd105} : s = 25;
	{8'd247,8'd106} : s = 99;
	{8'd247,8'd107} : s = 92;
	{8'd247,8'd108} : s = 218;
	{8'd247,8'd109} : s = 90;
	{8'd247,8'd110} : s = 217;
	{8'd247,8'd111} : s = 214;
	{8'd247,8'd112} : s = 373;
	{8'd247,8'd113} : s = 89;
	{8'd247,8'd114} : s = 213;
	{8'd247,8'd115} : s = 211;
	{8'd247,8'd116} : s = 371;
	{8'd247,8'd117} : s = 206;
	{8'd247,8'd118} : s = 366;
	{8'd247,8'd119} : s = 365;
	{8'd247,8'd120} : s = 478;
	{8'd247,8'd121} : s = 86;
	{8'd247,8'd122} : s = 205;
	{8'd247,8'd123} : s = 203;
	{8'd247,8'd124} : s = 363;
	{8'd247,8'd125} : s = 199;
	{8'd247,8'd126} : s = 359;
	{8'd247,8'd127} : s = 350;
	{8'd247,8'd128} : s = 477;
	{8'd247,8'd129} : s = 188;
	{8'd247,8'd130} : s = 349;
	{8'd247,8'd131} : s = 347;
	{8'd247,8'd132} : s = 475;
	{8'd247,8'd133} : s = 343;
	{8'd247,8'd134} : s = 471;
	{8'd247,8'd135} : s = 463;
	{8'd247,8'd136} : s = 509;
	{8'd247,8'd137} : s = 3;
	{8'd247,8'd138} : s = 22;
	{8'd247,8'd139} : s = 21;
	{8'd247,8'd140} : s = 85;
	{8'd247,8'd141} : s = 19;
	{8'd247,8'd142} : s = 83;
	{8'd247,8'd143} : s = 78;
	{8'd247,8'd144} : s = 186;
	{8'd247,8'd145} : s = 14;
	{8'd247,8'd146} : s = 77;
	{8'd247,8'd147} : s = 75;
	{8'd247,8'd148} : s = 185;
	{8'd247,8'd149} : s = 71;
	{8'd247,8'd150} : s = 182;
	{8'd247,8'd151} : s = 181;
	{8'd247,8'd152} : s = 335;
	{8'd247,8'd153} : s = 13;
	{8'd247,8'd154} : s = 60;
	{8'd247,8'd155} : s = 58;
	{8'd247,8'd156} : s = 179;
	{8'd247,8'd157} : s = 57;
	{8'd247,8'd158} : s = 174;
	{8'd247,8'd159} : s = 173;
	{8'd247,8'd160} : s = 318;
	{8'd247,8'd161} : s = 54;
	{8'd247,8'd162} : s = 171;
	{8'd247,8'd163} : s = 167;
	{8'd247,8'd164} : s = 317;
	{8'd247,8'd165} : s = 158;
	{8'd247,8'd166} : s = 315;
	{8'd247,8'd167} : s = 311;
	{8'd247,8'd168} : s = 446;
	{8'd247,8'd169} : s = 11;
	{8'd247,8'd170} : s = 53;
	{8'd247,8'd171} : s = 51;
	{8'd247,8'd172} : s = 157;
	{8'd247,8'd173} : s = 46;
	{8'd247,8'd174} : s = 155;
	{8'd247,8'd175} : s = 151;
	{8'd247,8'd176} : s = 303;
	{8'd247,8'd177} : s = 45;
	{8'd247,8'd178} : s = 143;
	{8'd247,8'd179} : s = 124;
	{8'd247,8'd180} : s = 287;
	{8'd247,8'd181} : s = 122;
	{8'd247,8'd182} : s = 252;
	{8'd247,8'd183} : s = 250;
	{8'd247,8'd184} : s = 445;
	{8'd247,8'd185} : s = 43;
	{8'd247,8'd186} : s = 121;
	{8'd247,8'd187} : s = 118;
	{8'd247,8'd188} : s = 249;
	{8'd247,8'd189} : s = 117;
	{8'd247,8'd190} : s = 246;
	{8'd247,8'd191} : s = 245;
	{8'd247,8'd192} : s = 443;
	{8'd247,8'd193} : s = 115;
	{8'd247,8'd194} : s = 243;
	{8'd247,8'd195} : s = 238;
	{8'd247,8'd196} : s = 439;
	{8'd247,8'd197} : s = 237;
	{8'd247,8'd198} : s = 431;
	{8'd247,8'd199} : s = 415;
	{8'd247,8'd200} : s = 507;
	{8'd247,8'd201} : s = 7;
	{8'd247,8'd202} : s = 39;
	{8'd247,8'd203} : s = 30;
	{8'd247,8'd204} : s = 110;
	{8'd247,8'd205} : s = 29;
	{8'd247,8'd206} : s = 109;
	{8'd247,8'd207} : s = 107;
	{8'd247,8'd208} : s = 235;
	{8'd247,8'd209} : s = 27;
	{8'd247,8'd210} : s = 103;
	{8'd247,8'd211} : s = 94;
	{8'd247,8'd212} : s = 231;
	{8'd247,8'd213} : s = 93;
	{8'd247,8'd214} : s = 222;
	{8'd247,8'd215} : s = 221;
	{8'd247,8'd216} : s = 382;
	{8'd247,8'd217} : s = 23;
	{8'd247,8'd218} : s = 91;
	{8'd247,8'd219} : s = 87;
	{8'd247,8'd220} : s = 219;
	{8'd247,8'd221} : s = 79;
	{8'd247,8'd222} : s = 215;
	{8'd247,8'd223} : s = 207;
	{8'd247,8'd224} : s = 381;
	{8'd247,8'd225} : s = 62;
	{8'd247,8'd226} : s = 190;
	{8'd247,8'd227} : s = 189;
	{8'd247,8'd228} : s = 379;
	{8'd247,8'd229} : s = 187;
	{8'd247,8'd230} : s = 375;
	{8'd247,8'd231} : s = 367;
	{8'd247,8'd232} : s = 503;
	{8'd247,8'd233} : s = 15;
	{8'd247,8'd234} : s = 61;
	{8'd247,8'd235} : s = 59;
	{8'd247,8'd236} : s = 183;
	{8'd247,8'd237} : s = 55;
	{8'd247,8'd238} : s = 175;
	{8'd247,8'd239} : s = 159;
	{8'd247,8'd240} : s = 351;
	{8'd247,8'd241} : s = 47;
	{8'd247,8'd242} : s = 126;
	{8'd247,8'd243} : s = 125;
	{8'd247,8'd244} : s = 319;
	{8'd247,8'd245} : s = 123;
	{8'd247,8'd246} : s = 254;
	{8'd247,8'd247} : s = 253;
	{8'd247,8'd248} : s = 479;
	{8'd247,8'd249} : s = 31;
	{8'd247,8'd250} : s = 119;
	{8'd247,8'd251} : s = 111;
	{8'd247,8'd252} : s = 251;
	{8'd247,8'd253} : s = 95;
	{8'd247,8'd254} : s = 247;
	{8'd247,8'd255} : s = 239;
	{8'd248,8'd0} : s = 316;
	{8'd248,8'd1} : s = 435;
	{8'd248,8'd2} : s = 430;
	{8'd248,8'd3} : s = 499;
	{8'd248,8'd4} : s = 429;
	{8'd248,8'd5} : s = 494;
	{8'd248,8'd6} : s = 493;
	{8'd248,8'd7} : s = 510;
	{8'd248,8'd8} : s = 1;
	{8'd248,8'd9} : s = 18;
	{8'd248,8'd10} : s = 17;
	{8'd248,8'd11} : s = 82;
	{8'd248,8'd12} : s = 12;
	{8'd248,8'd13} : s = 81;
	{8'd248,8'd14} : s = 76;
	{8'd248,8'd15} : s = 195;
	{8'd248,8'd16} : s = 10;
	{8'd248,8'd17} : s = 74;
	{8'd248,8'd18} : s = 73;
	{8'd248,8'd19} : s = 184;
	{8'd248,8'd20} : s = 70;
	{8'd248,8'd21} : s = 180;
	{8'd248,8'd22} : s = 178;
	{8'd248,8'd23} : s = 314;
	{8'd248,8'd24} : s = 9;
	{8'd248,8'd25} : s = 69;
	{8'd248,8'd26} : s = 67;
	{8'd248,8'd27} : s = 177;
	{8'd248,8'd28} : s = 56;
	{8'd248,8'd29} : s = 172;
	{8'd248,8'd30} : s = 170;
	{8'd248,8'd31} : s = 313;
	{8'd248,8'd32} : s = 52;
	{8'd248,8'd33} : s = 169;
	{8'd248,8'd34} : s = 166;
	{8'd248,8'd35} : s = 310;
	{8'd248,8'd36} : s = 165;
	{8'd248,8'd37} : s = 309;
	{8'd248,8'd38} : s = 307;
	{8'd248,8'd39} : s = 427;
	{8'd248,8'd40} : s = 6;
	{8'd248,8'd41} : s = 50;
	{8'd248,8'd42} : s = 49;
	{8'd248,8'd43} : s = 163;
	{8'd248,8'd44} : s = 44;
	{8'd248,8'd45} : s = 156;
	{8'd248,8'd46} : s = 154;
	{8'd248,8'd47} : s = 302;
	{8'd248,8'd48} : s = 42;
	{8'd248,8'd49} : s = 153;
	{8'd248,8'd50} : s = 150;
	{8'd248,8'd51} : s = 301;
	{8'd248,8'd52} : s = 149;
	{8'd248,8'd53} : s = 299;
	{8'd248,8'd54} : s = 295;
	{8'd248,8'd55} : s = 423;
	{8'd248,8'd56} : s = 41;
	{8'd248,8'd57} : s = 147;
	{8'd248,8'd58} : s = 142;
	{8'd248,8'd59} : s = 286;
	{8'd248,8'd60} : s = 141;
	{8'd248,8'd61} : s = 285;
	{8'd248,8'd62} : s = 283;
	{8'd248,8'd63} : s = 414;
	{8'd248,8'd64} : s = 139;
	{8'd248,8'd65} : s = 279;
	{8'd248,8'd66} : s = 271;
	{8'd248,8'd67} : s = 413;
	{8'd248,8'd68} : s = 248;
	{8'd248,8'd69} : s = 411;
	{8'd248,8'd70} : s = 407;
	{8'd248,8'd71} : s = 491;
	{8'd248,8'd72} : s = 5;
	{8'd248,8'd73} : s = 38;
	{8'd248,8'd74} : s = 37;
	{8'd248,8'd75} : s = 135;
	{8'd248,8'd76} : s = 35;
	{8'd248,8'd77} : s = 120;
	{8'd248,8'd78} : s = 116;
	{8'd248,8'd79} : s = 244;
	{8'd248,8'd80} : s = 28;
	{8'd248,8'd81} : s = 114;
	{8'd248,8'd82} : s = 113;
	{8'd248,8'd83} : s = 242;
	{8'd248,8'd84} : s = 108;
	{8'd248,8'd85} : s = 241;
	{8'd248,8'd86} : s = 236;
	{8'd248,8'd87} : s = 399;
	{8'd248,8'd88} : s = 26;
	{8'd248,8'd89} : s = 106;
	{8'd248,8'd90} : s = 105;
	{8'd248,8'd91} : s = 234;
	{8'd248,8'd92} : s = 102;
	{8'd248,8'd93} : s = 233;
	{8'd248,8'd94} : s = 230;
	{8'd248,8'd95} : s = 380;
	{8'd248,8'd96} : s = 101;
	{8'd248,8'd97} : s = 229;
	{8'd248,8'd98} : s = 227;
	{8'd248,8'd99} : s = 378;
	{8'd248,8'd100} : s = 220;
	{8'd248,8'd101} : s = 377;
	{8'd248,8'd102} : s = 374;
	{8'd248,8'd103} : s = 487;
	{8'd248,8'd104} : s = 25;
	{8'd248,8'd105} : s = 99;
	{8'd248,8'd106} : s = 92;
	{8'd248,8'd107} : s = 218;
	{8'd248,8'd108} : s = 90;
	{8'd248,8'd109} : s = 217;
	{8'd248,8'd110} : s = 214;
	{8'd248,8'd111} : s = 373;
	{8'd248,8'd112} : s = 89;
	{8'd248,8'd113} : s = 213;
	{8'd248,8'd114} : s = 211;
	{8'd248,8'd115} : s = 371;
	{8'd248,8'd116} : s = 206;
	{8'd248,8'd117} : s = 366;
	{8'd248,8'd118} : s = 365;
	{8'd248,8'd119} : s = 478;
	{8'd248,8'd120} : s = 86;
	{8'd248,8'd121} : s = 205;
	{8'd248,8'd122} : s = 203;
	{8'd248,8'd123} : s = 363;
	{8'd248,8'd124} : s = 199;
	{8'd248,8'd125} : s = 359;
	{8'd248,8'd126} : s = 350;
	{8'd248,8'd127} : s = 477;
	{8'd248,8'd128} : s = 188;
	{8'd248,8'd129} : s = 349;
	{8'd248,8'd130} : s = 347;
	{8'd248,8'd131} : s = 475;
	{8'd248,8'd132} : s = 343;
	{8'd248,8'd133} : s = 471;
	{8'd248,8'd134} : s = 463;
	{8'd248,8'd135} : s = 509;
	{8'd248,8'd136} : s = 3;
	{8'd248,8'd137} : s = 22;
	{8'd248,8'd138} : s = 21;
	{8'd248,8'd139} : s = 85;
	{8'd248,8'd140} : s = 19;
	{8'd248,8'd141} : s = 83;
	{8'd248,8'd142} : s = 78;
	{8'd248,8'd143} : s = 186;
	{8'd248,8'd144} : s = 14;
	{8'd248,8'd145} : s = 77;
	{8'd248,8'd146} : s = 75;
	{8'd248,8'd147} : s = 185;
	{8'd248,8'd148} : s = 71;
	{8'd248,8'd149} : s = 182;
	{8'd248,8'd150} : s = 181;
	{8'd248,8'd151} : s = 335;
	{8'd248,8'd152} : s = 13;
	{8'd248,8'd153} : s = 60;
	{8'd248,8'd154} : s = 58;
	{8'd248,8'd155} : s = 179;
	{8'd248,8'd156} : s = 57;
	{8'd248,8'd157} : s = 174;
	{8'd248,8'd158} : s = 173;
	{8'd248,8'd159} : s = 318;
	{8'd248,8'd160} : s = 54;
	{8'd248,8'd161} : s = 171;
	{8'd248,8'd162} : s = 167;
	{8'd248,8'd163} : s = 317;
	{8'd248,8'd164} : s = 158;
	{8'd248,8'd165} : s = 315;
	{8'd248,8'd166} : s = 311;
	{8'd248,8'd167} : s = 446;
	{8'd248,8'd168} : s = 11;
	{8'd248,8'd169} : s = 53;
	{8'd248,8'd170} : s = 51;
	{8'd248,8'd171} : s = 157;
	{8'd248,8'd172} : s = 46;
	{8'd248,8'd173} : s = 155;
	{8'd248,8'd174} : s = 151;
	{8'd248,8'd175} : s = 303;
	{8'd248,8'd176} : s = 45;
	{8'd248,8'd177} : s = 143;
	{8'd248,8'd178} : s = 124;
	{8'd248,8'd179} : s = 287;
	{8'd248,8'd180} : s = 122;
	{8'd248,8'd181} : s = 252;
	{8'd248,8'd182} : s = 250;
	{8'd248,8'd183} : s = 445;
	{8'd248,8'd184} : s = 43;
	{8'd248,8'd185} : s = 121;
	{8'd248,8'd186} : s = 118;
	{8'd248,8'd187} : s = 249;
	{8'd248,8'd188} : s = 117;
	{8'd248,8'd189} : s = 246;
	{8'd248,8'd190} : s = 245;
	{8'd248,8'd191} : s = 443;
	{8'd248,8'd192} : s = 115;
	{8'd248,8'd193} : s = 243;
	{8'd248,8'd194} : s = 238;
	{8'd248,8'd195} : s = 439;
	{8'd248,8'd196} : s = 237;
	{8'd248,8'd197} : s = 431;
	{8'd248,8'd198} : s = 415;
	{8'd248,8'd199} : s = 507;
	{8'd248,8'd200} : s = 7;
	{8'd248,8'd201} : s = 39;
	{8'd248,8'd202} : s = 30;
	{8'd248,8'd203} : s = 110;
	{8'd248,8'd204} : s = 29;
	{8'd248,8'd205} : s = 109;
	{8'd248,8'd206} : s = 107;
	{8'd248,8'd207} : s = 235;
	{8'd248,8'd208} : s = 27;
	{8'd248,8'd209} : s = 103;
	{8'd248,8'd210} : s = 94;
	{8'd248,8'd211} : s = 231;
	{8'd248,8'd212} : s = 93;
	{8'd248,8'd213} : s = 222;
	{8'd248,8'd214} : s = 221;
	{8'd248,8'd215} : s = 382;
	{8'd248,8'd216} : s = 23;
	{8'd248,8'd217} : s = 91;
	{8'd248,8'd218} : s = 87;
	{8'd248,8'd219} : s = 219;
	{8'd248,8'd220} : s = 79;
	{8'd248,8'd221} : s = 215;
	{8'd248,8'd222} : s = 207;
	{8'd248,8'd223} : s = 381;
	{8'd248,8'd224} : s = 62;
	{8'd248,8'd225} : s = 190;
	{8'd248,8'd226} : s = 189;
	{8'd248,8'd227} : s = 379;
	{8'd248,8'd228} : s = 187;
	{8'd248,8'd229} : s = 375;
	{8'd248,8'd230} : s = 367;
	{8'd248,8'd231} : s = 503;
	{8'd248,8'd232} : s = 15;
	{8'd248,8'd233} : s = 61;
	{8'd248,8'd234} : s = 59;
	{8'd248,8'd235} : s = 183;
	{8'd248,8'd236} : s = 55;
	{8'd248,8'd237} : s = 175;
	{8'd248,8'd238} : s = 159;
	{8'd248,8'd239} : s = 351;
	{8'd248,8'd240} : s = 47;
	{8'd248,8'd241} : s = 126;
	{8'd248,8'd242} : s = 125;
	{8'd248,8'd243} : s = 319;
	{8'd248,8'd244} : s = 123;
	{8'd248,8'd245} : s = 254;
	{8'd248,8'd246} : s = 253;
	{8'd248,8'd247} : s = 479;
	{8'd248,8'd248} : s = 31;
	{8'd248,8'd249} : s = 119;
	{8'd248,8'd250} : s = 111;
	{8'd248,8'd251} : s = 251;
	{8'd248,8'd252} : s = 95;
	{8'd248,8'd253} : s = 247;
	{8'd248,8'd254} : s = 239;
	{8'd248,8'd255} : s = 495;
	{8'd249,8'd0} : s = 435;
	{8'd249,8'd1} : s = 430;
	{8'd249,8'd2} : s = 499;
	{8'd249,8'd3} : s = 429;
	{8'd249,8'd4} : s = 494;
	{8'd249,8'd5} : s = 493;
	{8'd249,8'd6} : s = 510;
	{8'd249,8'd7} : s = 1;
	{8'd249,8'd8} : s = 18;
	{8'd249,8'd9} : s = 17;
	{8'd249,8'd10} : s = 82;
	{8'd249,8'd11} : s = 12;
	{8'd249,8'd12} : s = 81;
	{8'd249,8'd13} : s = 76;
	{8'd249,8'd14} : s = 195;
	{8'd249,8'd15} : s = 10;
	{8'd249,8'd16} : s = 74;
	{8'd249,8'd17} : s = 73;
	{8'd249,8'd18} : s = 184;
	{8'd249,8'd19} : s = 70;
	{8'd249,8'd20} : s = 180;
	{8'd249,8'd21} : s = 178;
	{8'd249,8'd22} : s = 314;
	{8'd249,8'd23} : s = 9;
	{8'd249,8'd24} : s = 69;
	{8'd249,8'd25} : s = 67;
	{8'd249,8'd26} : s = 177;
	{8'd249,8'd27} : s = 56;
	{8'd249,8'd28} : s = 172;
	{8'd249,8'd29} : s = 170;
	{8'd249,8'd30} : s = 313;
	{8'd249,8'd31} : s = 52;
	{8'd249,8'd32} : s = 169;
	{8'd249,8'd33} : s = 166;
	{8'd249,8'd34} : s = 310;
	{8'd249,8'd35} : s = 165;
	{8'd249,8'd36} : s = 309;
	{8'd249,8'd37} : s = 307;
	{8'd249,8'd38} : s = 427;
	{8'd249,8'd39} : s = 6;
	{8'd249,8'd40} : s = 50;
	{8'd249,8'd41} : s = 49;
	{8'd249,8'd42} : s = 163;
	{8'd249,8'd43} : s = 44;
	{8'd249,8'd44} : s = 156;
	{8'd249,8'd45} : s = 154;
	{8'd249,8'd46} : s = 302;
	{8'd249,8'd47} : s = 42;
	{8'd249,8'd48} : s = 153;
	{8'd249,8'd49} : s = 150;
	{8'd249,8'd50} : s = 301;
	{8'd249,8'd51} : s = 149;
	{8'd249,8'd52} : s = 299;
	{8'd249,8'd53} : s = 295;
	{8'd249,8'd54} : s = 423;
	{8'd249,8'd55} : s = 41;
	{8'd249,8'd56} : s = 147;
	{8'd249,8'd57} : s = 142;
	{8'd249,8'd58} : s = 286;
	{8'd249,8'd59} : s = 141;
	{8'd249,8'd60} : s = 285;
	{8'd249,8'd61} : s = 283;
	{8'd249,8'd62} : s = 414;
	{8'd249,8'd63} : s = 139;
	{8'd249,8'd64} : s = 279;
	{8'd249,8'd65} : s = 271;
	{8'd249,8'd66} : s = 413;
	{8'd249,8'd67} : s = 248;
	{8'd249,8'd68} : s = 411;
	{8'd249,8'd69} : s = 407;
	{8'd249,8'd70} : s = 491;
	{8'd249,8'd71} : s = 5;
	{8'd249,8'd72} : s = 38;
	{8'd249,8'd73} : s = 37;
	{8'd249,8'd74} : s = 135;
	{8'd249,8'd75} : s = 35;
	{8'd249,8'd76} : s = 120;
	{8'd249,8'd77} : s = 116;
	{8'd249,8'd78} : s = 244;
	{8'd249,8'd79} : s = 28;
	{8'd249,8'd80} : s = 114;
	{8'd249,8'd81} : s = 113;
	{8'd249,8'd82} : s = 242;
	{8'd249,8'd83} : s = 108;
	{8'd249,8'd84} : s = 241;
	{8'd249,8'd85} : s = 236;
	{8'd249,8'd86} : s = 399;
	{8'd249,8'd87} : s = 26;
	{8'd249,8'd88} : s = 106;
	{8'd249,8'd89} : s = 105;
	{8'd249,8'd90} : s = 234;
	{8'd249,8'd91} : s = 102;
	{8'd249,8'd92} : s = 233;
	{8'd249,8'd93} : s = 230;
	{8'd249,8'd94} : s = 380;
	{8'd249,8'd95} : s = 101;
	{8'd249,8'd96} : s = 229;
	{8'd249,8'd97} : s = 227;
	{8'd249,8'd98} : s = 378;
	{8'd249,8'd99} : s = 220;
	{8'd249,8'd100} : s = 377;
	{8'd249,8'd101} : s = 374;
	{8'd249,8'd102} : s = 487;
	{8'd249,8'd103} : s = 25;
	{8'd249,8'd104} : s = 99;
	{8'd249,8'd105} : s = 92;
	{8'd249,8'd106} : s = 218;
	{8'd249,8'd107} : s = 90;
	{8'd249,8'd108} : s = 217;
	{8'd249,8'd109} : s = 214;
	{8'd249,8'd110} : s = 373;
	{8'd249,8'd111} : s = 89;
	{8'd249,8'd112} : s = 213;
	{8'd249,8'd113} : s = 211;
	{8'd249,8'd114} : s = 371;
	{8'd249,8'd115} : s = 206;
	{8'd249,8'd116} : s = 366;
	{8'd249,8'd117} : s = 365;
	{8'd249,8'd118} : s = 478;
	{8'd249,8'd119} : s = 86;
	{8'd249,8'd120} : s = 205;
	{8'd249,8'd121} : s = 203;
	{8'd249,8'd122} : s = 363;
	{8'd249,8'd123} : s = 199;
	{8'd249,8'd124} : s = 359;
	{8'd249,8'd125} : s = 350;
	{8'd249,8'd126} : s = 477;
	{8'd249,8'd127} : s = 188;
	{8'd249,8'd128} : s = 349;
	{8'd249,8'd129} : s = 347;
	{8'd249,8'd130} : s = 475;
	{8'd249,8'd131} : s = 343;
	{8'd249,8'd132} : s = 471;
	{8'd249,8'd133} : s = 463;
	{8'd249,8'd134} : s = 509;
	{8'd249,8'd135} : s = 3;
	{8'd249,8'd136} : s = 22;
	{8'd249,8'd137} : s = 21;
	{8'd249,8'd138} : s = 85;
	{8'd249,8'd139} : s = 19;
	{8'd249,8'd140} : s = 83;
	{8'd249,8'd141} : s = 78;
	{8'd249,8'd142} : s = 186;
	{8'd249,8'd143} : s = 14;
	{8'd249,8'd144} : s = 77;
	{8'd249,8'd145} : s = 75;
	{8'd249,8'd146} : s = 185;
	{8'd249,8'd147} : s = 71;
	{8'd249,8'd148} : s = 182;
	{8'd249,8'd149} : s = 181;
	{8'd249,8'd150} : s = 335;
	{8'd249,8'd151} : s = 13;
	{8'd249,8'd152} : s = 60;
	{8'd249,8'd153} : s = 58;
	{8'd249,8'd154} : s = 179;
	{8'd249,8'd155} : s = 57;
	{8'd249,8'd156} : s = 174;
	{8'd249,8'd157} : s = 173;
	{8'd249,8'd158} : s = 318;
	{8'd249,8'd159} : s = 54;
	{8'd249,8'd160} : s = 171;
	{8'd249,8'd161} : s = 167;
	{8'd249,8'd162} : s = 317;
	{8'd249,8'd163} : s = 158;
	{8'd249,8'd164} : s = 315;
	{8'd249,8'd165} : s = 311;
	{8'd249,8'd166} : s = 446;
	{8'd249,8'd167} : s = 11;
	{8'd249,8'd168} : s = 53;
	{8'd249,8'd169} : s = 51;
	{8'd249,8'd170} : s = 157;
	{8'd249,8'd171} : s = 46;
	{8'd249,8'd172} : s = 155;
	{8'd249,8'd173} : s = 151;
	{8'd249,8'd174} : s = 303;
	{8'd249,8'd175} : s = 45;
	{8'd249,8'd176} : s = 143;
	{8'd249,8'd177} : s = 124;
	{8'd249,8'd178} : s = 287;
	{8'd249,8'd179} : s = 122;
	{8'd249,8'd180} : s = 252;
	{8'd249,8'd181} : s = 250;
	{8'd249,8'd182} : s = 445;
	{8'd249,8'd183} : s = 43;
	{8'd249,8'd184} : s = 121;
	{8'd249,8'd185} : s = 118;
	{8'd249,8'd186} : s = 249;
	{8'd249,8'd187} : s = 117;
	{8'd249,8'd188} : s = 246;
	{8'd249,8'd189} : s = 245;
	{8'd249,8'd190} : s = 443;
	{8'd249,8'd191} : s = 115;
	{8'd249,8'd192} : s = 243;
	{8'd249,8'd193} : s = 238;
	{8'd249,8'd194} : s = 439;
	{8'd249,8'd195} : s = 237;
	{8'd249,8'd196} : s = 431;
	{8'd249,8'd197} : s = 415;
	{8'd249,8'd198} : s = 507;
	{8'd249,8'd199} : s = 7;
	{8'd249,8'd200} : s = 39;
	{8'd249,8'd201} : s = 30;
	{8'd249,8'd202} : s = 110;
	{8'd249,8'd203} : s = 29;
	{8'd249,8'd204} : s = 109;
	{8'd249,8'd205} : s = 107;
	{8'd249,8'd206} : s = 235;
	{8'd249,8'd207} : s = 27;
	{8'd249,8'd208} : s = 103;
	{8'd249,8'd209} : s = 94;
	{8'd249,8'd210} : s = 231;
	{8'd249,8'd211} : s = 93;
	{8'd249,8'd212} : s = 222;
	{8'd249,8'd213} : s = 221;
	{8'd249,8'd214} : s = 382;
	{8'd249,8'd215} : s = 23;
	{8'd249,8'd216} : s = 91;
	{8'd249,8'd217} : s = 87;
	{8'd249,8'd218} : s = 219;
	{8'd249,8'd219} : s = 79;
	{8'd249,8'd220} : s = 215;
	{8'd249,8'd221} : s = 207;
	{8'd249,8'd222} : s = 381;
	{8'd249,8'd223} : s = 62;
	{8'd249,8'd224} : s = 190;
	{8'd249,8'd225} : s = 189;
	{8'd249,8'd226} : s = 379;
	{8'd249,8'd227} : s = 187;
	{8'd249,8'd228} : s = 375;
	{8'd249,8'd229} : s = 367;
	{8'd249,8'd230} : s = 503;
	{8'd249,8'd231} : s = 15;
	{8'd249,8'd232} : s = 61;
	{8'd249,8'd233} : s = 59;
	{8'd249,8'd234} : s = 183;
	{8'd249,8'd235} : s = 55;
	{8'd249,8'd236} : s = 175;
	{8'd249,8'd237} : s = 159;
	{8'd249,8'd238} : s = 351;
	{8'd249,8'd239} : s = 47;
	{8'd249,8'd240} : s = 126;
	{8'd249,8'd241} : s = 125;
	{8'd249,8'd242} : s = 319;
	{8'd249,8'd243} : s = 123;
	{8'd249,8'd244} : s = 254;
	{8'd249,8'd245} : s = 253;
	{8'd249,8'd246} : s = 479;
	{8'd249,8'd247} : s = 31;
	{8'd249,8'd248} : s = 119;
	{8'd249,8'd249} : s = 111;
	{8'd249,8'd250} : s = 251;
	{8'd249,8'd251} : s = 95;
	{8'd249,8'd252} : s = 247;
	{8'd249,8'd253} : s = 239;
	{8'd249,8'd254} : s = 495;
	{8'd249,8'd255} : s = 63;
	{8'd250,8'd0} : s = 430;
	{8'd250,8'd1} : s = 499;
	{8'd250,8'd2} : s = 429;
	{8'd250,8'd3} : s = 494;
	{8'd250,8'd4} : s = 493;
	{8'd250,8'd5} : s = 510;
	{8'd250,8'd6} : s = 1;
	{8'd250,8'd7} : s = 18;
	{8'd250,8'd8} : s = 17;
	{8'd250,8'd9} : s = 82;
	{8'd250,8'd10} : s = 12;
	{8'd250,8'd11} : s = 81;
	{8'd250,8'd12} : s = 76;
	{8'd250,8'd13} : s = 195;
	{8'd250,8'd14} : s = 10;
	{8'd250,8'd15} : s = 74;
	{8'd250,8'd16} : s = 73;
	{8'd250,8'd17} : s = 184;
	{8'd250,8'd18} : s = 70;
	{8'd250,8'd19} : s = 180;
	{8'd250,8'd20} : s = 178;
	{8'd250,8'd21} : s = 314;
	{8'd250,8'd22} : s = 9;
	{8'd250,8'd23} : s = 69;
	{8'd250,8'd24} : s = 67;
	{8'd250,8'd25} : s = 177;
	{8'd250,8'd26} : s = 56;
	{8'd250,8'd27} : s = 172;
	{8'd250,8'd28} : s = 170;
	{8'd250,8'd29} : s = 313;
	{8'd250,8'd30} : s = 52;
	{8'd250,8'd31} : s = 169;
	{8'd250,8'd32} : s = 166;
	{8'd250,8'd33} : s = 310;
	{8'd250,8'd34} : s = 165;
	{8'd250,8'd35} : s = 309;
	{8'd250,8'd36} : s = 307;
	{8'd250,8'd37} : s = 427;
	{8'd250,8'd38} : s = 6;
	{8'd250,8'd39} : s = 50;
	{8'd250,8'd40} : s = 49;
	{8'd250,8'd41} : s = 163;
	{8'd250,8'd42} : s = 44;
	{8'd250,8'd43} : s = 156;
	{8'd250,8'd44} : s = 154;
	{8'd250,8'd45} : s = 302;
	{8'd250,8'd46} : s = 42;
	{8'd250,8'd47} : s = 153;
	{8'd250,8'd48} : s = 150;
	{8'd250,8'd49} : s = 301;
	{8'd250,8'd50} : s = 149;
	{8'd250,8'd51} : s = 299;
	{8'd250,8'd52} : s = 295;
	{8'd250,8'd53} : s = 423;
	{8'd250,8'd54} : s = 41;
	{8'd250,8'd55} : s = 147;
	{8'd250,8'd56} : s = 142;
	{8'd250,8'd57} : s = 286;
	{8'd250,8'd58} : s = 141;
	{8'd250,8'd59} : s = 285;
	{8'd250,8'd60} : s = 283;
	{8'd250,8'd61} : s = 414;
	{8'd250,8'd62} : s = 139;
	{8'd250,8'd63} : s = 279;
	{8'd250,8'd64} : s = 271;
	{8'd250,8'd65} : s = 413;
	{8'd250,8'd66} : s = 248;
	{8'd250,8'd67} : s = 411;
	{8'd250,8'd68} : s = 407;
	{8'd250,8'd69} : s = 491;
	{8'd250,8'd70} : s = 5;
	{8'd250,8'd71} : s = 38;
	{8'd250,8'd72} : s = 37;
	{8'd250,8'd73} : s = 135;
	{8'd250,8'd74} : s = 35;
	{8'd250,8'd75} : s = 120;
	{8'd250,8'd76} : s = 116;
	{8'd250,8'd77} : s = 244;
	{8'd250,8'd78} : s = 28;
	{8'd250,8'd79} : s = 114;
	{8'd250,8'd80} : s = 113;
	{8'd250,8'd81} : s = 242;
	{8'd250,8'd82} : s = 108;
	{8'd250,8'd83} : s = 241;
	{8'd250,8'd84} : s = 236;
	{8'd250,8'd85} : s = 399;
	{8'd250,8'd86} : s = 26;
	{8'd250,8'd87} : s = 106;
	{8'd250,8'd88} : s = 105;
	{8'd250,8'd89} : s = 234;
	{8'd250,8'd90} : s = 102;
	{8'd250,8'd91} : s = 233;
	{8'd250,8'd92} : s = 230;
	{8'd250,8'd93} : s = 380;
	{8'd250,8'd94} : s = 101;
	{8'd250,8'd95} : s = 229;
	{8'd250,8'd96} : s = 227;
	{8'd250,8'd97} : s = 378;
	{8'd250,8'd98} : s = 220;
	{8'd250,8'd99} : s = 377;
	{8'd250,8'd100} : s = 374;
	{8'd250,8'd101} : s = 487;
	{8'd250,8'd102} : s = 25;
	{8'd250,8'd103} : s = 99;
	{8'd250,8'd104} : s = 92;
	{8'd250,8'd105} : s = 218;
	{8'd250,8'd106} : s = 90;
	{8'd250,8'd107} : s = 217;
	{8'd250,8'd108} : s = 214;
	{8'd250,8'd109} : s = 373;
	{8'd250,8'd110} : s = 89;
	{8'd250,8'd111} : s = 213;
	{8'd250,8'd112} : s = 211;
	{8'd250,8'd113} : s = 371;
	{8'd250,8'd114} : s = 206;
	{8'd250,8'd115} : s = 366;
	{8'd250,8'd116} : s = 365;
	{8'd250,8'd117} : s = 478;
	{8'd250,8'd118} : s = 86;
	{8'd250,8'd119} : s = 205;
	{8'd250,8'd120} : s = 203;
	{8'd250,8'd121} : s = 363;
	{8'd250,8'd122} : s = 199;
	{8'd250,8'd123} : s = 359;
	{8'd250,8'd124} : s = 350;
	{8'd250,8'd125} : s = 477;
	{8'd250,8'd126} : s = 188;
	{8'd250,8'd127} : s = 349;
	{8'd250,8'd128} : s = 347;
	{8'd250,8'd129} : s = 475;
	{8'd250,8'd130} : s = 343;
	{8'd250,8'd131} : s = 471;
	{8'd250,8'd132} : s = 463;
	{8'd250,8'd133} : s = 509;
	{8'd250,8'd134} : s = 3;
	{8'd250,8'd135} : s = 22;
	{8'd250,8'd136} : s = 21;
	{8'd250,8'd137} : s = 85;
	{8'd250,8'd138} : s = 19;
	{8'd250,8'd139} : s = 83;
	{8'd250,8'd140} : s = 78;
	{8'd250,8'd141} : s = 186;
	{8'd250,8'd142} : s = 14;
	{8'd250,8'd143} : s = 77;
	{8'd250,8'd144} : s = 75;
	{8'd250,8'd145} : s = 185;
	{8'd250,8'd146} : s = 71;
	{8'd250,8'd147} : s = 182;
	{8'd250,8'd148} : s = 181;
	{8'd250,8'd149} : s = 335;
	{8'd250,8'd150} : s = 13;
	{8'd250,8'd151} : s = 60;
	{8'd250,8'd152} : s = 58;
	{8'd250,8'd153} : s = 179;
	{8'd250,8'd154} : s = 57;
	{8'd250,8'd155} : s = 174;
	{8'd250,8'd156} : s = 173;
	{8'd250,8'd157} : s = 318;
	{8'd250,8'd158} : s = 54;
	{8'd250,8'd159} : s = 171;
	{8'd250,8'd160} : s = 167;
	{8'd250,8'd161} : s = 317;
	{8'd250,8'd162} : s = 158;
	{8'd250,8'd163} : s = 315;
	{8'd250,8'd164} : s = 311;
	{8'd250,8'd165} : s = 446;
	{8'd250,8'd166} : s = 11;
	{8'd250,8'd167} : s = 53;
	{8'd250,8'd168} : s = 51;
	{8'd250,8'd169} : s = 157;
	{8'd250,8'd170} : s = 46;
	{8'd250,8'd171} : s = 155;
	{8'd250,8'd172} : s = 151;
	{8'd250,8'd173} : s = 303;
	{8'd250,8'd174} : s = 45;
	{8'd250,8'd175} : s = 143;
	{8'd250,8'd176} : s = 124;
	{8'd250,8'd177} : s = 287;
	{8'd250,8'd178} : s = 122;
	{8'd250,8'd179} : s = 252;
	{8'd250,8'd180} : s = 250;
	{8'd250,8'd181} : s = 445;
	{8'd250,8'd182} : s = 43;
	{8'd250,8'd183} : s = 121;
	{8'd250,8'd184} : s = 118;
	{8'd250,8'd185} : s = 249;
	{8'd250,8'd186} : s = 117;
	{8'd250,8'd187} : s = 246;
	{8'd250,8'd188} : s = 245;
	{8'd250,8'd189} : s = 443;
	{8'd250,8'd190} : s = 115;
	{8'd250,8'd191} : s = 243;
	{8'd250,8'd192} : s = 238;
	{8'd250,8'd193} : s = 439;
	{8'd250,8'd194} : s = 237;
	{8'd250,8'd195} : s = 431;
	{8'd250,8'd196} : s = 415;
	{8'd250,8'd197} : s = 507;
	{8'd250,8'd198} : s = 7;
	{8'd250,8'd199} : s = 39;
	{8'd250,8'd200} : s = 30;
	{8'd250,8'd201} : s = 110;
	{8'd250,8'd202} : s = 29;
	{8'd250,8'd203} : s = 109;
	{8'd250,8'd204} : s = 107;
	{8'd250,8'd205} : s = 235;
	{8'd250,8'd206} : s = 27;
	{8'd250,8'd207} : s = 103;
	{8'd250,8'd208} : s = 94;
	{8'd250,8'd209} : s = 231;
	{8'd250,8'd210} : s = 93;
	{8'd250,8'd211} : s = 222;
	{8'd250,8'd212} : s = 221;
	{8'd250,8'd213} : s = 382;
	{8'd250,8'd214} : s = 23;
	{8'd250,8'd215} : s = 91;
	{8'd250,8'd216} : s = 87;
	{8'd250,8'd217} : s = 219;
	{8'd250,8'd218} : s = 79;
	{8'd250,8'd219} : s = 215;
	{8'd250,8'd220} : s = 207;
	{8'd250,8'd221} : s = 381;
	{8'd250,8'd222} : s = 62;
	{8'd250,8'd223} : s = 190;
	{8'd250,8'd224} : s = 189;
	{8'd250,8'd225} : s = 379;
	{8'd250,8'd226} : s = 187;
	{8'd250,8'd227} : s = 375;
	{8'd250,8'd228} : s = 367;
	{8'd250,8'd229} : s = 503;
	{8'd250,8'd230} : s = 15;
	{8'd250,8'd231} : s = 61;
	{8'd250,8'd232} : s = 59;
	{8'd250,8'd233} : s = 183;
	{8'd250,8'd234} : s = 55;
	{8'd250,8'd235} : s = 175;
	{8'd250,8'd236} : s = 159;
	{8'd250,8'd237} : s = 351;
	{8'd250,8'd238} : s = 47;
	{8'd250,8'd239} : s = 126;
	{8'd250,8'd240} : s = 125;
	{8'd250,8'd241} : s = 319;
	{8'd250,8'd242} : s = 123;
	{8'd250,8'd243} : s = 254;
	{8'd250,8'd244} : s = 253;
	{8'd250,8'd245} : s = 479;
	{8'd250,8'd246} : s = 31;
	{8'd250,8'd247} : s = 119;
	{8'd250,8'd248} : s = 111;
	{8'd250,8'd249} : s = 251;
	{8'd250,8'd250} : s = 95;
	{8'd250,8'd251} : s = 247;
	{8'd250,8'd252} : s = 239;
	{8'd250,8'd253} : s = 495;
	{8'd250,8'd254} : s = 63;
	{8'd250,8'd255} : s = 223;
	{8'd251,8'd0} : s = 499;
	{8'd251,8'd1} : s = 429;
	{8'd251,8'd2} : s = 494;
	{8'd251,8'd3} : s = 493;
	{8'd251,8'd4} : s = 510;
	{8'd251,8'd5} : s = 1;
	{8'd251,8'd6} : s = 18;
	{8'd251,8'd7} : s = 17;
	{8'd251,8'd8} : s = 82;
	{8'd251,8'd9} : s = 12;
	{8'd251,8'd10} : s = 81;
	{8'd251,8'd11} : s = 76;
	{8'd251,8'd12} : s = 195;
	{8'd251,8'd13} : s = 10;
	{8'd251,8'd14} : s = 74;
	{8'd251,8'd15} : s = 73;
	{8'd251,8'd16} : s = 184;
	{8'd251,8'd17} : s = 70;
	{8'd251,8'd18} : s = 180;
	{8'd251,8'd19} : s = 178;
	{8'd251,8'd20} : s = 314;
	{8'd251,8'd21} : s = 9;
	{8'd251,8'd22} : s = 69;
	{8'd251,8'd23} : s = 67;
	{8'd251,8'd24} : s = 177;
	{8'd251,8'd25} : s = 56;
	{8'd251,8'd26} : s = 172;
	{8'd251,8'd27} : s = 170;
	{8'd251,8'd28} : s = 313;
	{8'd251,8'd29} : s = 52;
	{8'd251,8'd30} : s = 169;
	{8'd251,8'd31} : s = 166;
	{8'd251,8'd32} : s = 310;
	{8'd251,8'd33} : s = 165;
	{8'd251,8'd34} : s = 309;
	{8'd251,8'd35} : s = 307;
	{8'd251,8'd36} : s = 427;
	{8'd251,8'd37} : s = 6;
	{8'd251,8'd38} : s = 50;
	{8'd251,8'd39} : s = 49;
	{8'd251,8'd40} : s = 163;
	{8'd251,8'd41} : s = 44;
	{8'd251,8'd42} : s = 156;
	{8'd251,8'd43} : s = 154;
	{8'd251,8'd44} : s = 302;
	{8'd251,8'd45} : s = 42;
	{8'd251,8'd46} : s = 153;
	{8'd251,8'd47} : s = 150;
	{8'd251,8'd48} : s = 301;
	{8'd251,8'd49} : s = 149;
	{8'd251,8'd50} : s = 299;
	{8'd251,8'd51} : s = 295;
	{8'd251,8'd52} : s = 423;
	{8'd251,8'd53} : s = 41;
	{8'd251,8'd54} : s = 147;
	{8'd251,8'd55} : s = 142;
	{8'd251,8'd56} : s = 286;
	{8'd251,8'd57} : s = 141;
	{8'd251,8'd58} : s = 285;
	{8'd251,8'd59} : s = 283;
	{8'd251,8'd60} : s = 414;
	{8'd251,8'd61} : s = 139;
	{8'd251,8'd62} : s = 279;
	{8'd251,8'd63} : s = 271;
	{8'd251,8'd64} : s = 413;
	{8'd251,8'd65} : s = 248;
	{8'd251,8'd66} : s = 411;
	{8'd251,8'd67} : s = 407;
	{8'd251,8'd68} : s = 491;
	{8'd251,8'd69} : s = 5;
	{8'd251,8'd70} : s = 38;
	{8'd251,8'd71} : s = 37;
	{8'd251,8'd72} : s = 135;
	{8'd251,8'd73} : s = 35;
	{8'd251,8'd74} : s = 120;
	{8'd251,8'd75} : s = 116;
	{8'd251,8'd76} : s = 244;
	{8'd251,8'd77} : s = 28;
	{8'd251,8'd78} : s = 114;
	{8'd251,8'd79} : s = 113;
	{8'd251,8'd80} : s = 242;
	{8'd251,8'd81} : s = 108;
	{8'd251,8'd82} : s = 241;
	{8'd251,8'd83} : s = 236;
	{8'd251,8'd84} : s = 399;
	{8'd251,8'd85} : s = 26;
	{8'd251,8'd86} : s = 106;
	{8'd251,8'd87} : s = 105;
	{8'd251,8'd88} : s = 234;
	{8'd251,8'd89} : s = 102;
	{8'd251,8'd90} : s = 233;
	{8'd251,8'd91} : s = 230;
	{8'd251,8'd92} : s = 380;
	{8'd251,8'd93} : s = 101;
	{8'd251,8'd94} : s = 229;
	{8'd251,8'd95} : s = 227;
	{8'd251,8'd96} : s = 378;
	{8'd251,8'd97} : s = 220;
	{8'd251,8'd98} : s = 377;
	{8'd251,8'd99} : s = 374;
	{8'd251,8'd100} : s = 487;
	{8'd251,8'd101} : s = 25;
	{8'd251,8'd102} : s = 99;
	{8'd251,8'd103} : s = 92;
	{8'd251,8'd104} : s = 218;
	{8'd251,8'd105} : s = 90;
	{8'd251,8'd106} : s = 217;
	{8'd251,8'd107} : s = 214;
	{8'd251,8'd108} : s = 373;
	{8'd251,8'd109} : s = 89;
	{8'd251,8'd110} : s = 213;
	{8'd251,8'd111} : s = 211;
	{8'd251,8'd112} : s = 371;
	{8'd251,8'd113} : s = 206;
	{8'd251,8'd114} : s = 366;
	{8'd251,8'd115} : s = 365;
	{8'd251,8'd116} : s = 478;
	{8'd251,8'd117} : s = 86;
	{8'd251,8'd118} : s = 205;
	{8'd251,8'd119} : s = 203;
	{8'd251,8'd120} : s = 363;
	{8'd251,8'd121} : s = 199;
	{8'd251,8'd122} : s = 359;
	{8'd251,8'd123} : s = 350;
	{8'd251,8'd124} : s = 477;
	{8'd251,8'd125} : s = 188;
	{8'd251,8'd126} : s = 349;
	{8'd251,8'd127} : s = 347;
	{8'd251,8'd128} : s = 475;
	{8'd251,8'd129} : s = 343;
	{8'd251,8'd130} : s = 471;
	{8'd251,8'd131} : s = 463;
	{8'd251,8'd132} : s = 509;
	{8'd251,8'd133} : s = 3;
	{8'd251,8'd134} : s = 22;
	{8'd251,8'd135} : s = 21;
	{8'd251,8'd136} : s = 85;
	{8'd251,8'd137} : s = 19;
	{8'd251,8'd138} : s = 83;
	{8'd251,8'd139} : s = 78;
	{8'd251,8'd140} : s = 186;
	{8'd251,8'd141} : s = 14;
	{8'd251,8'd142} : s = 77;
	{8'd251,8'd143} : s = 75;
	{8'd251,8'd144} : s = 185;
	{8'd251,8'd145} : s = 71;
	{8'd251,8'd146} : s = 182;
	{8'd251,8'd147} : s = 181;
	{8'd251,8'd148} : s = 335;
	{8'd251,8'd149} : s = 13;
	{8'd251,8'd150} : s = 60;
	{8'd251,8'd151} : s = 58;
	{8'd251,8'd152} : s = 179;
	{8'd251,8'd153} : s = 57;
	{8'd251,8'd154} : s = 174;
	{8'd251,8'd155} : s = 173;
	{8'd251,8'd156} : s = 318;
	{8'd251,8'd157} : s = 54;
	{8'd251,8'd158} : s = 171;
	{8'd251,8'd159} : s = 167;
	{8'd251,8'd160} : s = 317;
	{8'd251,8'd161} : s = 158;
	{8'd251,8'd162} : s = 315;
	{8'd251,8'd163} : s = 311;
	{8'd251,8'd164} : s = 446;
	{8'd251,8'd165} : s = 11;
	{8'd251,8'd166} : s = 53;
	{8'd251,8'd167} : s = 51;
	{8'd251,8'd168} : s = 157;
	{8'd251,8'd169} : s = 46;
	{8'd251,8'd170} : s = 155;
	{8'd251,8'd171} : s = 151;
	{8'd251,8'd172} : s = 303;
	{8'd251,8'd173} : s = 45;
	{8'd251,8'd174} : s = 143;
	{8'd251,8'd175} : s = 124;
	{8'd251,8'd176} : s = 287;
	{8'd251,8'd177} : s = 122;
	{8'd251,8'd178} : s = 252;
	{8'd251,8'd179} : s = 250;
	{8'd251,8'd180} : s = 445;
	{8'd251,8'd181} : s = 43;
	{8'd251,8'd182} : s = 121;
	{8'd251,8'd183} : s = 118;
	{8'd251,8'd184} : s = 249;
	{8'd251,8'd185} : s = 117;
	{8'd251,8'd186} : s = 246;
	{8'd251,8'd187} : s = 245;
	{8'd251,8'd188} : s = 443;
	{8'd251,8'd189} : s = 115;
	{8'd251,8'd190} : s = 243;
	{8'd251,8'd191} : s = 238;
	{8'd251,8'd192} : s = 439;
	{8'd251,8'd193} : s = 237;
	{8'd251,8'd194} : s = 431;
	{8'd251,8'd195} : s = 415;
	{8'd251,8'd196} : s = 507;
	{8'd251,8'd197} : s = 7;
	{8'd251,8'd198} : s = 39;
	{8'd251,8'd199} : s = 30;
	{8'd251,8'd200} : s = 110;
	{8'd251,8'd201} : s = 29;
	{8'd251,8'd202} : s = 109;
	{8'd251,8'd203} : s = 107;
	{8'd251,8'd204} : s = 235;
	{8'd251,8'd205} : s = 27;
	{8'd251,8'd206} : s = 103;
	{8'd251,8'd207} : s = 94;
	{8'd251,8'd208} : s = 231;
	{8'd251,8'd209} : s = 93;
	{8'd251,8'd210} : s = 222;
	{8'd251,8'd211} : s = 221;
	{8'd251,8'd212} : s = 382;
	{8'd251,8'd213} : s = 23;
	{8'd251,8'd214} : s = 91;
	{8'd251,8'd215} : s = 87;
	{8'd251,8'd216} : s = 219;
	{8'd251,8'd217} : s = 79;
	{8'd251,8'd218} : s = 215;
	{8'd251,8'd219} : s = 207;
	{8'd251,8'd220} : s = 381;
	{8'd251,8'd221} : s = 62;
	{8'd251,8'd222} : s = 190;
	{8'd251,8'd223} : s = 189;
	{8'd251,8'd224} : s = 379;
	{8'd251,8'd225} : s = 187;
	{8'd251,8'd226} : s = 375;
	{8'd251,8'd227} : s = 367;
	{8'd251,8'd228} : s = 503;
	{8'd251,8'd229} : s = 15;
	{8'd251,8'd230} : s = 61;
	{8'd251,8'd231} : s = 59;
	{8'd251,8'd232} : s = 183;
	{8'd251,8'd233} : s = 55;
	{8'd251,8'd234} : s = 175;
	{8'd251,8'd235} : s = 159;
	{8'd251,8'd236} : s = 351;
	{8'd251,8'd237} : s = 47;
	{8'd251,8'd238} : s = 126;
	{8'd251,8'd239} : s = 125;
	{8'd251,8'd240} : s = 319;
	{8'd251,8'd241} : s = 123;
	{8'd251,8'd242} : s = 254;
	{8'd251,8'd243} : s = 253;
	{8'd251,8'd244} : s = 479;
	{8'd251,8'd245} : s = 31;
	{8'd251,8'd246} : s = 119;
	{8'd251,8'd247} : s = 111;
	{8'd251,8'd248} : s = 251;
	{8'd251,8'd249} : s = 95;
	{8'd251,8'd250} : s = 247;
	{8'd251,8'd251} : s = 239;
	{8'd251,8'd252} : s = 495;
	{8'd251,8'd253} : s = 63;
	{8'd251,8'd254} : s = 223;
	{8'd251,8'd255} : s = 191;
	{8'd252,8'd0} : s = 429;
	{8'd252,8'd1} : s = 494;
	{8'd252,8'd2} : s = 493;
	{8'd252,8'd3} : s = 510;
	{8'd252,8'd4} : s = 1;
	{8'd252,8'd5} : s = 18;
	{8'd252,8'd6} : s = 17;
	{8'd252,8'd7} : s = 82;
	{8'd252,8'd8} : s = 12;
	{8'd252,8'd9} : s = 81;
	{8'd252,8'd10} : s = 76;
	{8'd252,8'd11} : s = 195;
	{8'd252,8'd12} : s = 10;
	{8'd252,8'd13} : s = 74;
	{8'd252,8'd14} : s = 73;
	{8'd252,8'd15} : s = 184;
	{8'd252,8'd16} : s = 70;
	{8'd252,8'd17} : s = 180;
	{8'd252,8'd18} : s = 178;
	{8'd252,8'd19} : s = 314;
	{8'd252,8'd20} : s = 9;
	{8'd252,8'd21} : s = 69;
	{8'd252,8'd22} : s = 67;
	{8'd252,8'd23} : s = 177;
	{8'd252,8'd24} : s = 56;
	{8'd252,8'd25} : s = 172;
	{8'd252,8'd26} : s = 170;
	{8'd252,8'd27} : s = 313;
	{8'd252,8'd28} : s = 52;
	{8'd252,8'd29} : s = 169;
	{8'd252,8'd30} : s = 166;
	{8'd252,8'd31} : s = 310;
	{8'd252,8'd32} : s = 165;
	{8'd252,8'd33} : s = 309;
	{8'd252,8'd34} : s = 307;
	{8'd252,8'd35} : s = 427;
	{8'd252,8'd36} : s = 6;
	{8'd252,8'd37} : s = 50;
	{8'd252,8'd38} : s = 49;
	{8'd252,8'd39} : s = 163;
	{8'd252,8'd40} : s = 44;
	{8'd252,8'd41} : s = 156;
	{8'd252,8'd42} : s = 154;
	{8'd252,8'd43} : s = 302;
	{8'd252,8'd44} : s = 42;
	{8'd252,8'd45} : s = 153;
	{8'd252,8'd46} : s = 150;
	{8'd252,8'd47} : s = 301;
	{8'd252,8'd48} : s = 149;
	{8'd252,8'd49} : s = 299;
	{8'd252,8'd50} : s = 295;
	{8'd252,8'd51} : s = 423;
	{8'd252,8'd52} : s = 41;
	{8'd252,8'd53} : s = 147;
	{8'd252,8'd54} : s = 142;
	{8'd252,8'd55} : s = 286;
	{8'd252,8'd56} : s = 141;
	{8'd252,8'd57} : s = 285;
	{8'd252,8'd58} : s = 283;
	{8'd252,8'd59} : s = 414;
	{8'd252,8'd60} : s = 139;
	{8'd252,8'd61} : s = 279;
	{8'd252,8'd62} : s = 271;
	{8'd252,8'd63} : s = 413;
	{8'd252,8'd64} : s = 248;
	{8'd252,8'd65} : s = 411;
	{8'd252,8'd66} : s = 407;
	{8'd252,8'd67} : s = 491;
	{8'd252,8'd68} : s = 5;
	{8'd252,8'd69} : s = 38;
	{8'd252,8'd70} : s = 37;
	{8'd252,8'd71} : s = 135;
	{8'd252,8'd72} : s = 35;
	{8'd252,8'd73} : s = 120;
	{8'd252,8'd74} : s = 116;
	{8'd252,8'd75} : s = 244;
	{8'd252,8'd76} : s = 28;
	{8'd252,8'd77} : s = 114;
	{8'd252,8'd78} : s = 113;
	{8'd252,8'd79} : s = 242;
	{8'd252,8'd80} : s = 108;
	{8'd252,8'd81} : s = 241;
	{8'd252,8'd82} : s = 236;
	{8'd252,8'd83} : s = 399;
	{8'd252,8'd84} : s = 26;
	{8'd252,8'd85} : s = 106;
	{8'd252,8'd86} : s = 105;
	{8'd252,8'd87} : s = 234;
	{8'd252,8'd88} : s = 102;
	{8'd252,8'd89} : s = 233;
	{8'd252,8'd90} : s = 230;
	{8'd252,8'd91} : s = 380;
	{8'd252,8'd92} : s = 101;
	{8'd252,8'd93} : s = 229;
	{8'd252,8'd94} : s = 227;
	{8'd252,8'd95} : s = 378;
	{8'd252,8'd96} : s = 220;
	{8'd252,8'd97} : s = 377;
	{8'd252,8'd98} : s = 374;
	{8'd252,8'd99} : s = 487;
	{8'd252,8'd100} : s = 25;
	{8'd252,8'd101} : s = 99;
	{8'd252,8'd102} : s = 92;
	{8'd252,8'd103} : s = 218;
	{8'd252,8'd104} : s = 90;
	{8'd252,8'd105} : s = 217;
	{8'd252,8'd106} : s = 214;
	{8'd252,8'd107} : s = 373;
	{8'd252,8'd108} : s = 89;
	{8'd252,8'd109} : s = 213;
	{8'd252,8'd110} : s = 211;
	{8'd252,8'd111} : s = 371;
	{8'd252,8'd112} : s = 206;
	{8'd252,8'd113} : s = 366;
	{8'd252,8'd114} : s = 365;
	{8'd252,8'd115} : s = 478;
	{8'd252,8'd116} : s = 86;
	{8'd252,8'd117} : s = 205;
	{8'd252,8'd118} : s = 203;
	{8'd252,8'd119} : s = 363;
	{8'd252,8'd120} : s = 199;
	{8'd252,8'd121} : s = 359;
	{8'd252,8'd122} : s = 350;
	{8'd252,8'd123} : s = 477;
	{8'd252,8'd124} : s = 188;
	{8'd252,8'd125} : s = 349;
	{8'd252,8'd126} : s = 347;
	{8'd252,8'd127} : s = 475;
	{8'd252,8'd128} : s = 343;
	{8'd252,8'd129} : s = 471;
	{8'd252,8'd130} : s = 463;
	{8'd252,8'd131} : s = 509;
	{8'd252,8'd132} : s = 3;
	{8'd252,8'd133} : s = 22;
	{8'd252,8'd134} : s = 21;
	{8'd252,8'd135} : s = 85;
	{8'd252,8'd136} : s = 19;
	{8'd252,8'd137} : s = 83;
	{8'd252,8'd138} : s = 78;
	{8'd252,8'd139} : s = 186;
	{8'd252,8'd140} : s = 14;
	{8'd252,8'd141} : s = 77;
	{8'd252,8'd142} : s = 75;
	{8'd252,8'd143} : s = 185;
	{8'd252,8'd144} : s = 71;
	{8'd252,8'd145} : s = 182;
	{8'd252,8'd146} : s = 181;
	{8'd252,8'd147} : s = 335;
	{8'd252,8'd148} : s = 13;
	{8'd252,8'd149} : s = 60;
	{8'd252,8'd150} : s = 58;
	{8'd252,8'd151} : s = 179;
	{8'd252,8'd152} : s = 57;
	{8'd252,8'd153} : s = 174;
	{8'd252,8'd154} : s = 173;
	{8'd252,8'd155} : s = 318;
	{8'd252,8'd156} : s = 54;
	{8'd252,8'd157} : s = 171;
	{8'd252,8'd158} : s = 167;
	{8'd252,8'd159} : s = 317;
	{8'd252,8'd160} : s = 158;
	{8'd252,8'd161} : s = 315;
	{8'd252,8'd162} : s = 311;
	{8'd252,8'd163} : s = 446;
	{8'd252,8'd164} : s = 11;
	{8'd252,8'd165} : s = 53;
	{8'd252,8'd166} : s = 51;
	{8'd252,8'd167} : s = 157;
	{8'd252,8'd168} : s = 46;
	{8'd252,8'd169} : s = 155;
	{8'd252,8'd170} : s = 151;
	{8'd252,8'd171} : s = 303;
	{8'd252,8'd172} : s = 45;
	{8'd252,8'd173} : s = 143;
	{8'd252,8'd174} : s = 124;
	{8'd252,8'd175} : s = 287;
	{8'd252,8'd176} : s = 122;
	{8'd252,8'd177} : s = 252;
	{8'd252,8'd178} : s = 250;
	{8'd252,8'd179} : s = 445;
	{8'd252,8'd180} : s = 43;
	{8'd252,8'd181} : s = 121;
	{8'd252,8'd182} : s = 118;
	{8'd252,8'd183} : s = 249;
	{8'd252,8'd184} : s = 117;
	{8'd252,8'd185} : s = 246;
	{8'd252,8'd186} : s = 245;
	{8'd252,8'd187} : s = 443;
	{8'd252,8'd188} : s = 115;
	{8'd252,8'd189} : s = 243;
	{8'd252,8'd190} : s = 238;
	{8'd252,8'd191} : s = 439;
	{8'd252,8'd192} : s = 237;
	{8'd252,8'd193} : s = 431;
	{8'd252,8'd194} : s = 415;
	{8'd252,8'd195} : s = 507;
	{8'd252,8'd196} : s = 7;
	{8'd252,8'd197} : s = 39;
	{8'd252,8'd198} : s = 30;
	{8'd252,8'd199} : s = 110;
	{8'd252,8'd200} : s = 29;
	{8'd252,8'd201} : s = 109;
	{8'd252,8'd202} : s = 107;
	{8'd252,8'd203} : s = 235;
	{8'd252,8'd204} : s = 27;
	{8'd252,8'd205} : s = 103;
	{8'd252,8'd206} : s = 94;
	{8'd252,8'd207} : s = 231;
	{8'd252,8'd208} : s = 93;
	{8'd252,8'd209} : s = 222;
	{8'd252,8'd210} : s = 221;
	{8'd252,8'd211} : s = 382;
	{8'd252,8'd212} : s = 23;
	{8'd252,8'd213} : s = 91;
	{8'd252,8'd214} : s = 87;
	{8'd252,8'd215} : s = 219;
	{8'd252,8'd216} : s = 79;
	{8'd252,8'd217} : s = 215;
	{8'd252,8'd218} : s = 207;
	{8'd252,8'd219} : s = 381;
	{8'd252,8'd220} : s = 62;
	{8'd252,8'd221} : s = 190;
	{8'd252,8'd222} : s = 189;
	{8'd252,8'd223} : s = 379;
	{8'd252,8'd224} : s = 187;
	{8'd252,8'd225} : s = 375;
	{8'd252,8'd226} : s = 367;
	{8'd252,8'd227} : s = 503;
	{8'd252,8'd228} : s = 15;
	{8'd252,8'd229} : s = 61;
	{8'd252,8'd230} : s = 59;
	{8'd252,8'd231} : s = 183;
	{8'd252,8'd232} : s = 55;
	{8'd252,8'd233} : s = 175;
	{8'd252,8'd234} : s = 159;
	{8'd252,8'd235} : s = 351;
	{8'd252,8'd236} : s = 47;
	{8'd252,8'd237} : s = 126;
	{8'd252,8'd238} : s = 125;
	{8'd252,8'd239} : s = 319;
	{8'd252,8'd240} : s = 123;
	{8'd252,8'd241} : s = 254;
	{8'd252,8'd242} : s = 253;
	{8'd252,8'd243} : s = 479;
	{8'd252,8'd244} : s = 31;
	{8'd252,8'd245} : s = 119;
	{8'd252,8'd246} : s = 111;
	{8'd252,8'd247} : s = 251;
	{8'd252,8'd248} : s = 95;
	{8'd252,8'd249} : s = 247;
	{8'd252,8'd250} : s = 239;
	{8'd252,8'd251} : s = 495;
	{8'd252,8'd252} : s = 63;
	{8'd252,8'd253} : s = 223;
	{8'd252,8'd254} : s = 191;
	{8'd252,8'd255} : s = 447;
	{8'd253,8'd0} : s = 494;
	{8'd253,8'd1} : s = 493;
	{8'd253,8'd2} : s = 510;
	{8'd253,8'd3} : s = 1;
	{8'd253,8'd4} : s = 18;
	{8'd253,8'd5} : s = 17;
	{8'd253,8'd6} : s = 82;
	{8'd253,8'd7} : s = 12;
	{8'd253,8'd8} : s = 81;
	{8'd253,8'd9} : s = 76;
	{8'd253,8'd10} : s = 195;
	{8'd253,8'd11} : s = 10;
	{8'd253,8'd12} : s = 74;
	{8'd253,8'd13} : s = 73;
	{8'd253,8'd14} : s = 184;
	{8'd253,8'd15} : s = 70;
	{8'd253,8'd16} : s = 180;
	{8'd253,8'd17} : s = 178;
	{8'd253,8'd18} : s = 314;
	{8'd253,8'd19} : s = 9;
	{8'd253,8'd20} : s = 69;
	{8'd253,8'd21} : s = 67;
	{8'd253,8'd22} : s = 177;
	{8'd253,8'd23} : s = 56;
	{8'd253,8'd24} : s = 172;
	{8'd253,8'd25} : s = 170;
	{8'd253,8'd26} : s = 313;
	{8'd253,8'd27} : s = 52;
	{8'd253,8'd28} : s = 169;
	{8'd253,8'd29} : s = 166;
	{8'd253,8'd30} : s = 310;
	{8'd253,8'd31} : s = 165;
	{8'd253,8'd32} : s = 309;
	{8'd253,8'd33} : s = 307;
	{8'd253,8'd34} : s = 427;
	{8'd253,8'd35} : s = 6;
	{8'd253,8'd36} : s = 50;
	{8'd253,8'd37} : s = 49;
	{8'd253,8'd38} : s = 163;
	{8'd253,8'd39} : s = 44;
	{8'd253,8'd40} : s = 156;
	{8'd253,8'd41} : s = 154;
	{8'd253,8'd42} : s = 302;
	{8'd253,8'd43} : s = 42;
	{8'd253,8'd44} : s = 153;
	{8'd253,8'd45} : s = 150;
	{8'd253,8'd46} : s = 301;
	{8'd253,8'd47} : s = 149;
	{8'd253,8'd48} : s = 299;
	{8'd253,8'd49} : s = 295;
	{8'd253,8'd50} : s = 423;
	{8'd253,8'd51} : s = 41;
	{8'd253,8'd52} : s = 147;
	{8'd253,8'd53} : s = 142;
	{8'd253,8'd54} : s = 286;
	{8'd253,8'd55} : s = 141;
	{8'd253,8'd56} : s = 285;
	{8'd253,8'd57} : s = 283;
	{8'd253,8'd58} : s = 414;
	{8'd253,8'd59} : s = 139;
	{8'd253,8'd60} : s = 279;
	{8'd253,8'd61} : s = 271;
	{8'd253,8'd62} : s = 413;
	{8'd253,8'd63} : s = 248;
	{8'd253,8'd64} : s = 411;
	{8'd253,8'd65} : s = 407;
	{8'd253,8'd66} : s = 491;
	{8'd253,8'd67} : s = 5;
	{8'd253,8'd68} : s = 38;
	{8'd253,8'd69} : s = 37;
	{8'd253,8'd70} : s = 135;
	{8'd253,8'd71} : s = 35;
	{8'd253,8'd72} : s = 120;
	{8'd253,8'd73} : s = 116;
	{8'd253,8'd74} : s = 244;
	{8'd253,8'd75} : s = 28;
	{8'd253,8'd76} : s = 114;
	{8'd253,8'd77} : s = 113;
	{8'd253,8'd78} : s = 242;
	{8'd253,8'd79} : s = 108;
	{8'd253,8'd80} : s = 241;
	{8'd253,8'd81} : s = 236;
	{8'd253,8'd82} : s = 399;
	{8'd253,8'd83} : s = 26;
	{8'd253,8'd84} : s = 106;
	{8'd253,8'd85} : s = 105;
	{8'd253,8'd86} : s = 234;
	{8'd253,8'd87} : s = 102;
	{8'd253,8'd88} : s = 233;
	{8'd253,8'd89} : s = 230;
	{8'd253,8'd90} : s = 380;
	{8'd253,8'd91} : s = 101;
	{8'd253,8'd92} : s = 229;
	{8'd253,8'd93} : s = 227;
	{8'd253,8'd94} : s = 378;
	{8'd253,8'd95} : s = 220;
	{8'd253,8'd96} : s = 377;
	{8'd253,8'd97} : s = 374;
	{8'd253,8'd98} : s = 487;
	{8'd253,8'd99} : s = 25;
	{8'd253,8'd100} : s = 99;
	{8'd253,8'd101} : s = 92;
	{8'd253,8'd102} : s = 218;
	{8'd253,8'd103} : s = 90;
	{8'd253,8'd104} : s = 217;
	{8'd253,8'd105} : s = 214;
	{8'd253,8'd106} : s = 373;
	{8'd253,8'd107} : s = 89;
	{8'd253,8'd108} : s = 213;
	{8'd253,8'd109} : s = 211;
	{8'd253,8'd110} : s = 371;
	{8'd253,8'd111} : s = 206;
	{8'd253,8'd112} : s = 366;
	{8'd253,8'd113} : s = 365;
	{8'd253,8'd114} : s = 478;
	{8'd253,8'd115} : s = 86;
	{8'd253,8'd116} : s = 205;
	{8'd253,8'd117} : s = 203;
	{8'd253,8'd118} : s = 363;
	{8'd253,8'd119} : s = 199;
	{8'd253,8'd120} : s = 359;
	{8'd253,8'd121} : s = 350;
	{8'd253,8'd122} : s = 477;
	{8'd253,8'd123} : s = 188;
	{8'd253,8'd124} : s = 349;
	{8'd253,8'd125} : s = 347;
	{8'd253,8'd126} : s = 475;
	{8'd253,8'd127} : s = 343;
	{8'd253,8'd128} : s = 471;
	{8'd253,8'd129} : s = 463;
	{8'd253,8'd130} : s = 509;
	{8'd253,8'd131} : s = 3;
	{8'd253,8'd132} : s = 22;
	{8'd253,8'd133} : s = 21;
	{8'd253,8'd134} : s = 85;
	{8'd253,8'd135} : s = 19;
	{8'd253,8'd136} : s = 83;
	{8'd253,8'd137} : s = 78;
	{8'd253,8'd138} : s = 186;
	{8'd253,8'd139} : s = 14;
	{8'd253,8'd140} : s = 77;
	{8'd253,8'd141} : s = 75;
	{8'd253,8'd142} : s = 185;
	{8'd253,8'd143} : s = 71;
	{8'd253,8'd144} : s = 182;
	{8'd253,8'd145} : s = 181;
	{8'd253,8'd146} : s = 335;
	{8'd253,8'd147} : s = 13;
	{8'd253,8'd148} : s = 60;
	{8'd253,8'd149} : s = 58;
	{8'd253,8'd150} : s = 179;
	{8'd253,8'd151} : s = 57;
	{8'd253,8'd152} : s = 174;
	{8'd253,8'd153} : s = 173;
	{8'd253,8'd154} : s = 318;
	{8'd253,8'd155} : s = 54;
	{8'd253,8'd156} : s = 171;
	{8'd253,8'd157} : s = 167;
	{8'd253,8'd158} : s = 317;
	{8'd253,8'd159} : s = 158;
	{8'd253,8'd160} : s = 315;
	{8'd253,8'd161} : s = 311;
	{8'd253,8'd162} : s = 446;
	{8'd253,8'd163} : s = 11;
	{8'd253,8'd164} : s = 53;
	{8'd253,8'd165} : s = 51;
	{8'd253,8'd166} : s = 157;
	{8'd253,8'd167} : s = 46;
	{8'd253,8'd168} : s = 155;
	{8'd253,8'd169} : s = 151;
	{8'd253,8'd170} : s = 303;
	{8'd253,8'd171} : s = 45;
	{8'd253,8'd172} : s = 143;
	{8'd253,8'd173} : s = 124;
	{8'd253,8'd174} : s = 287;
	{8'd253,8'd175} : s = 122;
	{8'd253,8'd176} : s = 252;
	{8'd253,8'd177} : s = 250;
	{8'd253,8'd178} : s = 445;
	{8'd253,8'd179} : s = 43;
	{8'd253,8'd180} : s = 121;
	{8'd253,8'd181} : s = 118;
	{8'd253,8'd182} : s = 249;
	{8'd253,8'd183} : s = 117;
	{8'd253,8'd184} : s = 246;
	{8'd253,8'd185} : s = 245;
	{8'd253,8'd186} : s = 443;
	{8'd253,8'd187} : s = 115;
	{8'd253,8'd188} : s = 243;
	{8'd253,8'd189} : s = 238;
	{8'd253,8'd190} : s = 439;
	{8'd253,8'd191} : s = 237;
	{8'd253,8'd192} : s = 431;
	{8'd253,8'd193} : s = 415;
	{8'd253,8'd194} : s = 507;
	{8'd253,8'd195} : s = 7;
	{8'd253,8'd196} : s = 39;
	{8'd253,8'd197} : s = 30;
	{8'd253,8'd198} : s = 110;
	{8'd253,8'd199} : s = 29;
	{8'd253,8'd200} : s = 109;
	{8'd253,8'd201} : s = 107;
	{8'd253,8'd202} : s = 235;
	{8'd253,8'd203} : s = 27;
	{8'd253,8'd204} : s = 103;
	{8'd253,8'd205} : s = 94;
	{8'd253,8'd206} : s = 231;
	{8'd253,8'd207} : s = 93;
	{8'd253,8'd208} : s = 222;
	{8'd253,8'd209} : s = 221;
	{8'd253,8'd210} : s = 382;
	{8'd253,8'd211} : s = 23;
	{8'd253,8'd212} : s = 91;
	{8'd253,8'd213} : s = 87;
	{8'd253,8'd214} : s = 219;
	{8'd253,8'd215} : s = 79;
	{8'd253,8'd216} : s = 215;
	{8'd253,8'd217} : s = 207;
	{8'd253,8'd218} : s = 381;
	{8'd253,8'd219} : s = 62;
	{8'd253,8'd220} : s = 190;
	{8'd253,8'd221} : s = 189;
	{8'd253,8'd222} : s = 379;
	{8'd253,8'd223} : s = 187;
	{8'd253,8'd224} : s = 375;
	{8'd253,8'd225} : s = 367;
	{8'd253,8'd226} : s = 503;
	{8'd253,8'd227} : s = 15;
	{8'd253,8'd228} : s = 61;
	{8'd253,8'd229} : s = 59;
	{8'd253,8'd230} : s = 183;
	{8'd253,8'd231} : s = 55;
	{8'd253,8'd232} : s = 175;
	{8'd253,8'd233} : s = 159;
	{8'd253,8'd234} : s = 351;
	{8'd253,8'd235} : s = 47;
	{8'd253,8'd236} : s = 126;
	{8'd253,8'd237} : s = 125;
	{8'd253,8'd238} : s = 319;
	{8'd253,8'd239} : s = 123;
	{8'd253,8'd240} : s = 254;
	{8'd253,8'd241} : s = 253;
	{8'd253,8'd242} : s = 479;
	{8'd253,8'd243} : s = 31;
	{8'd253,8'd244} : s = 119;
	{8'd253,8'd245} : s = 111;
	{8'd253,8'd246} : s = 251;
	{8'd253,8'd247} : s = 95;
	{8'd253,8'd248} : s = 247;
	{8'd253,8'd249} : s = 239;
	{8'd253,8'd250} : s = 495;
	{8'd253,8'd251} : s = 63;
	{8'd253,8'd252} : s = 223;
	{8'd253,8'd253} : s = 191;
	{8'd253,8'd254} : s = 447;
	{8'd253,8'd255} : s = 127;
	{8'd254,8'd0} : s = 493;
	{8'd254,8'd1} : s = 510;
	{8'd254,8'd2} : s = 1;
	{8'd254,8'd3} : s = 18;
	{8'd254,8'd4} : s = 17;
	{8'd254,8'd5} : s = 82;
	{8'd254,8'd6} : s = 12;
	{8'd254,8'd7} : s = 81;
	{8'd254,8'd8} : s = 76;
	{8'd254,8'd9} : s = 195;
	{8'd254,8'd10} : s = 10;
	{8'd254,8'd11} : s = 74;
	{8'd254,8'd12} : s = 73;
	{8'd254,8'd13} : s = 184;
	{8'd254,8'd14} : s = 70;
	{8'd254,8'd15} : s = 180;
	{8'd254,8'd16} : s = 178;
	{8'd254,8'd17} : s = 314;
	{8'd254,8'd18} : s = 9;
	{8'd254,8'd19} : s = 69;
	{8'd254,8'd20} : s = 67;
	{8'd254,8'd21} : s = 177;
	{8'd254,8'd22} : s = 56;
	{8'd254,8'd23} : s = 172;
	{8'd254,8'd24} : s = 170;
	{8'd254,8'd25} : s = 313;
	{8'd254,8'd26} : s = 52;
	{8'd254,8'd27} : s = 169;
	{8'd254,8'd28} : s = 166;
	{8'd254,8'd29} : s = 310;
	{8'd254,8'd30} : s = 165;
	{8'd254,8'd31} : s = 309;
	{8'd254,8'd32} : s = 307;
	{8'd254,8'd33} : s = 427;
	{8'd254,8'd34} : s = 6;
	{8'd254,8'd35} : s = 50;
	{8'd254,8'd36} : s = 49;
	{8'd254,8'd37} : s = 163;
	{8'd254,8'd38} : s = 44;
	{8'd254,8'd39} : s = 156;
	{8'd254,8'd40} : s = 154;
	{8'd254,8'd41} : s = 302;
	{8'd254,8'd42} : s = 42;
	{8'd254,8'd43} : s = 153;
	{8'd254,8'd44} : s = 150;
	{8'd254,8'd45} : s = 301;
	{8'd254,8'd46} : s = 149;
	{8'd254,8'd47} : s = 299;
	{8'd254,8'd48} : s = 295;
	{8'd254,8'd49} : s = 423;
	{8'd254,8'd50} : s = 41;
	{8'd254,8'd51} : s = 147;
	{8'd254,8'd52} : s = 142;
	{8'd254,8'd53} : s = 286;
	{8'd254,8'd54} : s = 141;
	{8'd254,8'd55} : s = 285;
	{8'd254,8'd56} : s = 283;
	{8'd254,8'd57} : s = 414;
	{8'd254,8'd58} : s = 139;
	{8'd254,8'd59} : s = 279;
	{8'd254,8'd60} : s = 271;
	{8'd254,8'd61} : s = 413;
	{8'd254,8'd62} : s = 248;
	{8'd254,8'd63} : s = 411;
	{8'd254,8'd64} : s = 407;
	{8'd254,8'd65} : s = 491;
	{8'd254,8'd66} : s = 5;
	{8'd254,8'd67} : s = 38;
	{8'd254,8'd68} : s = 37;
	{8'd254,8'd69} : s = 135;
	{8'd254,8'd70} : s = 35;
	{8'd254,8'd71} : s = 120;
	{8'd254,8'd72} : s = 116;
	{8'd254,8'd73} : s = 244;
	{8'd254,8'd74} : s = 28;
	{8'd254,8'd75} : s = 114;
	{8'd254,8'd76} : s = 113;
	{8'd254,8'd77} : s = 242;
	{8'd254,8'd78} : s = 108;
	{8'd254,8'd79} : s = 241;
	{8'd254,8'd80} : s = 236;
	{8'd254,8'd81} : s = 399;
	{8'd254,8'd82} : s = 26;
	{8'd254,8'd83} : s = 106;
	{8'd254,8'd84} : s = 105;
	{8'd254,8'd85} : s = 234;
	{8'd254,8'd86} : s = 102;
	{8'd254,8'd87} : s = 233;
	{8'd254,8'd88} : s = 230;
	{8'd254,8'd89} : s = 380;
	{8'd254,8'd90} : s = 101;
	{8'd254,8'd91} : s = 229;
	{8'd254,8'd92} : s = 227;
	{8'd254,8'd93} : s = 378;
	{8'd254,8'd94} : s = 220;
	{8'd254,8'd95} : s = 377;
	{8'd254,8'd96} : s = 374;
	{8'd254,8'd97} : s = 487;
	{8'd254,8'd98} : s = 25;
	{8'd254,8'd99} : s = 99;
	{8'd254,8'd100} : s = 92;
	{8'd254,8'd101} : s = 218;
	{8'd254,8'd102} : s = 90;
	{8'd254,8'd103} : s = 217;
	{8'd254,8'd104} : s = 214;
	{8'd254,8'd105} : s = 373;
	{8'd254,8'd106} : s = 89;
	{8'd254,8'd107} : s = 213;
	{8'd254,8'd108} : s = 211;
	{8'd254,8'd109} : s = 371;
	{8'd254,8'd110} : s = 206;
	{8'd254,8'd111} : s = 366;
	{8'd254,8'd112} : s = 365;
	{8'd254,8'd113} : s = 478;
	{8'd254,8'd114} : s = 86;
	{8'd254,8'd115} : s = 205;
	{8'd254,8'd116} : s = 203;
	{8'd254,8'd117} : s = 363;
	{8'd254,8'd118} : s = 199;
	{8'd254,8'd119} : s = 359;
	{8'd254,8'd120} : s = 350;
	{8'd254,8'd121} : s = 477;
	{8'd254,8'd122} : s = 188;
	{8'd254,8'd123} : s = 349;
	{8'd254,8'd124} : s = 347;
	{8'd254,8'd125} : s = 475;
	{8'd254,8'd126} : s = 343;
	{8'd254,8'd127} : s = 471;
	{8'd254,8'd128} : s = 463;
	{8'd254,8'd129} : s = 509;
	{8'd254,8'd130} : s = 3;
	{8'd254,8'd131} : s = 22;
	{8'd254,8'd132} : s = 21;
	{8'd254,8'd133} : s = 85;
	{8'd254,8'd134} : s = 19;
	{8'd254,8'd135} : s = 83;
	{8'd254,8'd136} : s = 78;
	{8'd254,8'd137} : s = 186;
	{8'd254,8'd138} : s = 14;
	{8'd254,8'd139} : s = 77;
	{8'd254,8'd140} : s = 75;
	{8'd254,8'd141} : s = 185;
	{8'd254,8'd142} : s = 71;
	{8'd254,8'd143} : s = 182;
	{8'd254,8'd144} : s = 181;
	{8'd254,8'd145} : s = 335;
	{8'd254,8'd146} : s = 13;
	{8'd254,8'd147} : s = 60;
	{8'd254,8'd148} : s = 58;
	{8'd254,8'd149} : s = 179;
	{8'd254,8'd150} : s = 57;
	{8'd254,8'd151} : s = 174;
	{8'd254,8'd152} : s = 173;
	{8'd254,8'd153} : s = 318;
	{8'd254,8'd154} : s = 54;
	{8'd254,8'd155} : s = 171;
	{8'd254,8'd156} : s = 167;
	{8'd254,8'd157} : s = 317;
	{8'd254,8'd158} : s = 158;
	{8'd254,8'd159} : s = 315;
	{8'd254,8'd160} : s = 311;
	{8'd254,8'd161} : s = 446;
	{8'd254,8'd162} : s = 11;
	{8'd254,8'd163} : s = 53;
	{8'd254,8'd164} : s = 51;
	{8'd254,8'd165} : s = 157;
	{8'd254,8'd166} : s = 46;
	{8'd254,8'd167} : s = 155;
	{8'd254,8'd168} : s = 151;
	{8'd254,8'd169} : s = 303;
	{8'd254,8'd170} : s = 45;
	{8'd254,8'd171} : s = 143;
	{8'd254,8'd172} : s = 124;
	{8'd254,8'd173} : s = 287;
	{8'd254,8'd174} : s = 122;
	{8'd254,8'd175} : s = 252;
	{8'd254,8'd176} : s = 250;
	{8'd254,8'd177} : s = 445;
	{8'd254,8'd178} : s = 43;
	{8'd254,8'd179} : s = 121;
	{8'd254,8'd180} : s = 118;
	{8'd254,8'd181} : s = 249;
	{8'd254,8'd182} : s = 117;
	{8'd254,8'd183} : s = 246;
	{8'd254,8'd184} : s = 245;
	{8'd254,8'd185} : s = 443;
	{8'd254,8'd186} : s = 115;
	{8'd254,8'd187} : s = 243;
	{8'd254,8'd188} : s = 238;
	{8'd254,8'd189} : s = 439;
	{8'd254,8'd190} : s = 237;
	{8'd254,8'd191} : s = 431;
	{8'd254,8'd192} : s = 415;
	{8'd254,8'd193} : s = 507;
	{8'd254,8'd194} : s = 7;
	{8'd254,8'd195} : s = 39;
	{8'd254,8'd196} : s = 30;
	{8'd254,8'd197} : s = 110;
	{8'd254,8'd198} : s = 29;
	{8'd254,8'd199} : s = 109;
	{8'd254,8'd200} : s = 107;
	{8'd254,8'd201} : s = 235;
	{8'd254,8'd202} : s = 27;
	{8'd254,8'd203} : s = 103;
	{8'd254,8'd204} : s = 94;
	{8'd254,8'd205} : s = 231;
	{8'd254,8'd206} : s = 93;
	{8'd254,8'd207} : s = 222;
	{8'd254,8'd208} : s = 221;
	{8'd254,8'd209} : s = 382;
	{8'd254,8'd210} : s = 23;
	{8'd254,8'd211} : s = 91;
	{8'd254,8'd212} : s = 87;
	{8'd254,8'd213} : s = 219;
	{8'd254,8'd214} : s = 79;
	{8'd254,8'd215} : s = 215;
	{8'd254,8'd216} : s = 207;
	{8'd254,8'd217} : s = 381;
	{8'd254,8'd218} : s = 62;
	{8'd254,8'd219} : s = 190;
	{8'd254,8'd220} : s = 189;
	{8'd254,8'd221} : s = 379;
	{8'd254,8'd222} : s = 187;
	{8'd254,8'd223} : s = 375;
	{8'd254,8'd224} : s = 367;
	{8'd254,8'd225} : s = 503;
	{8'd254,8'd226} : s = 15;
	{8'd254,8'd227} : s = 61;
	{8'd254,8'd228} : s = 59;
	{8'd254,8'd229} : s = 183;
	{8'd254,8'd230} : s = 55;
	{8'd254,8'd231} : s = 175;
	{8'd254,8'd232} : s = 159;
	{8'd254,8'd233} : s = 351;
	{8'd254,8'd234} : s = 47;
	{8'd254,8'd235} : s = 126;
	{8'd254,8'd236} : s = 125;
	{8'd254,8'd237} : s = 319;
	{8'd254,8'd238} : s = 123;
	{8'd254,8'd239} : s = 254;
	{8'd254,8'd240} : s = 253;
	{8'd254,8'd241} : s = 479;
	{8'd254,8'd242} : s = 31;
	{8'd254,8'd243} : s = 119;
	{8'd254,8'd244} : s = 111;
	{8'd254,8'd245} : s = 251;
	{8'd254,8'd246} : s = 95;
	{8'd254,8'd247} : s = 247;
	{8'd254,8'd248} : s = 239;
	{8'd254,8'd249} : s = 495;
	{8'd254,8'd250} : s = 63;
	{8'd254,8'd251} : s = 223;
	{8'd254,8'd252} : s = 191;
	{8'd254,8'd253} : s = 447;
	{8'd254,8'd254} : s = 127;
	{8'd254,8'd255} : s = 383;
	{8'd255,8'd0} : s = 510;
	{8'd255,8'd1} : s = 1;
	{8'd255,8'd2} : s = 18;
	{8'd255,8'd3} : s = 17;
	{8'd255,8'd4} : s = 82;
	{8'd255,8'd5} : s = 12;
	{8'd255,8'd6} : s = 81;
	{8'd255,8'd7} : s = 76;
	{8'd255,8'd8} : s = 195;
	{8'd255,8'd9} : s = 10;
	{8'd255,8'd10} : s = 74;
	{8'd255,8'd11} : s = 73;
	{8'd255,8'd12} : s = 184;
	{8'd255,8'd13} : s = 70;
	{8'd255,8'd14} : s = 180;
	{8'd255,8'd15} : s = 178;
	{8'd255,8'd16} : s = 314;
	{8'd255,8'd17} : s = 9;
	{8'd255,8'd18} : s = 69;
	{8'd255,8'd19} : s = 67;
	{8'd255,8'd20} : s = 177;
	{8'd255,8'd21} : s = 56;
	{8'd255,8'd22} : s = 172;
	{8'd255,8'd23} : s = 170;
	{8'd255,8'd24} : s = 313;
	{8'd255,8'd25} : s = 52;
	{8'd255,8'd26} : s = 169;
	{8'd255,8'd27} : s = 166;
	{8'd255,8'd28} : s = 310;
	{8'd255,8'd29} : s = 165;
	{8'd255,8'd30} : s = 309;
	{8'd255,8'd31} : s = 307;
	{8'd255,8'd32} : s = 427;
	{8'd255,8'd33} : s = 6;
	{8'd255,8'd34} : s = 50;
	{8'd255,8'd35} : s = 49;
	{8'd255,8'd36} : s = 163;
	{8'd255,8'd37} : s = 44;
	{8'd255,8'd38} : s = 156;
	{8'd255,8'd39} : s = 154;
	{8'd255,8'd40} : s = 302;
	{8'd255,8'd41} : s = 42;
	{8'd255,8'd42} : s = 153;
	{8'd255,8'd43} : s = 150;
	{8'd255,8'd44} : s = 301;
	{8'd255,8'd45} : s = 149;
	{8'd255,8'd46} : s = 299;
	{8'd255,8'd47} : s = 295;
	{8'd255,8'd48} : s = 423;
	{8'd255,8'd49} : s = 41;
	{8'd255,8'd50} : s = 147;
	{8'd255,8'd51} : s = 142;
	{8'd255,8'd52} : s = 286;
	{8'd255,8'd53} : s = 141;
	{8'd255,8'd54} : s = 285;
	{8'd255,8'd55} : s = 283;
	{8'd255,8'd56} : s = 414;
	{8'd255,8'd57} : s = 139;
	{8'd255,8'd58} : s = 279;
	{8'd255,8'd59} : s = 271;
	{8'd255,8'd60} : s = 413;
	{8'd255,8'd61} : s = 248;
	{8'd255,8'd62} : s = 411;
	{8'd255,8'd63} : s = 407;
	{8'd255,8'd64} : s = 491;
	{8'd255,8'd65} : s = 5;
	{8'd255,8'd66} : s = 38;
	{8'd255,8'd67} : s = 37;
	{8'd255,8'd68} : s = 135;
	{8'd255,8'd69} : s = 35;
	{8'd255,8'd70} : s = 120;
	{8'd255,8'd71} : s = 116;
	{8'd255,8'd72} : s = 244;
	{8'd255,8'd73} : s = 28;
	{8'd255,8'd74} : s = 114;
	{8'd255,8'd75} : s = 113;
	{8'd255,8'd76} : s = 242;
	{8'd255,8'd77} : s = 108;
	{8'd255,8'd78} : s = 241;
	{8'd255,8'd79} : s = 236;
	{8'd255,8'd80} : s = 399;
	{8'd255,8'd81} : s = 26;
	{8'd255,8'd82} : s = 106;
	{8'd255,8'd83} : s = 105;
	{8'd255,8'd84} : s = 234;
	{8'd255,8'd85} : s = 102;
	{8'd255,8'd86} : s = 233;
	{8'd255,8'd87} : s = 230;
	{8'd255,8'd88} : s = 380;
	{8'd255,8'd89} : s = 101;
	{8'd255,8'd90} : s = 229;
	{8'd255,8'd91} : s = 227;
	{8'd255,8'd92} : s = 378;
	{8'd255,8'd93} : s = 220;
	{8'd255,8'd94} : s = 377;
	{8'd255,8'd95} : s = 374;
	{8'd255,8'd96} : s = 487;
	{8'd255,8'd97} : s = 25;
	{8'd255,8'd98} : s = 99;
	{8'd255,8'd99} : s = 92;
	{8'd255,8'd100} : s = 218;
	{8'd255,8'd101} : s = 90;
	{8'd255,8'd102} : s = 217;
	{8'd255,8'd103} : s = 214;
	{8'd255,8'd104} : s = 373;
	{8'd255,8'd105} : s = 89;
	{8'd255,8'd106} : s = 213;
	{8'd255,8'd107} : s = 211;
	{8'd255,8'd108} : s = 371;
	{8'd255,8'd109} : s = 206;
	{8'd255,8'd110} : s = 366;
	{8'd255,8'd111} : s = 365;
	{8'd255,8'd112} : s = 478;
	{8'd255,8'd113} : s = 86;
	{8'd255,8'd114} : s = 205;
	{8'd255,8'd115} : s = 203;
	{8'd255,8'd116} : s = 363;
	{8'd255,8'd117} : s = 199;
	{8'd255,8'd118} : s = 359;
	{8'd255,8'd119} : s = 350;
	{8'd255,8'd120} : s = 477;
	{8'd255,8'd121} : s = 188;
	{8'd255,8'd122} : s = 349;
	{8'd255,8'd123} : s = 347;
	{8'd255,8'd124} : s = 475;
	{8'd255,8'd125} : s = 343;
	{8'd255,8'd126} : s = 471;
	{8'd255,8'd127} : s = 463;
	{8'd255,8'd128} : s = 509;
	{8'd255,8'd129} : s = 3;
	{8'd255,8'd130} : s = 22;
	{8'd255,8'd131} : s = 21;
	{8'd255,8'd132} : s = 85;
	{8'd255,8'd133} : s = 19;
	{8'd255,8'd134} : s = 83;
	{8'd255,8'd135} : s = 78;
	{8'd255,8'd136} : s = 186;
	{8'd255,8'd137} : s = 14;
	{8'd255,8'd138} : s = 77;
	{8'd255,8'd139} : s = 75;
	{8'd255,8'd140} : s = 185;
	{8'd255,8'd141} : s = 71;
	{8'd255,8'd142} : s = 182;
	{8'd255,8'd143} : s = 181;
	{8'd255,8'd144} : s = 335;
	{8'd255,8'd145} : s = 13;
	{8'd255,8'd146} : s = 60;
	{8'd255,8'd147} : s = 58;
	{8'd255,8'd148} : s = 179;
	{8'd255,8'd149} : s = 57;
	{8'd255,8'd150} : s = 174;
	{8'd255,8'd151} : s = 173;
	{8'd255,8'd152} : s = 318;
	{8'd255,8'd153} : s = 54;
	{8'd255,8'd154} : s = 171;
	{8'd255,8'd155} : s = 167;
	{8'd255,8'd156} : s = 317;
	{8'd255,8'd157} : s = 158;
	{8'd255,8'd158} : s = 315;
	{8'd255,8'd159} : s = 311;
	{8'd255,8'd160} : s = 446;
	{8'd255,8'd161} : s = 11;
	{8'd255,8'd162} : s = 53;
	{8'd255,8'd163} : s = 51;
	{8'd255,8'd164} : s = 157;
	{8'd255,8'd165} : s = 46;
	{8'd255,8'd166} : s = 155;
	{8'd255,8'd167} : s = 151;
	{8'd255,8'd168} : s = 303;
	{8'd255,8'd169} : s = 45;
	{8'd255,8'd170} : s = 143;
	{8'd255,8'd171} : s = 124;
	{8'd255,8'd172} : s = 287;
	{8'd255,8'd173} : s = 122;
	{8'd255,8'd174} : s = 252;
	{8'd255,8'd175} : s = 250;
	{8'd255,8'd176} : s = 445;
	{8'd255,8'd177} : s = 43;
	{8'd255,8'd178} : s = 121;
	{8'd255,8'd179} : s = 118;
	{8'd255,8'd180} : s = 249;
	{8'd255,8'd181} : s = 117;
	{8'd255,8'd182} : s = 246;
	{8'd255,8'd183} : s = 245;
	{8'd255,8'd184} : s = 443;
	{8'd255,8'd185} : s = 115;
	{8'd255,8'd186} : s = 243;
	{8'd255,8'd187} : s = 238;
	{8'd255,8'd188} : s = 439;
	{8'd255,8'd189} : s = 237;
	{8'd255,8'd190} : s = 431;
	{8'd255,8'd191} : s = 415;
	{8'd255,8'd192} : s = 507;
	{8'd255,8'd193} : s = 7;
	{8'd255,8'd194} : s = 39;
	{8'd255,8'd195} : s = 30;
	{8'd255,8'd196} : s = 110;
	{8'd255,8'd197} : s = 29;
	{8'd255,8'd198} : s = 109;
	{8'd255,8'd199} : s = 107;
	{8'd255,8'd200} : s = 235;
	{8'd255,8'd201} : s = 27;
	{8'd255,8'd202} : s = 103;
	{8'd255,8'd203} : s = 94;
	{8'd255,8'd204} : s = 231;
	{8'd255,8'd205} : s = 93;
	{8'd255,8'd206} : s = 222;
	{8'd255,8'd207} : s = 221;
	{8'd255,8'd208} : s = 382;
	{8'd255,8'd209} : s = 23;
	{8'd255,8'd210} : s = 91;
	{8'd255,8'd211} : s = 87;
	{8'd255,8'd212} : s = 219;
	{8'd255,8'd213} : s = 79;
	{8'd255,8'd214} : s = 215;
	{8'd255,8'd215} : s = 207;
	{8'd255,8'd216} : s = 381;
	{8'd255,8'd217} : s = 62;
	{8'd255,8'd218} : s = 190;
	{8'd255,8'd219} : s = 189;
	{8'd255,8'd220} : s = 379;
	{8'd255,8'd221} : s = 187;
	{8'd255,8'd222} : s = 375;
	{8'd255,8'd223} : s = 367;
	{8'd255,8'd224} : s = 503;
	{8'd255,8'd225} : s = 15;
	{8'd255,8'd226} : s = 61;
	{8'd255,8'd227} : s = 59;
	{8'd255,8'd228} : s = 183;
	{8'd255,8'd229} : s = 55;
	{8'd255,8'd230} : s = 175;
	{8'd255,8'd231} : s = 159;
	{8'd255,8'd232} : s = 351;
	{8'd255,8'd233} : s = 47;
	{8'd255,8'd234} : s = 126;
	{8'd255,8'd235} : s = 125;
	{8'd255,8'd236} : s = 319;
	{8'd255,8'd237} : s = 123;
	{8'd255,8'd238} : s = 254;
	{8'd255,8'd239} : s = 253;
	{8'd255,8'd240} : s = 479;
	{8'd255,8'd241} : s = 31;
	{8'd255,8'd242} : s = 119;
	{8'd255,8'd243} : s = 111;
	{8'd255,8'd244} : s = 251;
	{8'd255,8'd245} : s = 95;
	{8'd255,8'd246} : s = 247;
	{8'd255,8'd247} : s = 239;
	{8'd255,8'd248} : s = 495;
	{8'd255,8'd249} : s = 63;
	{8'd255,8'd250} : s = 223;
	{8'd255,8'd251} : s = 191;
	{8'd255,8'd252} : s = 447;
	{8'd255,8'd253} : s = 127;
	{8'd255,8'd254} : s = 383;
	{8'd255,8'd255} : s = 255;
    endcase
end
endmodule
