module adder8nit_mapped(a__0, a__1, a__2, a__3, a__4, a__5, a__6, a__7,b__0, b__1, b__2, b__3, b__4, b__5, b__6, b__7s__0, s__1, s__2, s__3, s__4, s__5, s__6, s__7):
  input a__0, a__1, a__2, a__3, a__4, a__5, a__6, a__7;
  input b__0, b__1, b__2, b__3, b__4, b__5, b__6, b__7;
  output s__0, s__1, s__2, s__3, s__4, s__5, s__6, s__7;
  input cin;
  output cout;
  wire   N0, N1, N2, N3, N4, N5, N6;
  assign s__0 = p__0 ^ cin;
  assign s__1 = p__1 ^ c__1;
  assign s__2 = p__2 ^ c__2;
  assign s__3 = p__3 ^ c__3;
  assign s__4 = p__4 ^ c__4;
  assign s__5 = p__5 ^ c__5;
  assign s__6 = p__6 ^ c__6;
  assign s__7 = p__7 ^ c__7;
  assign N6 = p__6 & c__6;
  assign c__7 = g__6 | N6;
  assign N5 = p__5 & c__5;
  assign c__6 = g__5 | N5;
  assign N4 = p__4 & c__4;
  assign c__5 = g__4 | N4;
  assign N3 = p__3 & c__3;
  assign c__4 = g__3 | N3;
  assign N2 = p__2 & c__2;
  assign c__3 = g__2 | N2;
  assign N1 = p__1 & c__1;
  assign c__2 = g__1 | N1;
  assign N0 = p__0 & cin;
  assign c__1 = g__0 | N0;
  assign p__0 = a__0 ^ b__0;
  assign p__1 = a__1 ^ b__1;
  assign p__2 = a__2 ^ b__2;
  assign p__3 = a__3 ^ b__3;
  assign p__4 = a__4 ^ b__4;
  assign p__5 = a__5 ^ b__5;
  assign p__6 = a__6 ^ b__6;
  assign p__7 = a__7 ^ b__7;
  assign g__0 = a__0 & b__0;
  assign g__1 = a__1 & b__1;
  assign g__2 = a__2 & b__2;
  assign g__3 = a__3 & b__3;
  assign g__4 = a__4 & b__4;
  assign g__5 = a__5 & b__5;
  assign g__6 = a__6 & b__6;
