
module gen_nonlinear_part ( a, b, c, n );
  input [6:0] a;
  input [6:0] b;
  output [500:0] n;
  input c;
  wire   n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654;

  INVD0 U716 ( .I(b[6]), .ZN(n423) );
  INVD0 U717 ( .I(b[6]), .ZN(n424) );
  INVD0 U718 ( .I(b[6]), .ZN(n425) );
  INVD0 U719 ( .I(b[6]), .ZN(n426) );
  INVD0 U720 ( .I(b[6]), .ZN(n427) );
  INVD0 U721 ( .I(b[6]), .ZN(n428) );
  INVD0 U722 ( .I(b[6]), .ZN(n429) );
  INVD0 U723 ( .I(b[6]), .ZN(n430) );
  INVD0 U724 ( .I(b[6]), .ZN(n431) );
  INVD0 U725 ( .I(b[6]), .ZN(n432) );
  INVD0 U726 ( .I(a[6]), .ZN(n433) );
  INVD0 U727 ( .I(a[6]), .ZN(n434) );
  INVD0 U728 ( .I(a[6]), .ZN(n435) );
  INVD0 U729 ( .I(a[6]), .ZN(n436) );
  INVD0 U730 ( .I(a[6]), .ZN(n437) );
  INVD0 U731 ( .I(a[6]), .ZN(n438) );
  INVD0 U732 ( .I(a[6]), .ZN(n439) );
  INVD0 U733 ( .I(a[6]), .ZN(n440) );
  INVD0 U734 ( .I(a[6]), .ZN(n441) );
  INVD0 U735 ( .I(a[6]), .ZN(n442) );
  NR2D0 U736 ( .A1(n443), .A2(n432), .ZN(n[500]) );
  NR2D0 U737 ( .A1(n432), .A2(n444), .ZN(n[499]) );
  NR2D0 U738 ( .A1(n432), .A2(n445), .ZN(n[498]) );
  NR2D0 U739 ( .A1(n432), .A2(n446), .ZN(n[497]) );
  NR2D0 U740 ( .A1(n432), .A2(n447), .ZN(n[496]) );
  NR2D0 U741 ( .A1(n432), .A2(n448), .ZN(n[495]) );
  NR2D0 U742 ( .A1(n432), .A2(n449), .ZN(n[494]) );
  NR2D0 U743 ( .A1(n432), .A2(n450), .ZN(n[493]) );
  NR2D0 U744 ( .A1(n432), .A2(n451), .ZN(n[492]) );
  NR2D0 U745 ( .A1(n432), .A2(n452), .ZN(n[491]) );
  NR2D0 U746 ( .A1(n432), .A2(n453), .ZN(n[490]) );
  NR2D0 U747 ( .A1(n431), .A2(n454), .ZN(n[489]) );
  NR2D0 U748 ( .A1(n431), .A2(n455), .ZN(n[488]) );
  NR2D0 U749 ( .A1(n431), .A2(n456), .ZN(n[487]) );
  NR2D0 U750 ( .A1(n431), .A2(n457), .ZN(n[486]) );
  NR2D0 U751 ( .A1(n431), .A2(n458), .ZN(n[485]) );
  NR2D0 U752 ( .A1(n431), .A2(n459), .ZN(n[484]) );
  NR2D0 U753 ( .A1(n431), .A2(n460), .ZN(n[483]) );
  NR2D0 U754 ( .A1(n431), .A2(n461), .ZN(n[482]) );
  NR2D0 U755 ( .A1(n431), .A2(n462), .ZN(n[481]) );
  NR2D0 U756 ( .A1(n431), .A2(n463), .ZN(n[480]) );
  NR2D0 U757 ( .A1(n431), .A2(n464), .ZN(n[479]) );
  NR2D0 U758 ( .A1(n431), .A2(n465), .ZN(n[478]) );
  NR2D0 U759 ( .A1(n431), .A2(n466), .ZN(n[477]) );
  NR2D0 U760 ( .A1(n430), .A2(n467), .ZN(n[476]) );
  NR2D0 U761 ( .A1(n430), .A2(n468), .ZN(n[475]) );
  NR2D0 U762 ( .A1(n430), .A2(n469), .ZN(n[474]) );
  NR2D0 U763 ( .A1(n430), .A2(n470), .ZN(n[473]) );
  NR2D0 U764 ( .A1(n430), .A2(n471), .ZN(n[472]) );
  NR2D0 U765 ( .A1(n430), .A2(n472), .ZN(n[471]) );
  NR2D0 U766 ( .A1(n430), .A2(n473), .ZN(n[470]) );
  NR2D0 U767 ( .A1(n430), .A2(n474), .ZN(n[469]) );
  NR2D0 U768 ( .A1(n430), .A2(n475), .ZN(n[468]) );
  NR2D0 U769 ( .A1(n430), .A2(n476), .ZN(n[467]) );
  NR2D0 U770 ( .A1(n430), .A2(n477), .ZN(n[466]) );
  NR2D0 U771 ( .A1(n430), .A2(n478), .ZN(n[465]) );
  NR2D0 U772 ( .A1(n430), .A2(n479), .ZN(n[464]) );
  NR2D0 U773 ( .A1(n429), .A2(n480), .ZN(n[463]) );
  NR2D0 U774 ( .A1(n429), .A2(n481), .ZN(n[462]) );
  NR2D0 U775 ( .A1(n429), .A2(n482), .ZN(n[461]) );
  NR2D0 U776 ( .A1(n429), .A2(n483), .ZN(n[460]) );
  NR2D0 U777 ( .A1(n429), .A2(n484), .ZN(n[459]) );
  NR2D0 U778 ( .A1(n429), .A2(n485), .ZN(n[458]) );
  NR2D0 U779 ( .A1(n429), .A2(n486), .ZN(n[457]) );
  NR2D0 U780 ( .A1(n429), .A2(n487), .ZN(n[456]) );
  NR2D0 U781 ( .A1(n429), .A2(n488), .ZN(n[455]) );
  NR2D0 U782 ( .A1(n429), .A2(n489), .ZN(n[454]) );
  NR2D0 U783 ( .A1(n429), .A2(n490), .ZN(n[453]) );
  NR2D0 U784 ( .A1(n429), .A2(n491), .ZN(n[452]) );
  NR2D0 U785 ( .A1(n429), .A2(n492), .ZN(n[451]) );
  NR2D0 U786 ( .A1(n428), .A2(n493), .ZN(n[450]) );
  NR2D0 U787 ( .A1(n428), .A2(n494), .ZN(n[449]) );
  NR2D0 U788 ( .A1(n428), .A2(n495), .ZN(n[448]) );
  NR2D0 U789 ( .A1(n428), .A2(n496), .ZN(n[447]) );
  NR2D0 U790 ( .A1(n428), .A2(n497), .ZN(n[446]) );
  NR2D0 U791 ( .A1(n428), .A2(n498), .ZN(n[445]) );
  NR2D0 U792 ( .A1(n428), .A2(n499), .ZN(n[444]) );
  NR2D0 U793 ( .A1(n428), .A2(n500), .ZN(n[443]) );
  NR2D0 U794 ( .A1(n428), .A2(n501), .ZN(n[442]) );
  NR2D0 U795 ( .A1(n428), .A2(n502), .ZN(n[441]) );
  NR2D0 U796 ( .A1(n428), .A2(n503), .ZN(n[440]) );
  NR2D0 U797 ( .A1(n428), .A2(n504), .ZN(n[439]) );
  NR2D0 U798 ( .A1(n428), .A2(n505), .ZN(n[438]) );
  NR2D0 U799 ( .A1(n427), .A2(n506), .ZN(n[437]) );
  NR2D0 U800 ( .A1(n427), .A2(n507), .ZN(n[436]) );
  NR2D0 U801 ( .A1(n427), .A2(n508), .ZN(n[435]) );
  NR2D0 U802 ( .A1(n427), .A2(n509), .ZN(n[434]) );
  NR2D0 U803 ( .A1(n427), .A2(n510), .ZN(n[433]) );
  NR2D0 U804 ( .A1(n427), .A2(n511), .ZN(n[432]) );
  NR2D0 U805 ( .A1(n427), .A2(n512), .ZN(n[431]) );
  NR2D0 U806 ( .A1(n427), .A2(n513), .ZN(n[430]) );
  NR2D0 U807 ( .A1(n427), .A2(n514), .ZN(n[429]) );
  NR2D0 U808 ( .A1(n427), .A2(n515), .ZN(n[428]) );
  NR2D0 U809 ( .A1(n427), .A2(n516), .ZN(n[427]) );
  NR2D0 U810 ( .A1(n427), .A2(n517), .ZN(n[426]) );
  NR2D0 U811 ( .A1(n427), .A2(n518), .ZN(n[425]) );
  NR2D0 U812 ( .A1(n426), .A2(n519), .ZN(n[424]) );
  NR2D0 U813 ( .A1(n426), .A2(n520), .ZN(n[423]) );
  NR2D0 U814 ( .A1(n426), .A2(n521), .ZN(n[422]) );
  NR2D0 U815 ( .A1(n426), .A2(n522), .ZN(n[421]) );
  NR2D0 U816 ( .A1(n426), .A2(n523), .ZN(n[420]) );
  NR2D0 U817 ( .A1(n426), .A2(n524), .ZN(n[419]) );
  NR2D0 U818 ( .A1(n426), .A2(n525), .ZN(n[418]) );
  NR2D0 U819 ( .A1(n426), .A2(n526), .ZN(n[417]) );
  NR2D0 U820 ( .A1(n426), .A2(n527), .ZN(n[416]) );
  NR2D0 U821 ( .A1(n426), .A2(n528), .ZN(n[415]) );
  NR2D0 U822 ( .A1(n426), .A2(n529), .ZN(n[414]) );
  NR2D0 U823 ( .A1(n426), .A2(n530), .ZN(n[413]) );
  NR2D0 U824 ( .A1(n426), .A2(n531), .ZN(n[412]) );
  NR2D0 U825 ( .A1(n425), .A2(n532), .ZN(n[411]) );
  NR2D0 U826 ( .A1(n425), .A2(n533), .ZN(n[410]) );
  NR2D0 U827 ( .A1(n425), .A2(n534), .ZN(n[409]) );
  NR2D0 U828 ( .A1(n425), .A2(n535), .ZN(n[408]) );
  NR2D0 U829 ( .A1(n425), .A2(n536), .ZN(n[407]) );
  NR2D0 U830 ( .A1(n425), .A2(n537), .ZN(n[406]) );
  NR2D0 U831 ( .A1(n425), .A2(n538), .ZN(n[405]) );
  NR2D0 U832 ( .A1(n425), .A2(n539), .ZN(n[404]) );
  NR2D0 U833 ( .A1(n425), .A2(n540), .ZN(n[403]) );
  NR2D0 U834 ( .A1(n425), .A2(n541), .ZN(n[402]) );
  NR2D0 U835 ( .A1(n425), .A2(n542), .ZN(n[401]) );
  NR2D0 U836 ( .A1(n425), .A2(n543), .ZN(n[400]) );
  NR2D0 U837 ( .A1(n425), .A2(n544), .ZN(n[399]) );
  NR2D0 U838 ( .A1(n424), .A2(n545), .ZN(n[398]) );
  NR2D0 U839 ( .A1(n424), .A2(n546), .ZN(n[397]) );
  NR2D0 U840 ( .A1(n424), .A2(n547), .ZN(n[396]) );
  NR2D0 U841 ( .A1(n424), .A2(n548), .ZN(n[395]) );
  NR2D0 U842 ( .A1(n424), .A2(n549), .ZN(n[394]) );
  NR2D0 U843 ( .A1(n424), .A2(n550), .ZN(n[393]) );
  NR2D0 U844 ( .A1(n424), .A2(n551), .ZN(n[392]) );
  NR2D0 U845 ( .A1(n424), .A2(n552), .ZN(n[391]) );
  NR2D0 U846 ( .A1(n424), .A2(n553), .ZN(n[390]) );
  NR2D0 U847 ( .A1(n424), .A2(n554), .ZN(n[389]) );
  NR2D0 U848 ( .A1(n424), .A2(n555), .ZN(n[388]) );
  NR2D0 U849 ( .A1(n424), .A2(n556), .ZN(n[387]) );
  NR2D0 U850 ( .A1(n424), .A2(n557), .ZN(n[386]) );
  NR2D0 U851 ( .A1(n423), .A2(n558), .ZN(n[385]) );
  NR2D0 U852 ( .A1(n423), .A2(n559), .ZN(n[384]) );
  NR2D0 U853 ( .A1(n423), .A2(n560), .ZN(n[383]) );
  NR2D0 U854 ( .A1(n423), .A2(n561), .ZN(n[382]) );
  NR2D0 U855 ( .A1(n423), .A2(n562), .ZN(n[381]) );
  NR2D0 U856 ( .A1(n423), .A2(n563), .ZN(n[380]) );
  NR2D0 U857 ( .A1(n423), .A2(n564), .ZN(n[379]) );
  NR2D0 U858 ( .A1(n423), .A2(n565), .ZN(n[378]) );
  NR2D0 U859 ( .A1(n423), .A2(n566), .ZN(n[377]) );
  NR2D0 U860 ( .A1(n423), .A2(n567), .ZN(n[376]) );
  NR2D0 U861 ( .A1(n423), .A2(n568), .ZN(n[375]) );
  NR2D0 U862 ( .A1(n423), .A2(n569), .ZN(n[374]) );
  NR2D0 U863 ( .A1(n443), .A2(n442), .ZN(n[373]) );
  NR2D0 U864 ( .A1(n444), .A2(n442), .ZN(n[372]) );
  NR2D0 U865 ( .A1(n445), .A2(n442), .ZN(n[371]) );
  NR2D0 U866 ( .A1(n446), .A2(n442), .ZN(n[370]) );
  NR2D0 U867 ( .A1(n447), .A2(n442), .ZN(n[369]) );
  NR2D0 U868 ( .A1(n448), .A2(n442), .ZN(n[368]) );
  NR2D0 U869 ( .A1(n449), .A2(n442), .ZN(n[367]) );
  NR2D0 U870 ( .A1(n450), .A2(n442), .ZN(n[366]) );
  NR2D0 U871 ( .A1(n451), .A2(n442), .ZN(n[365]) );
  NR2D0 U872 ( .A1(n452), .A2(n442), .ZN(n[364]) );
  NR2D0 U873 ( .A1(n453), .A2(n442), .ZN(n[363]) );
  NR2D0 U874 ( .A1(n454), .A2(n441), .ZN(n[362]) );
  NR2D0 U875 ( .A1(n455), .A2(n441), .ZN(n[361]) );
  NR2D0 U876 ( .A1(n456), .A2(n441), .ZN(n[360]) );
  NR2D0 U877 ( .A1(n457), .A2(n441), .ZN(n[359]) );
  NR2D0 U878 ( .A1(n458), .A2(n441), .ZN(n[358]) );
  NR2D0 U879 ( .A1(n459), .A2(n441), .ZN(n[357]) );
  NR2D0 U880 ( .A1(n460), .A2(n441), .ZN(n[356]) );
  NR2D0 U881 ( .A1(n461), .A2(n441), .ZN(n[355]) );
  NR2D0 U882 ( .A1(n462), .A2(n441), .ZN(n[354]) );
  NR2D0 U883 ( .A1(n463), .A2(n441), .ZN(n[353]) );
  NR2D0 U884 ( .A1(n464), .A2(n441), .ZN(n[352]) );
  NR2D0 U885 ( .A1(n465), .A2(n441), .ZN(n[351]) );
  NR2D0 U886 ( .A1(n466), .A2(n441), .ZN(n[350]) );
  NR2D0 U887 ( .A1(n467), .A2(n440), .ZN(n[349]) );
  NR2D0 U888 ( .A1(n468), .A2(n440), .ZN(n[348]) );
  NR2D0 U889 ( .A1(n469), .A2(n440), .ZN(n[347]) );
  NR2D0 U890 ( .A1(n470), .A2(n440), .ZN(n[346]) );
  NR2D0 U891 ( .A1(n471), .A2(n440), .ZN(n[345]) );
  NR2D0 U892 ( .A1(n472), .A2(n440), .ZN(n[344]) );
  NR2D0 U893 ( .A1(n473), .A2(n440), .ZN(n[343]) );
  NR2D0 U894 ( .A1(n474), .A2(n440), .ZN(n[342]) );
  NR2D0 U895 ( .A1(n475), .A2(n440), .ZN(n[341]) );
  NR2D0 U896 ( .A1(n476), .A2(n440), .ZN(n[340]) );
  NR2D0 U897 ( .A1(n477), .A2(n440), .ZN(n[339]) );
  NR2D0 U898 ( .A1(n478), .A2(n440), .ZN(n[338]) );
  NR2D0 U899 ( .A1(n479), .A2(n440), .ZN(n[337]) );
  NR2D0 U900 ( .A1(n480), .A2(n439), .ZN(n[336]) );
  NR2D0 U901 ( .A1(n481), .A2(n439), .ZN(n[335]) );
  NR2D0 U902 ( .A1(n482), .A2(n439), .ZN(n[334]) );
  NR2D0 U903 ( .A1(n483), .A2(n439), .ZN(n[333]) );
  NR2D0 U904 ( .A1(n484), .A2(n439), .ZN(n[332]) );
  NR2D0 U905 ( .A1(n485), .A2(n439), .ZN(n[331]) );
  NR2D0 U906 ( .A1(n486), .A2(n439), .ZN(n[330]) );
  NR2D0 U907 ( .A1(n487), .A2(n439), .ZN(n[329]) );
  NR2D0 U908 ( .A1(n488), .A2(n439), .ZN(n[328]) );
  NR2D0 U909 ( .A1(n489), .A2(n439), .ZN(n[327]) );
  NR2D0 U910 ( .A1(n490), .A2(n439), .ZN(n[326]) );
  NR2D0 U911 ( .A1(n491), .A2(n439), .ZN(n[325]) );
  NR2D0 U912 ( .A1(n492), .A2(n439), .ZN(n[324]) );
  NR2D0 U913 ( .A1(n493), .A2(n438), .ZN(n[323]) );
  NR2D0 U914 ( .A1(n494), .A2(n438), .ZN(n[322]) );
  NR2D0 U915 ( .A1(n495), .A2(n438), .ZN(n[321]) );
  NR2D0 U916 ( .A1(n496), .A2(n438), .ZN(n[320]) );
  NR2D0 U917 ( .A1(n497), .A2(n438), .ZN(n[319]) );
  NR2D0 U918 ( .A1(n498), .A2(n438), .ZN(n[318]) );
  NR2D0 U919 ( .A1(n499), .A2(n438), .ZN(n[317]) );
  NR2D0 U920 ( .A1(n500), .A2(n438), .ZN(n[316]) );
  NR2D0 U921 ( .A1(n501), .A2(n438), .ZN(n[315]) );
  NR2D0 U922 ( .A1(n502), .A2(n438), .ZN(n[314]) );
  NR2D0 U923 ( .A1(n503), .A2(n438), .ZN(n[313]) );
  NR2D0 U924 ( .A1(n504), .A2(n438), .ZN(n[312]) );
  NR2D0 U925 ( .A1(n505), .A2(n438), .ZN(n[311]) );
  NR2D0 U926 ( .A1(n506), .A2(n437), .ZN(n[310]) );
  NR2D0 U927 ( .A1(n507), .A2(n437), .ZN(n[309]) );
  NR2D0 U928 ( .A1(n508), .A2(n437), .ZN(n[308]) );
  NR2D0 U929 ( .A1(n509), .A2(n437), .ZN(n[307]) );
  NR2D0 U930 ( .A1(n510), .A2(n437), .ZN(n[306]) );
  NR2D0 U931 ( .A1(n511), .A2(n437), .ZN(n[305]) );
  NR2D0 U932 ( .A1(n512), .A2(n437), .ZN(n[304]) );
  NR2D0 U933 ( .A1(n513), .A2(n437), .ZN(n[303]) );
  NR2D0 U934 ( .A1(n514), .A2(n437), .ZN(n[302]) );
  NR2D0 U935 ( .A1(n515), .A2(n437), .ZN(n[301]) );
  NR2D0 U936 ( .A1(n516), .A2(n437), .ZN(n[300]) );
  INVD0 U937 ( .I(n570), .ZN(n[2]) );
  NR2D0 U938 ( .A1(n517), .A2(n437), .ZN(n[299]) );
  NR2D0 U939 ( .A1(n518), .A2(n437), .ZN(n[298]) );
  NR2D0 U940 ( .A1(n519), .A2(n436), .ZN(n[297]) );
  NR2D0 U941 ( .A1(n520), .A2(n436), .ZN(n[296]) );
  NR2D0 U942 ( .A1(n521), .A2(n436), .ZN(n[295]) );
  NR2D0 U943 ( .A1(n522), .A2(n436), .ZN(n[294]) );
  NR2D0 U944 ( .A1(n523), .A2(n436), .ZN(n[293]) );
  NR2D0 U945 ( .A1(n524), .A2(n436), .ZN(n[292]) );
  NR2D0 U946 ( .A1(n525), .A2(n436), .ZN(n[291]) );
  NR2D0 U947 ( .A1(n526), .A2(n436), .ZN(n[290]) );
  NR2D0 U948 ( .A1(n527), .A2(n436), .ZN(n[289]) );
  NR2D0 U949 ( .A1(n528), .A2(n436), .ZN(n[288]) );
  NR2D0 U950 ( .A1(n529), .A2(n436), .ZN(n[287]) );
  NR2D0 U951 ( .A1(n530), .A2(n436), .ZN(n[286]) );
  NR2D0 U952 ( .A1(n531), .A2(n436), .ZN(n[285]) );
  NR2D0 U953 ( .A1(n532), .A2(n435), .ZN(n[284]) );
  NR2D0 U954 ( .A1(n533), .A2(n435), .ZN(n[283]) );
  NR2D0 U955 ( .A1(n534), .A2(n435), .ZN(n[282]) );
  NR2D0 U956 ( .A1(n535), .A2(n435), .ZN(n[281]) );
  NR2D0 U957 ( .A1(n536), .A2(n435), .ZN(n[280]) );
  NR2D0 U958 ( .A1(n537), .A2(n435), .ZN(n[279]) );
  NR2D0 U959 ( .A1(n538), .A2(n435), .ZN(n[278]) );
  NR2D0 U960 ( .A1(n539), .A2(n435), .ZN(n[277]) );
  NR2D0 U961 ( .A1(n540), .A2(n435), .ZN(n[276]) );
  NR2D0 U962 ( .A1(n541), .A2(n435), .ZN(n[275]) );
  NR2D0 U963 ( .A1(n542), .A2(n435), .ZN(n[274]) );
  NR2D0 U964 ( .A1(n543), .A2(n435), .ZN(n[273]) );
  NR2D0 U965 ( .A1(n544), .A2(n435), .ZN(n[272]) );
  NR2D0 U966 ( .A1(n545), .A2(n434), .ZN(n[271]) );
  NR2D0 U967 ( .A1(n546), .A2(n434), .ZN(n[270]) );
  NR2D0 U968 ( .A1(n547), .A2(n434), .ZN(n[269]) );
  NR2D0 U969 ( .A1(n548), .A2(n434), .ZN(n[268]) );
  NR2D0 U970 ( .A1(n549), .A2(n434), .ZN(n[267]) );
  NR2D0 U971 ( .A1(n550), .A2(n434), .ZN(n[266]) );
  NR2D0 U972 ( .A1(n551), .A2(n434), .ZN(n[265]) );
  NR2D0 U973 ( .A1(n552), .A2(n434), .ZN(n[264]) );
  NR2D0 U974 ( .A1(n553), .A2(n434), .ZN(n[263]) );
  NR2D0 U975 ( .A1(n554), .A2(n434), .ZN(n[262]) );
  NR2D0 U976 ( .A1(n555), .A2(n434), .ZN(n[261]) );
  NR2D0 U977 ( .A1(n556), .A2(n434), .ZN(n[260]) );
  NR2D0 U978 ( .A1(n557), .A2(n434), .ZN(n[259]) );
  NR2D0 U979 ( .A1(n558), .A2(n433), .ZN(n[258]) );
  NR2D0 U980 ( .A1(n559), .A2(n433), .ZN(n[257]) );
  NR2D0 U981 ( .A1(n560), .A2(n433), .ZN(n[256]) );
  NR2D0 U982 ( .A1(n561), .A2(n433), .ZN(n[255]) );
  NR2D0 U983 ( .A1(n562), .A2(n433), .ZN(n[254]) );
  NR2D0 U984 ( .A1(n563), .A2(n433), .ZN(n[253]) );
  NR2D0 U985 ( .A1(n564), .A2(n433), .ZN(n[252]) );
  NR2D0 U986 ( .A1(n565), .A2(n433), .ZN(n[251]) );
  NR2D0 U987 ( .A1(n566), .A2(n433), .ZN(n[250]) );
  INVD0 U988 ( .I(n571), .ZN(n[24]) );
  NR2D0 U989 ( .A1(n567), .A2(n433), .ZN(n[249]) );
  NR2D0 U990 ( .A1(n568), .A2(n433), .ZN(n[248]) );
  NR2D0 U991 ( .A1(n569), .A2(n433), .ZN(n[247]) );
  NR2D0 U992 ( .A1(n423), .A2(n433), .ZN(n[246]) );
  INVD0 U993 ( .I(n443), .ZN(n[245]) );
  ND2D0 U994 ( .A1(b[5]), .A2(n[118]), .ZN(n443) );
  INVD0 U995 ( .I(n444), .ZN(n[244]) );
  ND2D0 U996 ( .A1(n[117]), .A2(b[5]), .ZN(n444) );
  INVD0 U997 ( .I(n445), .ZN(n[243]) );
  ND2D0 U998 ( .A1(n[116]), .A2(b[5]), .ZN(n445) );
  INVD0 U999 ( .I(n446), .ZN(n[242]) );
  ND2D0 U1000 ( .A1(n[115]), .A2(b[5]), .ZN(n446) );
  INVD0 U1001 ( .I(n447), .ZN(n[241]) );
  ND2D0 U1002 ( .A1(n[114]), .A2(b[5]), .ZN(n447) );
  INVD0 U1003 ( .I(n448), .ZN(n[240]) );
  ND2D0 U1004 ( .A1(n[113]), .A2(b[5]), .ZN(n448) );
  INVD0 U1005 ( .I(n572), .ZN(n[23]) );
  INVD0 U1006 ( .I(n449), .ZN(n[239]) );
  ND2D0 U1007 ( .A1(n[112]), .A2(b[5]), .ZN(n449) );
  INVD0 U1008 ( .I(n450), .ZN(n[238]) );
  ND2D0 U1009 ( .A1(n[111]), .A2(b[5]), .ZN(n450) );
  INVD0 U1010 ( .I(n451), .ZN(n[237]) );
  ND2D0 U1011 ( .A1(n[110]), .A2(b[5]), .ZN(n451) );
  INVD0 U1012 ( .I(n452), .ZN(n[236]) );
  ND2D0 U1013 ( .A1(n[109]), .A2(b[5]), .ZN(n452) );
  INVD0 U1014 ( .I(n453), .ZN(n[235]) );
  ND2D0 U1015 ( .A1(n[108]), .A2(b[5]), .ZN(n453) );
  INVD0 U1016 ( .I(n454), .ZN(n[234]) );
  ND2D0 U1017 ( .A1(n[107]), .A2(b[5]), .ZN(n454) );
  INVD0 U1018 ( .I(n455), .ZN(n[233]) );
  ND2D0 U1019 ( .A1(n[106]), .A2(b[5]), .ZN(n455) );
  INVD0 U1020 ( .I(n456), .ZN(n[232]) );
  ND2D0 U1021 ( .A1(n[105]), .A2(b[5]), .ZN(n456) );
  INVD0 U1022 ( .I(n457), .ZN(n[231]) );
  ND2D0 U1023 ( .A1(n[104]), .A2(b[5]), .ZN(n457) );
  INVD0 U1024 ( .I(n458), .ZN(n[230]) );
  ND2D0 U1025 ( .A1(n[103]), .A2(b[5]), .ZN(n458) );
  INVD0 U1026 ( .I(n573), .ZN(n[22]) );
  INVD0 U1027 ( .I(n459), .ZN(n[229]) );
  ND2D0 U1028 ( .A1(n[102]), .A2(b[5]), .ZN(n459) );
  INVD0 U1029 ( .I(n460), .ZN(n[228]) );
  ND2D0 U1030 ( .A1(n[101]), .A2(b[5]), .ZN(n460) );
  INVD0 U1031 ( .I(n461), .ZN(n[227]) );
  ND2D0 U1032 ( .A1(n[100]), .A2(b[5]), .ZN(n461) );
  INVD0 U1033 ( .I(n462), .ZN(n[226]) );
  ND2D0 U1034 ( .A1(n[99]), .A2(b[5]), .ZN(n462) );
  INVD0 U1035 ( .I(n463), .ZN(n[225]) );
  ND2D0 U1036 ( .A1(n[98]), .A2(b[5]), .ZN(n463) );
  INVD0 U1037 ( .I(n464), .ZN(n[224]) );
  ND2D0 U1038 ( .A1(n[97]), .A2(b[5]), .ZN(n464) );
  INVD0 U1039 ( .I(n465), .ZN(n[223]) );
  ND2D0 U1040 ( .A1(n[96]), .A2(b[5]), .ZN(n465) );
  INVD0 U1041 ( .I(n466), .ZN(n[222]) );
  ND2D0 U1042 ( .A1(n[95]), .A2(b[5]), .ZN(n466) );
  INVD0 U1043 ( .I(n467), .ZN(n[221]) );
  ND2D0 U1044 ( .A1(n[94]), .A2(b[5]), .ZN(n467) );
  INVD0 U1045 ( .I(n468), .ZN(n[220]) );
  ND2D0 U1046 ( .A1(n[93]), .A2(b[5]), .ZN(n468) );
  INVD0 U1047 ( .I(n574), .ZN(n[21]) );
  INVD0 U1048 ( .I(n469), .ZN(n[219]) );
  ND2D0 U1049 ( .A1(n[92]), .A2(b[5]), .ZN(n469) );
  INVD0 U1050 ( .I(n470), .ZN(n[218]) );
  ND2D0 U1051 ( .A1(n[91]), .A2(b[5]), .ZN(n470) );
  INVD0 U1052 ( .I(n471), .ZN(n[217]) );
  ND2D0 U1053 ( .A1(n[90]), .A2(b[5]), .ZN(n471) );
  INVD0 U1054 ( .I(n472), .ZN(n[216]) );
  ND2D0 U1055 ( .A1(n[89]), .A2(b[5]), .ZN(n472) );
  INVD0 U1056 ( .I(n473), .ZN(n[215]) );
  ND2D0 U1057 ( .A1(n[88]), .A2(b[5]), .ZN(n473) );
  INVD0 U1058 ( .I(n474), .ZN(n[214]) );
  ND2D0 U1059 ( .A1(n[87]), .A2(b[5]), .ZN(n474) );
  INVD0 U1060 ( .I(n475), .ZN(n[213]) );
  ND2D0 U1061 ( .A1(n[86]), .A2(b[5]), .ZN(n475) );
  INVD0 U1062 ( .I(n476), .ZN(n[212]) );
  ND2D0 U1063 ( .A1(n[85]), .A2(b[5]), .ZN(n476) );
  INVD0 U1064 ( .I(n477), .ZN(n[211]) );
  ND2D0 U1065 ( .A1(n[84]), .A2(b[5]), .ZN(n477) );
  INVD0 U1066 ( .I(n478), .ZN(n[210]) );
  ND2D0 U1067 ( .A1(n[83]), .A2(b[5]), .ZN(n478) );
  INVD0 U1068 ( .I(n575), .ZN(n[20]) );
  INVD0 U1069 ( .I(n479), .ZN(n[209]) );
  ND2D0 U1070 ( .A1(n[82]), .A2(b[5]), .ZN(n479) );
  INVD0 U1071 ( .I(n480), .ZN(n[208]) );
  ND2D0 U1072 ( .A1(n[81]), .A2(b[5]), .ZN(n480) );
  INVD0 U1073 ( .I(n481), .ZN(n[207]) );
  ND2D0 U1074 ( .A1(n[80]), .A2(b[5]), .ZN(n481) );
  INVD0 U1075 ( .I(n482), .ZN(n[206]) );
  ND2D0 U1076 ( .A1(n[79]), .A2(b[5]), .ZN(n482) );
  INVD0 U1077 ( .I(n483), .ZN(n[205]) );
  ND2D0 U1078 ( .A1(n[78]), .A2(b[5]), .ZN(n483) );
  INVD0 U1079 ( .I(n484), .ZN(n[204]) );
  ND2D0 U1080 ( .A1(n[77]), .A2(b[5]), .ZN(n484) );
  INVD0 U1081 ( .I(n485), .ZN(n[203]) );
  ND2D0 U1082 ( .A1(n[76]), .A2(b[5]), .ZN(n485) );
  INVD0 U1083 ( .I(n486), .ZN(n[202]) );
  ND2D0 U1084 ( .A1(n[75]), .A2(b[5]), .ZN(n486) );
  INVD0 U1085 ( .I(n487), .ZN(n[201]) );
  ND2D0 U1086 ( .A1(n[74]), .A2(b[5]), .ZN(n487) );
  INVD0 U1087 ( .I(n488), .ZN(n[200]) );
  ND2D0 U1088 ( .A1(n[73]), .A2(b[5]), .ZN(n488) );
  INVD0 U1089 ( .I(n576), .ZN(n[1]) );
  INVD0 U1090 ( .I(n577), .ZN(n[19]) );
  INVD0 U1091 ( .I(n489), .ZN(n[199]) );
  ND2D0 U1092 ( .A1(n[72]), .A2(b[5]), .ZN(n489) );
  INVD0 U1093 ( .I(n490), .ZN(n[198]) );
  ND2D0 U1094 ( .A1(n[71]), .A2(b[5]), .ZN(n490) );
  INVD0 U1095 ( .I(n491), .ZN(n[197]) );
  ND2D0 U1096 ( .A1(n[70]), .A2(b[5]), .ZN(n491) );
  INVD0 U1097 ( .I(n492), .ZN(n[196]) );
  ND2D0 U1098 ( .A1(n[69]), .A2(b[5]), .ZN(n492) );
  INVD0 U1099 ( .I(n493), .ZN(n[195]) );
  ND2D0 U1100 ( .A1(n[68]), .A2(b[5]), .ZN(n493) );
  INVD0 U1101 ( .I(n494), .ZN(n[194]) );
  ND2D0 U1102 ( .A1(n[67]), .A2(b[5]), .ZN(n494) );
  INVD0 U1103 ( .I(n495), .ZN(n[193]) );
  ND2D0 U1104 ( .A1(n[66]), .A2(b[5]), .ZN(n495) );
  INVD0 U1105 ( .I(n496), .ZN(n[192]) );
  ND2D0 U1106 ( .A1(n[65]), .A2(b[5]), .ZN(n496) );
  INVD0 U1107 ( .I(n497), .ZN(n[191]) );
  ND2D0 U1108 ( .A1(n[64]), .A2(b[5]), .ZN(n497) );
  INVD0 U1109 ( .I(n498), .ZN(n[190]) );
  ND2D0 U1110 ( .A1(n[63]), .A2(b[5]), .ZN(n498) );
  INVD0 U1111 ( .I(n578), .ZN(n[18]) );
  INVD0 U1112 ( .I(n499), .ZN(n[189]) );
  ND2D0 U1113 ( .A1(n[62]), .A2(b[5]), .ZN(n499) );
  INVD0 U1114 ( .I(n500), .ZN(n[188]) );
  ND2D0 U1115 ( .A1(n[61]), .A2(b[5]), .ZN(n500) );
  INVD0 U1116 ( .I(n501), .ZN(n[187]) );
  ND2D0 U1117 ( .A1(n[60]), .A2(b[5]), .ZN(n501) );
  INVD0 U1118 ( .I(n502), .ZN(n[186]) );
  ND2D0 U1119 ( .A1(n[59]), .A2(b[5]), .ZN(n502) );
  INVD0 U1120 ( .I(n503), .ZN(n[185]) );
  ND2D0 U1121 ( .A1(n[58]), .A2(b[5]), .ZN(n503) );
  INVD0 U1122 ( .I(n504), .ZN(n[184]) );
  ND2D0 U1123 ( .A1(n[57]), .A2(b[5]), .ZN(n504) );
  INVD0 U1124 ( .I(n505), .ZN(n[183]) );
  ND2D0 U1125 ( .A1(n[56]), .A2(b[5]), .ZN(n505) );
  INVD0 U1126 ( .I(n506), .ZN(n[182]) );
  ND2D0 U1127 ( .A1(a[5]), .A2(n[118]), .ZN(n506) );
  INVD0 U1128 ( .I(n507), .ZN(n[181]) );
  ND2D0 U1129 ( .A1(a[5]), .A2(n[117]), .ZN(n507) );
  INVD0 U1130 ( .I(n508), .ZN(n[180]) );
  ND2D0 U1131 ( .A1(a[5]), .A2(n[116]), .ZN(n508) );
  INVD0 U1132 ( .I(n579), .ZN(n[17]) );
  INVD0 U1133 ( .I(n509), .ZN(n[179]) );
  ND2D0 U1134 ( .A1(a[5]), .A2(n[115]), .ZN(n509) );
  INVD0 U1135 ( .I(n510), .ZN(n[178]) );
  ND2D0 U1136 ( .A1(a[5]), .A2(n[114]), .ZN(n510) );
  INVD0 U1137 ( .I(n511), .ZN(n[177]) );
  ND2D0 U1138 ( .A1(a[5]), .A2(n[113]), .ZN(n511) );
  INVD0 U1139 ( .I(n512), .ZN(n[176]) );
  ND2D0 U1140 ( .A1(a[5]), .A2(n[112]), .ZN(n512) );
  INVD0 U1141 ( .I(n513), .ZN(n[175]) );
  ND2D0 U1142 ( .A1(a[5]), .A2(n[111]), .ZN(n513) );
  INVD0 U1143 ( .I(n514), .ZN(n[174]) );
  ND2D0 U1144 ( .A1(a[5]), .A2(n[110]), .ZN(n514) );
  INVD0 U1145 ( .I(n515), .ZN(n[173]) );
  ND2D0 U1146 ( .A1(a[5]), .A2(n[109]), .ZN(n515) );
  INVD0 U1147 ( .I(n516), .ZN(n[172]) );
  ND2D0 U1148 ( .A1(a[5]), .A2(n[108]), .ZN(n516) );
  INVD0 U1149 ( .I(n517), .ZN(n[171]) );
  ND2D0 U1150 ( .A1(a[5]), .A2(n[107]), .ZN(n517) );
  INVD0 U1151 ( .I(n518), .ZN(n[170]) );
  ND2D0 U1152 ( .A1(a[5]), .A2(n[106]), .ZN(n518) );
  INVD0 U1153 ( .I(n580), .ZN(n[16]) );
  INVD0 U1154 ( .I(n519), .ZN(n[169]) );
  ND2D0 U1155 ( .A1(a[5]), .A2(n[105]), .ZN(n519) );
  INVD0 U1156 ( .I(n520), .ZN(n[168]) );
  ND2D0 U1157 ( .A1(a[5]), .A2(n[104]), .ZN(n520) );
  INVD0 U1158 ( .I(n521), .ZN(n[167]) );
  ND2D0 U1159 ( .A1(a[5]), .A2(n[103]), .ZN(n521) );
  INVD0 U1160 ( .I(n522), .ZN(n[166]) );
  ND2D0 U1161 ( .A1(a[5]), .A2(n[102]), .ZN(n522) );
  INVD0 U1162 ( .I(n523), .ZN(n[165]) );
  ND2D0 U1163 ( .A1(a[5]), .A2(n[101]), .ZN(n523) );
  INVD0 U1164 ( .I(n524), .ZN(n[164]) );
  ND2D0 U1165 ( .A1(a[5]), .A2(n[100]), .ZN(n524) );
  INVD0 U1166 ( .I(n525), .ZN(n[163]) );
  ND2D0 U1167 ( .A1(a[5]), .A2(n[99]), .ZN(n525) );
  INVD0 U1168 ( .I(n581), .ZN(n[99]) );
  ND2D0 U1169 ( .A1(b[4]), .A2(n[36]), .ZN(n581) );
  INVD0 U1170 ( .I(n526), .ZN(n[162]) );
  ND2D0 U1171 ( .A1(a[5]), .A2(n[98]), .ZN(n526) );
  INVD0 U1172 ( .I(n582), .ZN(n[98]) );
  ND2D0 U1173 ( .A1(n[35]), .A2(b[4]), .ZN(n582) );
  INVD0 U1174 ( .I(n527), .ZN(n[161]) );
  ND2D0 U1175 ( .A1(a[5]), .A2(n[97]), .ZN(n527) );
  INVD0 U1176 ( .I(n583), .ZN(n[97]) );
  ND2D0 U1177 ( .A1(n[34]), .A2(b[4]), .ZN(n583) );
  INVD0 U1178 ( .I(n528), .ZN(n[160]) );
  ND2D0 U1179 ( .A1(a[5]), .A2(n[96]), .ZN(n528) );
  INVD0 U1180 ( .I(n584), .ZN(n[96]) );
  ND2D0 U1181 ( .A1(n[33]), .A2(b[4]), .ZN(n584) );
  INVD0 U1182 ( .I(n585), .ZN(n[15]) );
  INVD0 U1183 ( .I(n529), .ZN(n[159]) );
  ND2D0 U1184 ( .A1(a[5]), .A2(n[95]), .ZN(n529) );
  INVD0 U1185 ( .I(n586), .ZN(n[95]) );
  ND2D0 U1186 ( .A1(n[32]), .A2(b[4]), .ZN(n586) );
  INVD0 U1187 ( .I(n530), .ZN(n[158]) );
  ND2D0 U1188 ( .A1(a[5]), .A2(n[94]), .ZN(n530) );
  INVD0 U1189 ( .I(n587), .ZN(n[94]) );
  ND2D0 U1190 ( .A1(n[31]), .A2(b[4]), .ZN(n587) );
  INVD0 U1191 ( .I(n531), .ZN(n[157]) );
  ND2D0 U1192 ( .A1(a[5]), .A2(n[93]), .ZN(n531) );
  INVD0 U1193 ( .I(n588), .ZN(n[93]) );
  ND2D0 U1194 ( .A1(n[30]), .A2(b[4]), .ZN(n588) );
  INVD0 U1195 ( .I(n532), .ZN(n[156]) );
  ND2D0 U1196 ( .A1(a[5]), .A2(n[92]), .ZN(n532) );
  INVD0 U1197 ( .I(n589), .ZN(n[92]) );
  ND2D0 U1198 ( .A1(n[29]), .A2(b[4]), .ZN(n589) );
  INVD0 U1199 ( .I(n533), .ZN(n[155]) );
  ND2D0 U1200 ( .A1(a[5]), .A2(n[91]), .ZN(n533) );
  INVD0 U1201 ( .I(n590), .ZN(n[91]) );
  ND2D0 U1202 ( .A1(n[28]), .A2(b[4]), .ZN(n590) );
  INVD0 U1203 ( .I(n534), .ZN(n[154]) );
  ND2D0 U1204 ( .A1(a[5]), .A2(n[90]), .ZN(n534) );
  INVD0 U1205 ( .I(n591), .ZN(n[90]) );
  ND2D0 U1206 ( .A1(n[27]), .A2(b[4]), .ZN(n591) );
  INVD0 U1207 ( .I(n535), .ZN(n[153]) );
  ND2D0 U1208 ( .A1(a[5]), .A2(n[89]), .ZN(n535) );
  INVD0 U1209 ( .I(n592), .ZN(n[89]) );
  ND2D0 U1210 ( .A1(n[26]), .A2(b[4]), .ZN(n592) );
  INVD0 U1211 ( .I(n536), .ZN(n[152]) );
  ND2D0 U1212 ( .A1(a[5]), .A2(n[88]), .ZN(n536) );
  INVD0 U1213 ( .I(n593), .ZN(n[88]) );
  ND2D0 U1214 ( .A1(n[25]), .A2(b[4]), .ZN(n593) );
  INVD0 U1215 ( .I(n537), .ZN(n[151]) );
  ND2D0 U1216 ( .A1(a[5]), .A2(n[87]), .ZN(n537) );
  INVD0 U1217 ( .I(n594), .ZN(n[87]) );
  ND2D0 U1218 ( .A1(a[4]), .A2(n[55]), .ZN(n594) );
  INVD0 U1219 ( .I(n538), .ZN(n[150]) );
  ND2D0 U1220 ( .A1(a[5]), .A2(n[86]), .ZN(n538) );
  INVD0 U1221 ( .I(n595), .ZN(n[86]) );
  ND2D0 U1222 ( .A1(n[54]), .A2(a[4]), .ZN(n595) );
  INVD0 U1223 ( .I(n596), .ZN(n[14]) );
  INVD0 U1224 ( .I(n539), .ZN(n[149]) );
  ND2D0 U1225 ( .A1(a[5]), .A2(n[85]), .ZN(n539) );
  INVD0 U1226 ( .I(n597), .ZN(n[85]) );
  ND2D0 U1227 ( .A1(n[53]), .A2(a[4]), .ZN(n597) );
  INVD0 U1228 ( .I(n540), .ZN(n[148]) );
  ND2D0 U1229 ( .A1(a[5]), .A2(n[84]), .ZN(n540) );
  INVD0 U1230 ( .I(n598), .ZN(n[84]) );
  ND2D0 U1231 ( .A1(n[52]), .A2(a[4]), .ZN(n598) );
  INVD0 U1232 ( .I(n541), .ZN(n[147]) );
  ND2D0 U1233 ( .A1(a[5]), .A2(n[83]), .ZN(n541) );
  INVD0 U1234 ( .I(n599), .ZN(n[83]) );
  ND2D0 U1235 ( .A1(n[51]), .A2(a[4]), .ZN(n599) );
  INVD0 U1236 ( .I(n542), .ZN(n[146]) );
  ND2D0 U1237 ( .A1(a[5]), .A2(n[82]), .ZN(n542) );
  INVD0 U1238 ( .I(n600), .ZN(n[82]) );
  ND2D0 U1239 ( .A1(n[50]), .A2(a[4]), .ZN(n600) );
  INVD0 U1240 ( .I(n543), .ZN(n[145]) );
  ND2D0 U1241 ( .A1(a[5]), .A2(n[81]), .ZN(n543) );
  INVD0 U1242 ( .I(n601), .ZN(n[81]) );
  ND2D0 U1243 ( .A1(n[49]), .A2(a[4]), .ZN(n601) );
  INVD0 U1244 ( .I(n544), .ZN(n[144]) );
  ND2D0 U1245 ( .A1(a[5]), .A2(n[80]), .ZN(n544) );
  INVD0 U1246 ( .I(n602), .ZN(n[80]) );
  ND2D0 U1247 ( .A1(n[48]), .A2(a[4]), .ZN(n602) );
  INVD0 U1248 ( .I(n545), .ZN(n[143]) );
  ND2D0 U1249 ( .A1(a[5]), .A2(n[79]), .ZN(n545) );
  INVD0 U1250 ( .I(n603), .ZN(n[79]) );
  ND2D0 U1251 ( .A1(n[47]), .A2(a[4]), .ZN(n603) );
  INVD0 U1252 ( .I(n546), .ZN(n[142]) );
  ND2D0 U1253 ( .A1(a[5]), .A2(n[78]), .ZN(n546) );
  INVD0 U1254 ( .I(n604), .ZN(n[78]) );
  ND2D0 U1255 ( .A1(n[46]), .A2(a[4]), .ZN(n604) );
  INVD0 U1256 ( .I(n547), .ZN(n[141]) );
  ND2D0 U1257 ( .A1(a[5]), .A2(n[77]), .ZN(n547) );
  INVD0 U1258 ( .I(n605), .ZN(n[77]) );
  ND2D0 U1259 ( .A1(n[45]), .A2(a[4]), .ZN(n605) );
  INVD0 U1260 ( .I(n548), .ZN(n[140]) );
  ND2D0 U1261 ( .A1(a[5]), .A2(n[76]), .ZN(n548) );
  INVD0 U1262 ( .I(n606), .ZN(n[76]) );
  ND2D0 U1263 ( .A1(n[44]), .A2(a[4]), .ZN(n606) );
  INVD0 U1264 ( .I(n607), .ZN(n[13]) );
  INVD0 U1265 ( .I(n549), .ZN(n[139]) );
  ND2D0 U1266 ( .A1(a[5]), .A2(n[75]), .ZN(n549) );
  INVD0 U1267 ( .I(n608), .ZN(n[75]) );
  ND2D0 U1268 ( .A1(n[43]), .A2(a[4]), .ZN(n608) );
  INVD0 U1269 ( .I(n550), .ZN(n[138]) );
  ND2D0 U1270 ( .A1(a[5]), .A2(n[74]), .ZN(n550) );
  INVD0 U1271 ( .I(n609), .ZN(n[74]) );
  ND2D0 U1272 ( .A1(n[42]), .A2(a[4]), .ZN(n609) );
  INVD0 U1273 ( .I(n551), .ZN(n[137]) );
  ND2D0 U1274 ( .A1(a[5]), .A2(n[73]), .ZN(n551) );
  INVD0 U1275 ( .I(n610), .ZN(n[73]) );
  ND2D0 U1276 ( .A1(n[41]), .A2(a[4]), .ZN(n610) );
  INVD0 U1277 ( .I(n552), .ZN(n[136]) );
  ND2D0 U1278 ( .A1(a[5]), .A2(n[72]), .ZN(n552) );
  INVD0 U1279 ( .I(n611), .ZN(n[72]) );
  ND2D0 U1280 ( .A1(n[40]), .A2(a[4]), .ZN(n611) );
  INVD0 U1281 ( .I(n553), .ZN(n[135]) );
  ND2D0 U1282 ( .A1(a[5]), .A2(n[71]), .ZN(n553) );
  INVD0 U1283 ( .I(n612), .ZN(n[71]) );
  ND2D0 U1284 ( .A1(n[39]), .A2(a[4]), .ZN(n612) );
  INVD0 U1285 ( .I(n554), .ZN(n[134]) );
  ND2D0 U1286 ( .A1(a[5]), .A2(n[70]), .ZN(n554) );
  INVD0 U1287 ( .I(n613), .ZN(n[70]) );
  ND2D0 U1288 ( .A1(n[38]), .A2(a[4]), .ZN(n613) );
  INVD0 U1289 ( .I(n555), .ZN(n[133]) );
  ND2D0 U1290 ( .A1(a[5]), .A2(n[69]), .ZN(n555) );
  INVD0 U1291 ( .I(n614), .ZN(n[69]) );
  ND2D0 U1292 ( .A1(n[37]), .A2(a[4]), .ZN(n614) );
  INVD0 U1293 ( .I(n556), .ZN(n[132]) );
  ND2D0 U1294 ( .A1(a[5]), .A2(n[68]), .ZN(n556) );
  INVD0 U1295 ( .I(n615), .ZN(n[68]) );
  ND2D0 U1296 ( .A1(a[4]), .A2(n[36]), .ZN(n615) );
  NR2D0 U1297 ( .A1(n616), .A2(n575), .ZN(n[36]) );
  INVD0 U1298 ( .I(n557), .ZN(n[131]) );
  ND2D0 U1299 ( .A1(a[5]), .A2(n[67]), .ZN(n557) );
  INVD0 U1300 ( .I(n617), .ZN(n[67]) );
  ND2D0 U1301 ( .A1(a[4]), .A2(n[35]), .ZN(n617) );
  NR2D0 U1302 ( .A1(n577), .A2(n616), .ZN(n[35]) );
  INVD0 U1303 ( .I(n558), .ZN(n[130]) );
  ND2D0 U1304 ( .A1(a[5]), .A2(n[66]), .ZN(n558) );
  INVD0 U1305 ( .I(n618), .ZN(n[66]) );
  ND2D0 U1306 ( .A1(a[4]), .A2(n[34]), .ZN(n618) );
  NR2D0 U1307 ( .A1(n578), .A2(n616), .ZN(n[34]) );
  INVD0 U1308 ( .I(n619), .ZN(n[12]) );
  INVD0 U1309 ( .I(n559), .ZN(n[129]) );
  ND2D0 U1310 ( .A1(a[5]), .A2(n[65]), .ZN(n559) );
  INVD0 U1311 ( .I(n620), .ZN(n[65]) );
  ND2D0 U1312 ( .A1(a[4]), .A2(n[33]), .ZN(n620) );
  NR2D0 U1313 ( .A1(n579), .A2(n616), .ZN(n[33]) );
  INVD0 U1314 ( .I(n560), .ZN(n[128]) );
  ND2D0 U1315 ( .A1(a[5]), .A2(n[64]), .ZN(n560) );
  INVD0 U1316 ( .I(n621), .ZN(n[64]) );
  ND2D0 U1317 ( .A1(a[4]), .A2(n[32]), .ZN(n621) );
  NR2D0 U1318 ( .A1(n580), .A2(n616), .ZN(n[32]) );
  INVD0 U1319 ( .I(n561), .ZN(n[127]) );
  ND2D0 U1320 ( .A1(a[5]), .A2(n[63]), .ZN(n561) );
  INVD0 U1321 ( .I(n622), .ZN(n[63]) );
  ND2D0 U1322 ( .A1(a[4]), .A2(n[31]), .ZN(n622) );
  NR2D0 U1323 ( .A1(n585), .A2(n616), .ZN(n[31]) );
  INVD0 U1324 ( .I(n562), .ZN(n[126]) );
  ND2D0 U1325 ( .A1(a[5]), .A2(n[62]), .ZN(n562) );
  INVD0 U1326 ( .I(n623), .ZN(n[62]) );
  ND2D0 U1327 ( .A1(a[4]), .A2(n[30]), .ZN(n623) );
  NR2D0 U1328 ( .A1(n596), .A2(n616), .ZN(n[30]) );
  INVD0 U1329 ( .I(n563), .ZN(n[125]) );
  ND2D0 U1330 ( .A1(a[5]), .A2(n[61]), .ZN(n563) );
  INVD0 U1331 ( .I(n624), .ZN(n[61]) );
  ND2D0 U1332 ( .A1(a[4]), .A2(n[29]), .ZN(n624) );
  NR2D0 U1333 ( .A1(n607), .A2(n616), .ZN(n[29]) );
  INVD0 U1334 ( .I(n564), .ZN(n[124]) );
  ND2D0 U1335 ( .A1(a[5]), .A2(n[60]), .ZN(n564) );
  INVD0 U1336 ( .I(n625), .ZN(n[60]) );
  ND2D0 U1337 ( .A1(a[4]), .A2(n[28]), .ZN(n625) );
  NR2D0 U1338 ( .A1(n619), .A2(n616), .ZN(n[28]) );
  INVD0 U1339 ( .I(n565), .ZN(n[123]) );
  ND2D0 U1340 ( .A1(a[5]), .A2(n[59]), .ZN(n565) );
  INVD0 U1341 ( .I(n626), .ZN(n[59]) );
  ND2D0 U1342 ( .A1(a[4]), .A2(n[27]), .ZN(n626) );
  NR2D0 U1343 ( .A1(n627), .A2(n616), .ZN(n[27]) );
  INVD0 U1344 ( .I(n566), .ZN(n[122]) );
  ND2D0 U1345 ( .A1(a[5]), .A2(n[58]), .ZN(n566) );
  INVD0 U1346 ( .I(n628), .ZN(n[58]) );
  ND2D0 U1347 ( .A1(a[4]), .A2(n[26]), .ZN(n628) );
  NR2D0 U1348 ( .A1(n629), .A2(n616), .ZN(n[26]) );
  INVD0 U1349 ( .I(n567), .ZN(n[121]) );
  ND2D0 U1350 ( .A1(a[5]), .A2(n[57]), .ZN(n567) );
  INVD0 U1351 ( .I(n630), .ZN(n[57]) );
  ND2D0 U1352 ( .A1(a[4]), .A2(n[25]), .ZN(n630) );
  NR2D0 U1353 ( .A1(n631), .A2(n616), .ZN(n[25]) );
  INVD0 U1354 ( .I(n568), .ZN(n[120]) );
  ND2D0 U1355 ( .A1(a[5]), .A2(n[56]), .ZN(n568) );
  INVD0 U1356 ( .I(n632), .ZN(n[56]) );
  ND2D0 U1357 ( .A1(a[4]), .A2(b[4]), .ZN(n632) );
  INVD0 U1358 ( .I(n627), .ZN(n[11]) );
  INVD0 U1359 ( .I(n569), .ZN(n[119]) );
  ND2D0 U1360 ( .A1(a[5]), .A2(b[5]), .ZN(n569) );
  INVD0 U1361 ( .I(n633), .ZN(n[118]) );
  ND2D0 U1362 ( .A1(n[55]), .A2(b[4]), .ZN(n633) );
  NR2D0 U1363 ( .A1(n571), .A2(n631), .ZN(n[55]) );
  INVD0 U1364 ( .I(n634), .ZN(n[117]) );
  ND2D0 U1365 ( .A1(n[54]), .A2(b[4]), .ZN(n634) );
  NR2D0 U1366 ( .A1(n572), .A2(n631), .ZN(n[54]) );
  INVD0 U1367 ( .I(n635), .ZN(n[116]) );
  ND2D0 U1368 ( .A1(n[53]), .A2(b[4]), .ZN(n635) );
  NR2D0 U1369 ( .A1(n573), .A2(n631), .ZN(n[53]) );
  INVD0 U1370 ( .I(n636), .ZN(n[115]) );
  ND2D0 U1371 ( .A1(n[52]), .A2(b[4]), .ZN(n636) );
  NR2D0 U1372 ( .A1(n574), .A2(n631), .ZN(n[52]) );
  INVD0 U1373 ( .I(n637), .ZN(n[114]) );
  ND2D0 U1374 ( .A1(n[51]), .A2(b[4]), .ZN(n637) );
  NR2D0 U1375 ( .A1(n631), .A2(n575), .ZN(n[51]) );
  ND2D0 U1376 ( .A1(b[2]), .A2(n[5]), .ZN(n575) );
  INVD0 U1377 ( .I(n638), .ZN(n[113]) );
  ND2D0 U1378 ( .A1(n[50]), .A2(b[4]), .ZN(n638) );
  NR2D0 U1379 ( .A1(n631), .A2(n577), .ZN(n[50]) );
  ND2D0 U1380 ( .A1(n[4]), .A2(b[2]), .ZN(n577) );
  INVD0 U1381 ( .I(n639), .ZN(n[112]) );
  ND2D0 U1382 ( .A1(n[49]), .A2(b[4]), .ZN(n639) );
  NR2D0 U1383 ( .A1(n631), .A2(n578), .ZN(n[49]) );
  ND2D0 U1384 ( .A1(n[3]), .A2(b[2]), .ZN(n578) );
  INVD0 U1385 ( .I(n640), .ZN(n[111]) );
  ND2D0 U1386 ( .A1(n[48]), .A2(b[4]), .ZN(n640) );
  NR2D0 U1387 ( .A1(n631), .A2(n579), .ZN(n[48]) );
  ND2D0 U1388 ( .A1(a[2]), .A2(n[9]), .ZN(n579) );
  INVD0 U1389 ( .I(n641), .ZN(n[110]) );
  ND2D0 U1390 ( .A1(n[47]), .A2(b[4]), .ZN(n641) );
  NR2D0 U1391 ( .A1(n631), .A2(n580), .ZN(n[47]) );
  ND2D0 U1392 ( .A1(n[8]), .A2(a[2]), .ZN(n580) );
  INVD0 U1393 ( .I(n629), .ZN(n[10]) );
  INVD0 U1394 ( .I(n642), .ZN(n[109]) );
  ND2D0 U1395 ( .A1(n[46]), .A2(b[4]), .ZN(n642) );
  NR2D0 U1396 ( .A1(n631), .A2(n585), .ZN(n[46]) );
  ND2D0 U1397 ( .A1(n[7]), .A2(a[2]), .ZN(n585) );
  INVD0 U1398 ( .I(n643), .ZN(n[108]) );
  ND2D0 U1399 ( .A1(n[45]), .A2(b[4]), .ZN(n643) );
  NR2D0 U1400 ( .A1(n631), .A2(n596), .ZN(n[45]) );
  ND2D0 U1401 ( .A1(n[6]), .A2(a[2]), .ZN(n596) );
  INVD0 U1402 ( .I(n644), .ZN(n[107]) );
  ND2D0 U1403 ( .A1(n[44]), .A2(b[4]), .ZN(n644) );
  NR2D0 U1404 ( .A1(n631), .A2(n607), .ZN(n[44]) );
  ND2D0 U1405 ( .A1(a[2]), .A2(n[5]), .ZN(n607) );
  NR2D0 U1406 ( .A1(n645), .A2(n576), .ZN(n[5]) );
  INVD0 U1407 ( .I(n646), .ZN(n[106]) );
  ND2D0 U1408 ( .A1(n[43]), .A2(b[4]), .ZN(n646) );
  NR2D0 U1409 ( .A1(n631), .A2(n619), .ZN(n[43]) );
  ND2D0 U1410 ( .A1(a[2]), .A2(n[4]), .ZN(n619) );
  NR2D0 U1411 ( .A1(n647), .A2(n645), .ZN(n[4]) );
  INVD0 U1412 ( .I(n648), .ZN(n[105]) );
  ND2D0 U1413 ( .A1(n[42]), .A2(b[4]), .ZN(n648) );
  NR2D0 U1414 ( .A1(n631), .A2(n627), .ZN(n[42]) );
  ND2D0 U1415 ( .A1(a[2]), .A2(n[3]), .ZN(n627) );
  NR2D0 U1416 ( .A1(n645), .A2(n649), .ZN(n[3]) );
  INVD0 U1417 ( .I(n650), .ZN(n[104]) );
  ND2D0 U1418 ( .A1(n[41]), .A2(b[4]), .ZN(n650) );
  NR2D0 U1419 ( .A1(n631), .A2(n629), .ZN(n[41]) );
  ND2D0 U1420 ( .A1(a[2]), .A2(b[2]), .ZN(n629) );
  INVD0 U1421 ( .I(b[3]), .ZN(n631) );
  INVD0 U1422 ( .I(n651), .ZN(n[103]) );
  ND2D0 U1423 ( .A1(n[40]), .A2(b[4]), .ZN(n651) );
  NR2D0 U1424 ( .A1(n571), .A2(n616), .ZN(n[40]) );
  ND2D0 U1425 ( .A1(n[9]), .A2(b[2]), .ZN(n571) );
  NR2D0 U1426 ( .A1(n649), .A2(n570), .ZN(n[9]) );
  INVD0 U1427 ( .I(n652), .ZN(n[102]) );
  ND2D0 U1428 ( .A1(n[39]), .A2(b[4]), .ZN(n652) );
  NR2D0 U1429 ( .A1(n572), .A2(n616), .ZN(n[39]) );
  ND2D0 U1430 ( .A1(n[8]), .A2(b[2]), .ZN(n572) );
  NR2D0 U1431 ( .A1(n576), .A2(n649), .ZN(n[8]) );
  ND2D0 U1432 ( .A1(a[0]), .A2(c), .ZN(n576) );
  INVD0 U1433 ( .I(n653), .ZN(n[101]) );
  ND2D0 U1434 ( .A1(n[38]), .A2(b[4]), .ZN(n653) );
  NR2D0 U1435 ( .A1(n573), .A2(n616), .ZN(n[38]) );
  ND2D0 U1436 ( .A1(n[7]), .A2(b[2]), .ZN(n573) );
  NR2D0 U1437 ( .A1(n647), .A2(n649), .ZN(n[7]) );
  INVD0 U1438 ( .I(b[1]), .ZN(n649) );
  INVD0 U1439 ( .I(n654), .ZN(n[100]) );
  ND2D0 U1440 ( .A1(n[37]), .A2(b[4]), .ZN(n654) );
  NR2D0 U1441 ( .A1(n574), .A2(n616), .ZN(n[37]) );
  INVD0 U1442 ( .I(a[3]), .ZN(n616) );
  ND2D0 U1443 ( .A1(n[6]), .A2(b[2]), .ZN(n574) );
  NR2D0 U1444 ( .A1(n645), .A2(n570), .ZN(n[6]) );
  ND2D0 U1445 ( .A1(c), .A2(b[0]), .ZN(n570) );
  INVD0 U1446 ( .I(a[1]), .ZN(n645) );
  INVD0 U1447 ( .I(n647), .ZN(n[0]) );
  ND2D0 U1448 ( .A1(a[0]), .A2(b[0]), .ZN(n647) );
endmodule

