module gen_linear_part(a,b,n,s);

input  [11:0] a, b; //adder inputs
input [8176:0] n; // non-linear outputs
output [11:0] s;

wire [8176:0] t; // non-linear outputs
//asigning bit 0
assign s[0] = (a[0] ^ b[0]);
//asigning bit 1
assign t[0] = n[0];
assign t[1] = t[0] ^ n[1];
assign t[2] = t[1] ^ n[2];

assign s[1] = ( a[1] ^ b [1] ) ^ t[2];

//asigning bit 2
assign t[3] = n[3];
assign t[4] = t[3] ^ n[4];
assign t[5] = t[4] ^ n[5];
assign t[6] = t[5] ^ n[6];
assign t[7] = t[6] ^ n[7];
assign t[8] = t[7] ^ n[8];
assign t[9] = t[8] ^ n[9];

assign s[2] = ( a[2] ^ b [2] ) ^ t[9];

//asigning bit 3
assign t[10] = n[10];
assign t[11] = t[10] ^ n[11];
assign t[12] = t[11] ^ n[12];
assign t[13] = t[12] ^ n[13];
assign t[14] = t[13] ^ n[14];
assign t[15] = t[14] ^ n[15];
assign t[16] = t[15] ^ n[16];
assign t[17] = t[16] ^ n[17];
assign t[18] = t[17] ^ n[18];
assign t[19] = t[18] ^ n[19];
assign t[20] = t[19] ^ n[20];
assign t[21] = t[20] ^ n[21];
assign t[22] = t[21] ^ n[22];
assign t[23] = t[22] ^ n[23];
assign t[24] = t[23] ^ n[24];

assign s[3] = ( a[3] ^ b [3] ) ^ t[24];

//asigning bit 4
assign t[25] = n[25];
assign t[26] = t[25] ^ n[26];
assign t[27] = t[26] ^ n[27];
assign t[28] = t[27] ^ n[28];
assign t[29] = t[28] ^ n[29];
assign t[30] = t[29] ^ n[30];
assign t[31] = t[30] ^ n[31];
assign t[32] = t[31] ^ n[32];
assign t[33] = t[32] ^ n[33];
assign t[34] = t[33] ^ n[34];
assign t[35] = t[34] ^ n[35];
assign t[36] = t[35] ^ n[36];
assign t[37] = t[36] ^ n[37];
assign t[38] = t[37] ^ n[38];
assign t[39] = t[38] ^ n[39];
assign t[40] = t[39] ^ n[40];
assign t[41] = t[40] ^ n[41];
assign t[42] = t[41] ^ n[42];
assign t[43] = t[42] ^ n[43];
assign t[44] = t[43] ^ n[44];
assign t[45] = t[44] ^ n[45];
assign t[46] = t[45] ^ n[46];
assign t[47] = t[46] ^ n[47];
assign t[48] = t[47] ^ n[48];
assign t[49] = t[48] ^ n[49];
assign t[50] = t[49] ^ n[50];
assign t[51] = t[50] ^ n[51];
assign t[52] = t[51] ^ n[52];
assign t[53] = t[52] ^ n[53];
assign t[54] = t[53] ^ n[54];
assign t[55] = t[54] ^ n[55];

assign s[4] = ( a[4] ^ b [4] ) ^ t[55];

//asigning bit 5
assign t[56] = n[56];
assign t[57] = t[56] ^ n[57];
assign t[58] = t[57] ^ n[58];
assign t[59] = t[58] ^ n[59];
assign t[60] = t[59] ^ n[60];
assign t[61] = t[60] ^ n[61];
assign t[62] = t[61] ^ n[62];
assign t[63] = t[62] ^ n[63];
assign t[64] = t[63] ^ n[64];
assign t[65] = t[64] ^ n[65];
assign t[66] = t[65] ^ n[66];
assign t[67] = t[66] ^ n[67];
assign t[68] = t[67] ^ n[68];
assign t[69] = t[68] ^ n[69];
assign t[70] = t[69] ^ n[70];
assign t[71] = t[70] ^ n[71];
assign t[72] = t[71] ^ n[72];
assign t[73] = t[72] ^ n[73];
assign t[74] = t[73] ^ n[74];
assign t[75] = t[74] ^ n[75];
assign t[76] = t[75] ^ n[76];
assign t[77] = t[76] ^ n[77];
assign t[78] = t[77] ^ n[78];
assign t[79] = t[78] ^ n[79];
assign t[80] = t[79] ^ n[80];
assign t[81] = t[80] ^ n[81];
assign t[82] = t[81] ^ n[82];
assign t[83] = t[82] ^ n[83];
assign t[84] = t[83] ^ n[84];
assign t[85] = t[84] ^ n[85];
assign t[86] = t[85] ^ n[86];
assign t[87] = t[86] ^ n[87];
assign t[88] = t[87] ^ n[88];
assign t[89] = t[88] ^ n[89];
assign t[90] = t[89] ^ n[90];
assign t[91] = t[90] ^ n[91];
assign t[92] = t[91] ^ n[92];
assign t[93] = t[92] ^ n[93];
assign t[94] = t[93] ^ n[94];
assign t[95] = t[94] ^ n[95];
assign t[96] = t[95] ^ n[96];
assign t[97] = t[96] ^ n[97];
assign t[98] = t[97] ^ n[98];
assign t[99] = t[98] ^ n[99];
assign t[100] = t[99] ^ n[100];
assign t[101] = t[100] ^ n[101];
assign t[102] = t[101] ^ n[102];
assign t[103] = t[102] ^ n[103];
assign t[104] = t[103] ^ n[104];
assign t[105] = t[104] ^ n[105];
assign t[106] = t[105] ^ n[106];
assign t[107] = t[106] ^ n[107];
assign t[108] = t[107] ^ n[108];
assign t[109] = t[108] ^ n[109];
assign t[110] = t[109] ^ n[110];
assign t[111] = t[110] ^ n[111];
assign t[112] = t[111] ^ n[112];
assign t[113] = t[112] ^ n[113];
assign t[114] = t[113] ^ n[114];
assign t[115] = t[114] ^ n[115];
assign t[116] = t[115] ^ n[116];
assign t[117] = t[116] ^ n[117];
assign t[118] = t[117] ^ n[118];

assign s[5] = ( a[5] ^ b [5] ) ^ t[118];

//asigning bit 6
assign t[119] = n[119];
assign t[120] = t[119] ^ n[120];
assign t[121] = t[120] ^ n[121];
assign t[122] = t[121] ^ n[122];
assign t[123] = t[122] ^ n[123];
assign t[124] = t[123] ^ n[124];
assign t[125] = t[124] ^ n[125];
assign t[126] = t[125] ^ n[126];
assign t[127] = t[126] ^ n[127];
assign t[128] = t[127] ^ n[128];
assign t[129] = t[128] ^ n[129];
assign t[130] = t[129] ^ n[130];
assign t[131] = t[130] ^ n[131];
assign t[132] = t[131] ^ n[132];
assign t[133] = t[132] ^ n[133];
assign t[134] = t[133] ^ n[134];
assign t[135] = t[134] ^ n[135];
assign t[136] = t[135] ^ n[136];
assign t[137] = t[136] ^ n[137];
assign t[138] = t[137] ^ n[138];
assign t[139] = t[138] ^ n[139];
assign t[140] = t[139] ^ n[140];
assign t[141] = t[140] ^ n[141];
assign t[142] = t[141] ^ n[142];
assign t[143] = t[142] ^ n[143];
assign t[144] = t[143] ^ n[144];
assign t[145] = t[144] ^ n[145];
assign t[146] = t[145] ^ n[146];
assign t[147] = t[146] ^ n[147];
assign t[148] = t[147] ^ n[148];
assign t[149] = t[148] ^ n[149];
assign t[150] = t[149] ^ n[150];
assign t[151] = t[150] ^ n[151];
assign t[152] = t[151] ^ n[152];
assign t[153] = t[152] ^ n[153];
assign t[154] = t[153] ^ n[154];
assign t[155] = t[154] ^ n[155];
assign t[156] = t[155] ^ n[156];
assign t[157] = t[156] ^ n[157];
assign t[158] = t[157] ^ n[158];
assign t[159] = t[158] ^ n[159];
assign t[160] = t[159] ^ n[160];
assign t[161] = t[160] ^ n[161];
assign t[162] = t[161] ^ n[162];
assign t[163] = t[162] ^ n[163];
assign t[164] = t[163] ^ n[164];
assign t[165] = t[164] ^ n[165];
assign t[166] = t[165] ^ n[166];
assign t[167] = t[166] ^ n[167];
assign t[168] = t[167] ^ n[168];
assign t[169] = t[168] ^ n[169];
assign t[170] = t[169] ^ n[170];
assign t[171] = t[170] ^ n[171];
assign t[172] = t[171] ^ n[172];
assign t[173] = t[172] ^ n[173];
assign t[174] = t[173] ^ n[174];
assign t[175] = t[174] ^ n[175];
assign t[176] = t[175] ^ n[176];
assign t[177] = t[176] ^ n[177];
assign t[178] = t[177] ^ n[178];
assign t[179] = t[178] ^ n[179];
assign t[180] = t[179] ^ n[180];
assign t[181] = t[180] ^ n[181];
assign t[182] = t[181] ^ n[182];
assign t[183] = t[182] ^ n[183];
assign t[184] = t[183] ^ n[184];
assign t[185] = t[184] ^ n[185];
assign t[186] = t[185] ^ n[186];
assign t[187] = t[186] ^ n[187];
assign t[188] = t[187] ^ n[188];
assign t[189] = t[188] ^ n[189];
assign t[190] = t[189] ^ n[190];
assign t[191] = t[190] ^ n[191];
assign t[192] = t[191] ^ n[192];
assign t[193] = t[192] ^ n[193];
assign t[194] = t[193] ^ n[194];
assign t[195] = t[194] ^ n[195];
assign t[196] = t[195] ^ n[196];
assign t[197] = t[196] ^ n[197];
assign t[198] = t[197] ^ n[198];
assign t[199] = t[198] ^ n[199];
assign t[200] = t[199] ^ n[200];
assign t[201] = t[200] ^ n[201];
assign t[202] = t[201] ^ n[202];
assign t[203] = t[202] ^ n[203];
assign t[204] = t[203] ^ n[204];
assign t[205] = t[204] ^ n[205];
assign t[206] = t[205] ^ n[206];
assign t[207] = t[206] ^ n[207];
assign t[208] = t[207] ^ n[208];
assign t[209] = t[208] ^ n[209];
assign t[210] = t[209] ^ n[210];
assign t[211] = t[210] ^ n[211];
assign t[212] = t[211] ^ n[212];
assign t[213] = t[212] ^ n[213];
assign t[214] = t[213] ^ n[214];
assign t[215] = t[214] ^ n[215];
assign t[216] = t[215] ^ n[216];
assign t[217] = t[216] ^ n[217];
assign t[218] = t[217] ^ n[218];
assign t[219] = t[218] ^ n[219];
assign t[220] = t[219] ^ n[220];
assign t[221] = t[220] ^ n[221];
assign t[222] = t[221] ^ n[222];
assign t[223] = t[222] ^ n[223];
assign t[224] = t[223] ^ n[224];
assign t[225] = t[224] ^ n[225];
assign t[226] = t[225] ^ n[226];
assign t[227] = t[226] ^ n[227];
assign t[228] = t[227] ^ n[228];
assign t[229] = t[228] ^ n[229];
assign t[230] = t[229] ^ n[230];
assign t[231] = t[230] ^ n[231];
assign t[232] = t[231] ^ n[232];
assign t[233] = t[232] ^ n[233];
assign t[234] = t[233] ^ n[234];
assign t[235] = t[234] ^ n[235];
assign t[236] = t[235] ^ n[236];
assign t[237] = t[236] ^ n[237];
assign t[238] = t[237] ^ n[238];
assign t[239] = t[238] ^ n[239];
assign t[240] = t[239] ^ n[240];
assign t[241] = t[240] ^ n[241];
assign t[242] = t[241] ^ n[242];
assign t[243] = t[242] ^ n[243];
assign t[244] = t[243] ^ n[244];
assign t[245] = t[244] ^ n[245];

assign s[6] = ( a[6] ^ b [6] ) ^ t[245];

//asigning bit 7
assign t[246] = n[246];
assign t[247] = t[246] ^ n[247];
assign t[248] = t[247] ^ n[248];
assign t[249] = t[248] ^ n[249];
assign t[250] = t[249] ^ n[250];
assign t[251] = t[250] ^ n[251];
assign t[252] = t[251] ^ n[252];
assign t[253] = t[252] ^ n[253];
assign t[254] = t[253] ^ n[254];
assign t[255] = t[254] ^ n[255];
assign t[256] = t[255] ^ n[256];
assign t[257] = t[256] ^ n[257];
assign t[258] = t[257] ^ n[258];
assign t[259] = t[258] ^ n[259];
assign t[260] = t[259] ^ n[260];
assign t[261] = t[260] ^ n[261];
assign t[262] = t[261] ^ n[262];
assign t[263] = t[262] ^ n[263];
assign t[264] = t[263] ^ n[264];
assign t[265] = t[264] ^ n[265];
assign t[266] = t[265] ^ n[266];
assign t[267] = t[266] ^ n[267];
assign t[268] = t[267] ^ n[268];
assign t[269] = t[268] ^ n[269];
assign t[270] = t[269] ^ n[270];
assign t[271] = t[270] ^ n[271];
assign t[272] = t[271] ^ n[272];
assign t[273] = t[272] ^ n[273];
assign t[274] = t[273] ^ n[274];
assign t[275] = t[274] ^ n[275];
assign t[276] = t[275] ^ n[276];
assign t[277] = t[276] ^ n[277];
assign t[278] = t[277] ^ n[278];
assign t[279] = t[278] ^ n[279];
assign t[280] = t[279] ^ n[280];
assign t[281] = t[280] ^ n[281];
assign t[282] = t[281] ^ n[282];
assign t[283] = t[282] ^ n[283];
assign t[284] = t[283] ^ n[284];
assign t[285] = t[284] ^ n[285];
assign t[286] = t[285] ^ n[286];
assign t[287] = t[286] ^ n[287];
assign t[288] = t[287] ^ n[288];
assign t[289] = t[288] ^ n[289];
assign t[290] = t[289] ^ n[290];
assign t[291] = t[290] ^ n[291];
assign t[292] = t[291] ^ n[292];
assign t[293] = t[292] ^ n[293];
assign t[294] = t[293] ^ n[294];
assign t[295] = t[294] ^ n[295];
assign t[296] = t[295] ^ n[296];
assign t[297] = t[296] ^ n[297];
assign t[298] = t[297] ^ n[298];
assign t[299] = t[298] ^ n[299];
assign t[300] = t[299] ^ n[300];
assign t[301] = t[300] ^ n[301];
assign t[302] = t[301] ^ n[302];
assign t[303] = t[302] ^ n[303];
assign t[304] = t[303] ^ n[304];
assign t[305] = t[304] ^ n[305];
assign t[306] = t[305] ^ n[306];
assign t[307] = t[306] ^ n[307];
assign t[308] = t[307] ^ n[308];
assign t[309] = t[308] ^ n[309];
assign t[310] = t[309] ^ n[310];
assign t[311] = t[310] ^ n[311];
assign t[312] = t[311] ^ n[312];
assign t[313] = t[312] ^ n[313];
assign t[314] = t[313] ^ n[314];
assign t[315] = t[314] ^ n[315];
assign t[316] = t[315] ^ n[316];
assign t[317] = t[316] ^ n[317];
assign t[318] = t[317] ^ n[318];
assign t[319] = t[318] ^ n[319];
assign t[320] = t[319] ^ n[320];
assign t[321] = t[320] ^ n[321];
assign t[322] = t[321] ^ n[322];
assign t[323] = t[322] ^ n[323];
assign t[324] = t[323] ^ n[324];
assign t[325] = t[324] ^ n[325];
assign t[326] = t[325] ^ n[326];
assign t[327] = t[326] ^ n[327];
assign t[328] = t[327] ^ n[328];
assign t[329] = t[328] ^ n[329];
assign t[330] = t[329] ^ n[330];
assign t[331] = t[330] ^ n[331];
assign t[332] = t[331] ^ n[332];
assign t[333] = t[332] ^ n[333];
assign t[334] = t[333] ^ n[334];
assign t[335] = t[334] ^ n[335];
assign t[336] = t[335] ^ n[336];
assign t[337] = t[336] ^ n[337];
assign t[338] = t[337] ^ n[338];
assign t[339] = t[338] ^ n[339];
assign t[340] = t[339] ^ n[340];
assign t[341] = t[340] ^ n[341];
assign t[342] = t[341] ^ n[342];
assign t[343] = t[342] ^ n[343];
assign t[344] = t[343] ^ n[344];
assign t[345] = t[344] ^ n[345];
assign t[346] = t[345] ^ n[346];
assign t[347] = t[346] ^ n[347];
assign t[348] = t[347] ^ n[348];
assign t[349] = t[348] ^ n[349];
assign t[350] = t[349] ^ n[350];
assign t[351] = t[350] ^ n[351];
assign t[352] = t[351] ^ n[352];
assign t[353] = t[352] ^ n[353];
assign t[354] = t[353] ^ n[354];
assign t[355] = t[354] ^ n[355];
assign t[356] = t[355] ^ n[356];
assign t[357] = t[356] ^ n[357];
assign t[358] = t[357] ^ n[358];
assign t[359] = t[358] ^ n[359];
assign t[360] = t[359] ^ n[360];
assign t[361] = t[360] ^ n[361];
assign t[362] = t[361] ^ n[362];
assign t[363] = t[362] ^ n[363];
assign t[364] = t[363] ^ n[364];
assign t[365] = t[364] ^ n[365];
assign t[366] = t[365] ^ n[366];
assign t[367] = t[366] ^ n[367];
assign t[368] = t[367] ^ n[368];
assign t[369] = t[368] ^ n[369];
assign t[370] = t[369] ^ n[370];
assign t[371] = t[370] ^ n[371];
assign t[372] = t[371] ^ n[372];
assign t[373] = t[372] ^ n[373];
assign t[374] = t[373] ^ n[374];
assign t[375] = t[374] ^ n[375];
assign t[376] = t[375] ^ n[376];
assign t[377] = t[376] ^ n[377];
assign t[378] = t[377] ^ n[378];
assign t[379] = t[378] ^ n[379];
assign t[380] = t[379] ^ n[380];
assign t[381] = t[380] ^ n[381];
assign t[382] = t[381] ^ n[382];
assign t[383] = t[382] ^ n[383];
assign t[384] = t[383] ^ n[384];
assign t[385] = t[384] ^ n[385];
assign t[386] = t[385] ^ n[386];
assign t[387] = t[386] ^ n[387];
assign t[388] = t[387] ^ n[388];
assign t[389] = t[388] ^ n[389];
assign t[390] = t[389] ^ n[390];
assign t[391] = t[390] ^ n[391];
assign t[392] = t[391] ^ n[392];
assign t[393] = t[392] ^ n[393];
assign t[394] = t[393] ^ n[394];
assign t[395] = t[394] ^ n[395];
assign t[396] = t[395] ^ n[396];
assign t[397] = t[396] ^ n[397];
assign t[398] = t[397] ^ n[398];
assign t[399] = t[398] ^ n[399];
assign t[400] = t[399] ^ n[400];
assign t[401] = t[400] ^ n[401];
assign t[402] = t[401] ^ n[402];
assign t[403] = t[402] ^ n[403];
assign t[404] = t[403] ^ n[404];
assign t[405] = t[404] ^ n[405];
assign t[406] = t[405] ^ n[406];
assign t[407] = t[406] ^ n[407];
assign t[408] = t[407] ^ n[408];
assign t[409] = t[408] ^ n[409];
assign t[410] = t[409] ^ n[410];
assign t[411] = t[410] ^ n[411];
assign t[412] = t[411] ^ n[412];
assign t[413] = t[412] ^ n[413];
assign t[414] = t[413] ^ n[414];
assign t[415] = t[414] ^ n[415];
assign t[416] = t[415] ^ n[416];
assign t[417] = t[416] ^ n[417];
assign t[418] = t[417] ^ n[418];
assign t[419] = t[418] ^ n[419];
assign t[420] = t[419] ^ n[420];
assign t[421] = t[420] ^ n[421];
assign t[422] = t[421] ^ n[422];
assign t[423] = t[422] ^ n[423];
assign t[424] = t[423] ^ n[424];
assign t[425] = t[424] ^ n[425];
assign t[426] = t[425] ^ n[426];
assign t[427] = t[426] ^ n[427];
assign t[428] = t[427] ^ n[428];
assign t[429] = t[428] ^ n[429];
assign t[430] = t[429] ^ n[430];
assign t[431] = t[430] ^ n[431];
assign t[432] = t[431] ^ n[432];
assign t[433] = t[432] ^ n[433];
assign t[434] = t[433] ^ n[434];
assign t[435] = t[434] ^ n[435];
assign t[436] = t[435] ^ n[436];
assign t[437] = t[436] ^ n[437];
assign t[438] = t[437] ^ n[438];
assign t[439] = t[438] ^ n[439];
assign t[440] = t[439] ^ n[440];
assign t[441] = t[440] ^ n[441];
assign t[442] = t[441] ^ n[442];
assign t[443] = t[442] ^ n[443];
assign t[444] = t[443] ^ n[444];
assign t[445] = t[444] ^ n[445];
assign t[446] = t[445] ^ n[446];
assign t[447] = t[446] ^ n[447];
assign t[448] = t[447] ^ n[448];
assign t[449] = t[448] ^ n[449];
assign t[450] = t[449] ^ n[450];
assign t[451] = t[450] ^ n[451];
assign t[452] = t[451] ^ n[452];
assign t[453] = t[452] ^ n[453];
assign t[454] = t[453] ^ n[454];
assign t[455] = t[454] ^ n[455];
assign t[456] = t[455] ^ n[456];
assign t[457] = t[456] ^ n[457];
assign t[458] = t[457] ^ n[458];
assign t[459] = t[458] ^ n[459];
assign t[460] = t[459] ^ n[460];
assign t[461] = t[460] ^ n[461];
assign t[462] = t[461] ^ n[462];
assign t[463] = t[462] ^ n[463];
assign t[464] = t[463] ^ n[464];
assign t[465] = t[464] ^ n[465];
assign t[466] = t[465] ^ n[466];
assign t[467] = t[466] ^ n[467];
assign t[468] = t[467] ^ n[468];
assign t[469] = t[468] ^ n[469];
assign t[470] = t[469] ^ n[470];
assign t[471] = t[470] ^ n[471];
assign t[472] = t[471] ^ n[472];
assign t[473] = t[472] ^ n[473];
assign t[474] = t[473] ^ n[474];
assign t[475] = t[474] ^ n[475];
assign t[476] = t[475] ^ n[476];
assign t[477] = t[476] ^ n[477];
assign t[478] = t[477] ^ n[478];
assign t[479] = t[478] ^ n[479];
assign t[480] = t[479] ^ n[480];
assign t[481] = t[480] ^ n[481];
assign t[482] = t[481] ^ n[482];
assign t[483] = t[482] ^ n[483];
assign t[484] = t[483] ^ n[484];
assign t[485] = t[484] ^ n[485];
assign t[486] = t[485] ^ n[486];
assign t[487] = t[486] ^ n[487];
assign t[488] = t[487] ^ n[488];
assign t[489] = t[488] ^ n[489];
assign t[490] = t[489] ^ n[490];
assign t[491] = t[490] ^ n[491];
assign t[492] = t[491] ^ n[492];
assign t[493] = t[492] ^ n[493];
assign t[494] = t[493] ^ n[494];
assign t[495] = t[494] ^ n[495];
assign t[496] = t[495] ^ n[496];
assign t[497] = t[496] ^ n[497];
assign t[498] = t[497] ^ n[498];
assign t[499] = t[498] ^ n[499];
assign t[500] = t[499] ^ n[500];

assign s[7] = ( a[7] ^ b [7] ) ^ t[500];

//asigning bit 8
assign t[501] = n[501];
assign t[502] = t[501] ^ n[502];
assign t[503] = t[502] ^ n[503];
assign t[504] = t[503] ^ n[504];
assign t[505] = t[504] ^ n[505];
assign t[506] = t[505] ^ n[506];
assign t[507] = t[506] ^ n[507];
assign t[508] = t[507] ^ n[508];
assign t[509] = t[508] ^ n[509];
assign t[510] = t[509] ^ n[510];
assign t[511] = t[510] ^ n[511];
assign t[512] = t[511] ^ n[512];
assign t[513] = t[512] ^ n[513];
assign t[514] = t[513] ^ n[514];
assign t[515] = t[514] ^ n[515];
assign t[516] = t[515] ^ n[516];
assign t[517] = t[516] ^ n[517];
assign t[518] = t[517] ^ n[518];
assign t[519] = t[518] ^ n[519];
assign t[520] = t[519] ^ n[520];
assign t[521] = t[520] ^ n[521];
assign t[522] = t[521] ^ n[522];
assign t[523] = t[522] ^ n[523];
assign t[524] = t[523] ^ n[524];
assign t[525] = t[524] ^ n[525];
assign t[526] = t[525] ^ n[526];
assign t[527] = t[526] ^ n[527];
assign t[528] = t[527] ^ n[528];
assign t[529] = t[528] ^ n[529];
assign t[530] = t[529] ^ n[530];
assign t[531] = t[530] ^ n[531];
assign t[532] = t[531] ^ n[532];
assign t[533] = t[532] ^ n[533];
assign t[534] = t[533] ^ n[534];
assign t[535] = t[534] ^ n[535];
assign t[536] = t[535] ^ n[536];
assign t[537] = t[536] ^ n[537];
assign t[538] = t[537] ^ n[538];
assign t[539] = t[538] ^ n[539];
assign t[540] = t[539] ^ n[540];
assign t[541] = t[540] ^ n[541];
assign t[542] = t[541] ^ n[542];
assign t[543] = t[542] ^ n[543];
assign t[544] = t[543] ^ n[544];
assign t[545] = t[544] ^ n[545];
assign t[546] = t[545] ^ n[546];
assign t[547] = t[546] ^ n[547];
assign t[548] = t[547] ^ n[548];
assign t[549] = t[548] ^ n[549];
assign t[550] = t[549] ^ n[550];
assign t[551] = t[550] ^ n[551];
assign t[552] = t[551] ^ n[552];
assign t[553] = t[552] ^ n[553];
assign t[554] = t[553] ^ n[554];
assign t[555] = t[554] ^ n[555];
assign t[556] = t[555] ^ n[556];
assign t[557] = t[556] ^ n[557];
assign t[558] = t[557] ^ n[558];
assign t[559] = t[558] ^ n[559];
assign t[560] = t[559] ^ n[560];
assign t[561] = t[560] ^ n[561];
assign t[562] = t[561] ^ n[562];
assign t[563] = t[562] ^ n[563];
assign t[564] = t[563] ^ n[564];
assign t[565] = t[564] ^ n[565];
assign t[566] = t[565] ^ n[566];
assign t[567] = t[566] ^ n[567];
assign t[568] = t[567] ^ n[568];
assign t[569] = t[568] ^ n[569];
assign t[570] = t[569] ^ n[570];
assign t[571] = t[570] ^ n[571];
assign t[572] = t[571] ^ n[572];
assign t[573] = t[572] ^ n[573];
assign t[574] = t[573] ^ n[574];
assign t[575] = t[574] ^ n[575];
assign t[576] = t[575] ^ n[576];
assign t[577] = t[576] ^ n[577];
assign t[578] = t[577] ^ n[578];
assign t[579] = t[578] ^ n[579];
assign t[580] = t[579] ^ n[580];
assign t[581] = t[580] ^ n[581];
assign t[582] = t[581] ^ n[582];
assign t[583] = t[582] ^ n[583];
assign t[584] = t[583] ^ n[584];
assign t[585] = t[584] ^ n[585];
assign t[586] = t[585] ^ n[586];
assign t[587] = t[586] ^ n[587];
assign t[588] = t[587] ^ n[588];
assign t[589] = t[588] ^ n[589];
assign t[590] = t[589] ^ n[590];
assign t[591] = t[590] ^ n[591];
assign t[592] = t[591] ^ n[592];
assign t[593] = t[592] ^ n[593];
assign t[594] = t[593] ^ n[594];
assign t[595] = t[594] ^ n[595];
assign t[596] = t[595] ^ n[596];
assign t[597] = t[596] ^ n[597];
assign t[598] = t[597] ^ n[598];
assign t[599] = t[598] ^ n[599];
assign t[600] = t[599] ^ n[600];
assign t[601] = t[600] ^ n[601];
assign t[602] = t[601] ^ n[602];
assign t[603] = t[602] ^ n[603];
assign t[604] = t[603] ^ n[604];
assign t[605] = t[604] ^ n[605];
assign t[606] = t[605] ^ n[606];
assign t[607] = t[606] ^ n[607];
assign t[608] = t[607] ^ n[608];
assign t[609] = t[608] ^ n[609];
assign t[610] = t[609] ^ n[610];
assign t[611] = t[610] ^ n[611];
assign t[612] = t[611] ^ n[612];
assign t[613] = t[612] ^ n[613];
assign t[614] = t[613] ^ n[614];
assign t[615] = t[614] ^ n[615];
assign t[616] = t[615] ^ n[616];
assign t[617] = t[616] ^ n[617];
assign t[618] = t[617] ^ n[618];
assign t[619] = t[618] ^ n[619];
assign t[620] = t[619] ^ n[620];
assign t[621] = t[620] ^ n[621];
assign t[622] = t[621] ^ n[622];
assign t[623] = t[622] ^ n[623];
assign t[624] = t[623] ^ n[624];
assign t[625] = t[624] ^ n[625];
assign t[626] = t[625] ^ n[626];
assign t[627] = t[626] ^ n[627];
assign t[628] = t[627] ^ n[628];
assign t[629] = t[628] ^ n[629];
assign t[630] = t[629] ^ n[630];
assign t[631] = t[630] ^ n[631];
assign t[632] = t[631] ^ n[632];
assign t[633] = t[632] ^ n[633];
assign t[634] = t[633] ^ n[634];
assign t[635] = t[634] ^ n[635];
assign t[636] = t[635] ^ n[636];
assign t[637] = t[636] ^ n[637];
assign t[638] = t[637] ^ n[638];
assign t[639] = t[638] ^ n[639];
assign t[640] = t[639] ^ n[640];
assign t[641] = t[640] ^ n[641];
assign t[642] = t[641] ^ n[642];
assign t[643] = t[642] ^ n[643];
assign t[644] = t[643] ^ n[644];
assign t[645] = t[644] ^ n[645];
assign t[646] = t[645] ^ n[646];
assign t[647] = t[646] ^ n[647];
assign t[648] = t[647] ^ n[648];
assign t[649] = t[648] ^ n[649];
assign t[650] = t[649] ^ n[650];
assign t[651] = t[650] ^ n[651];
assign t[652] = t[651] ^ n[652];
assign t[653] = t[652] ^ n[653];
assign t[654] = t[653] ^ n[654];
assign t[655] = t[654] ^ n[655];
assign t[656] = t[655] ^ n[656];
assign t[657] = t[656] ^ n[657];
assign t[658] = t[657] ^ n[658];
assign t[659] = t[658] ^ n[659];
assign t[660] = t[659] ^ n[660];
assign t[661] = t[660] ^ n[661];
assign t[662] = t[661] ^ n[662];
assign t[663] = t[662] ^ n[663];
assign t[664] = t[663] ^ n[664];
assign t[665] = t[664] ^ n[665];
assign t[666] = t[665] ^ n[666];
assign t[667] = t[666] ^ n[667];
assign t[668] = t[667] ^ n[668];
assign t[669] = t[668] ^ n[669];
assign t[670] = t[669] ^ n[670];
assign t[671] = t[670] ^ n[671];
assign t[672] = t[671] ^ n[672];
assign t[673] = t[672] ^ n[673];
assign t[674] = t[673] ^ n[674];
assign t[675] = t[674] ^ n[675];
assign t[676] = t[675] ^ n[676];
assign t[677] = t[676] ^ n[677];
assign t[678] = t[677] ^ n[678];
assign t[679] = t[678] ^ n[679];
assign t[680] = t[679] ^ n[680];
assign t[681] = t[680] ^ n[681];
assign t[682] = t[681] ^ n[682];
assign t[683] = t[682] ^ n[683];
assign t[684] = t[683] ^ n[684];
assign t[685] = t[684] ^ n[685];
assign t[686] = t[685] ^ n[686];
assign t[687] = t[686] ^ n[687];
assign t[688] = t[687] ^ n[688];
assign t[689] = t[688] ^ n[689];
assign t[690] = t[689] ^ n[690];
assign t[691] = t[690] ^ n[691];
assign t[692] = t[691] ^ n[692];
assign t[693] = t[692] ^ n[693];
assign t[694] = t[693] ^ n[694];
assign t[695] = t[694] ^ n[695];
assign t[696] = t[695] ^ n[696];
assign t[697] = t[696] ^ n[697];
assign t[698] = t[697] ^ n[698];
assign t[699] = t[698] ^ n[699];
assign t[700] = t[699] ^ n[700];
assign t[701] = t[700] ^ n[701];
assign t[702] = t[701] ^ n[702];
assign t[703] = t[702] ^ n[703];
assign t[704] = t[703] ^ n[704];
assign t[705] = t[704] ^ n[705];
assign t[706] = t[705] ^ n[706];
assign t[707] = t[706] ^ n[707];
assign t[708] = t[707] ^ n[708];
assign t[709] = t[708] ^ n[709];
assign t[710] = t[709] ^ n[710];
assign t[711] = t[710] ^ n[711];
assign t[712] = t[711] ^ n[712];
assign t[713] = t[712] ^ n[713];
assign t[714] = t[713] ^ n[714];
assign t[715] = t[714] ^ n[715];
assign t[716] = t[715] ^ n[716];
assign t[717] = t[716] ^ n[717];
assign t[718] = t[717] ^ n[718];
assign t[719] = t[718] ^ n[719];
assign t[720] = t[719] ^ n[720];
assign t[721] = t[720] ^ n[721];
assign t[722] = t[721] ^ n[722];
assign t[723] = t[722] ^ n[723];
assign t[724] = t[723] ^ n[724];
assign t[725] = t[724] ^ n[725];
assign t[726] = t[725] ^ n[726];
assign t[727] = t[726] ^ n[727];
assign t[728] = t[727] ^ n[728];
assign t[729] = t[728] ^ n[729];
assign t[730] = t[729] ^ n[730];
assign t[731] = t[730] ^ n[731];
assign t[732] = t[731] ^ n[732];
assign t[733] = t[732] ^ n[733];
assign t[734] = t[733] ^ n[734];
assign t[735] = t[734] ^ n[735];
assign t[736] = t[735] ^ n[736];
assign t[737] = t[736] ^ n[737];
assign t[738] = t[737] ^ n[738];
assign t[739] = t[738] ^ n[739];
assign t[740] = t[739] ^ n[740];
assign t[741] = t[740] ^ n[741];
assign t[742] = t[741] ^ n[742];
assign t[743] = t[742] ^ n[743];
assign t[744] = t[743] ^ n[744];
assign t[745] = t[744] ^ n[745];
assign t[746] = t[745] ^ n[746];
assign t[747] = t[746] ^ n[747];
assign t[748] = t[747] ^ n[748];
assign t[749] = t[748] ^ n[749];
assign t[750] = t[749] ^ n[750];
assign t[751] = t[750] ^ n[751];
assign t[752] = t[751] ^ n[752];
assign t[753] = t[752] ^ n[753];
assign t[754] = t[753] ^ n[754];
assign t[755] = t[754] ^ n[755];
assign t[756] = t[755] ^ n[756];
assign t[757] = t[756] ^ n[757];
assign t[758] = t[757] ^ n[758];
assign t[759] = t[758] ^ n[759];
assign t[760] = t[759] ^ n[760];
assign t[761] = t[760] ^ n[761];
assign t[762] = t[761] ^ n[762];
assign t[763] = t[762] ^ n[763];
assign t[764] = t[763] ^ n[764];
assign t[765] = t[764] ^ n[765];
assign t[766] = t[765] ^ n[766];
assign t[767] = t[766] ^ n[767];
assign t[768] = t[767] ^ n[768];
assign t[769] = t[768] ^ n[769];
assign t[770] = t[769] ^ n[770];
assign t[771] = t[770] ^ n[771];
assign t[772] = t[771] ^ n[772];
assign t[773] = t[772] ^ n[773];
assign t[774] = t[773] ^ n[774];
assign t[775] = t[774] ^ n[775];
assign t[776] = t[775] ^ n[776];
assign t[777] = t[776] ^ n[777];
assign t[778] = t[777] ^ n[778];
assign t[779] = t[778] ^ n[779];
assign t[780] = t[779] ^ n[780];
assign t[781] = t[780] ^ n[781];
assign t[782] = t[781] ^ n[782];
assign t[783] = t[782] ^ n[783];
assign t[784] = t[783] ^ n[784];
assign t[785] = t[784] ^ n[785];
assign t[786] = t[785] ^ n[786];
assign t[787] = t[786] ^ n[787];
assign t[788] = t[787] ^ n[788];
assign t[789] = t[788] ^ n[789];
assign t[790] = t[789] ^ n[790];
assign t[791] = t[790] ^ n[791];
assign t[792] = t[791] ^ n[792];
assign t[793] = t[792] ^ n[793];
assign t[794] = t[793] ^ n[794];
assign t[795] = t[794] ^ n[795];
assign t[796] = t[795] ^ n[796];
assign t[797] = t[796] ^ n[797];
assign t[798] = t[797] ^ n[798];
assign t[799] = t[798] ^ n[799];
assign t[800] = t[799] ^ n[800];
assign t[801] = t[800] ^ n[801];
assign t[802] = t[801] ^ n[802];
assign t[803] = t[802] ^ n[803];
assign t[804] = t[803] ^ n[804];
assign t[805] = t[804] ^ n[805];
assign t[806] = t[805] ^ n[806];
assign t[807] = t[806] ^ n[807];
assign t[808] = t[807] ^ n[808];
assign t[809] = t[808] ^ n[809];
assign t[810] = t[809] ^ n[810];
assign t[811] = t[810] ^ n[811];
assign t[812] = t[811] ^ n[812];
assign t[813] = t[812] ^ n[813];
assign t[814] = t[813] ^ n[814];
assign t[815] = t[814] ^ n[815];
assign t[816] = t[815] ^ n[816];
assign t[817] = t[816] ^ n[817];
assign t[818] = t[817] ^ n[818];
assign t[819] = t[818] ^ n[819];
assign t[820] = t[819] ^ n[820];
assign t[821] = t[820] ^ n[821];
assign t[822] = t[821] ^ n[822];
assign t[823] = t[822] ^ n[823];
assign t[824] = t[823] ^ n[824];
assign t[825] = t[824] ^ n[825];
assign t[826] = t[825] ^ n[826];
assign t[827] = t[826] ^ n[827];
assign t[828] = t[827] ^ n[828];
assign t[829] = t[828] ^ n[829];
assign t[830] = t[829] ^ n[830];
assign t[831] = t[830] ^ n[831];
assign t[832] = t[831] ^ n[832];
assign t[833] = t[832] ^ n[833];
assign t[834] = t[833] ^ n[834];
assign t[835] = t[834] ^ n[835];
assign t[836] = t[835] ^ n[836];
assign t[837] = t[836] ^ n[837];
assign t[838] = t[837] ^ n[838];
assign t[839] = t[838] ^ n[839];
assign t[840] = t[839] ^ n[840];
assign t[841] = t[840] ^ n[841];
assign t[842] = t[841] ^ n[842];
assign t[843] = t[842] ^ n[843];
assign t[844] = t[843] ^ n[844];
assign t[845] = t[844] ^ n[845];
assign t[846] = t[845] ^ n[846];
assign t[847] = t[846] ^ n[847];
assign t[848] = t[847] ^ n[848];
assign t[849] = t[848] ^ n[849];
assign t[850] = t[849] ^ n[850];
assign t[851] = t[850] ^ n[851];
assign t[852] = t[851] ^ n[852];
assign t[853] = t[852] ^ n[853];
assign t[854] = t[853] ^ n[854];
assign t[855] = t[854] ^ n[855];
assign t[856] = t[855] ^ n[856];
assign t[857] = t[856] ^ n[857];
assign t[858] = t[857] ^ n[858];
assign t[859] = t[858] ^ n[859];
assign t[860] = t[859] ^ n[860];
assign t[861] = t[860] ^ n[861];
assign t[862] = t[861] ^ n[862];
assign t[863] = t[862] ^ n[863];
assign t[864] = t[863] ^ n[864];
assign t[865] = t[864] ^ n[865];
assign t[866] = t[865] ^ n[866];
assign t[867] = t[866] ^ n[867];
assign t[868] = t[867] ^ n[868];
assign t[869] = t[868] ^ n[869];
assign t[870] = t[869] ^ n[870];
assign t[871] = t[870] ^ n[871];
assign t[872] = t[871] ^ n[872];
assign t[873] = t[872] ^ n[873];
assign t[874] = t[873] ^ n[874];
assign t[875] = t[874] ^ n[875];
assign t[876] = t[875] ^ n[876];
assign t[877] = t[876] ^ n[877];
assign t[878] = t[877] ^ n[878];
assign t[879] = t[878] ^ n[879];
assign t[880] = t[879] ^ n[880];
assign t[881] = t[880] ^ n[881];
assign t[882] = t[881] ^ n[882];
assign t[883] = t[882] ^ n[883];
assign t[884] = t[883] ^ n[884];
assign t[885] = t[884] ^ n[885];
assign t[886] = t[885] ^ n[886];
assign t[887] = t[886] ^ n[887];
assign t[888] = t[887] ^ n[888];
assign t[889] = t[888] ^ n[889];
assign t[890] = t[889] ^ n[890];
assign t[891] = t[890] ^ n[891];
assign t[892] = t[891] ^ n[892];
assign t[893] = t[892] ^ n[893];
assign t[894] = t[893] ^ n[894];
assign t[895] = t[894] ^ n[895];
assign t[896] = t[895] ^ n[896];
assign t[897] = t[896] ^ n[897];
assign t[898] = t[897] ^ n[898];
assign t[899] = t[898] ^ n[899];
assign t[900] = t[899] ^ n[900];
assign t[901] = t[900] ^ n[901];
assign t[902] = t[901] ^ n[902];
assign t[903] = t[902] ^ n[903];
assign t[904] = t[903] ^ n[904];
assign t[905] = t[904] ^ n[905];
assign t[906] = t[905] ^ n[906];
assign t[907] = t[906] ^ n[907];
assign t[908] = t[907] ^ n[908];
assign t[909] = t[908] ^ n[909];
assign t[910] = t[909] ^ n[910];
assign t[911] = t[910] ^ n[911];
assign t[912] = t[911] ^ n[912];
assign t[913] = t[912] ^ n[913];
assign t[914] = t[913] ^ n[914];
assign t[915] = t[914] ^ n[915];
assign t[916] = t[915] ^ n[916];
assign t[917] = t[916] ^ n[917];
assign t[918] = t[917] ^ n[918];
assign t[919] = t[918] ^ n[919];
assign t[920] = t[919] ^ n[920];
assign t[921] = t[920] ^ n[921];
assign t[922] = t[921] ^ n[922];
assign t[923] = t[922] ^ n[923];
assign t[924] = t[923] ^ n[924];
assign t[925] = t[924] ^ n[925];
assign t[926] = t[925] ^ n[926];
assign t[927] = t[926] ^ n[927];
assign t[928] = t[927] ^ n[928];
assign t[929] = t[928] ^ n[929];
assign t[930] = t[929] ^ n[930];
assign t[931] = t[930] ^ n[931];
assign t[932] = t[931] ^ n[932];
assign t[933] = t[932] ^ n[933];
assign t[934] = t[933] ^ n[934];
assign t[935] = t[934] ^ n[935];
assign t[936] = t[935] ^ n[936];
assign t[937] = t[936] ^ n[937];
assign t[938] = t[937] ^ n[938];
assign t[939] = t[938] ^ n[939];
assign t[940] = t[939] ^ n[940];
assign t[941] = t[940] ^ n[941];
assign t[942] = t[941] ^ n[942];
assign t[943] = t[942] ^ n[943];
assign t[944] = t[943] ^ n[944];
assign t[945] = t[944] ^ n[945];
assign t[946] = t[945] ^ n[946];
assign t[947] = t[946] ^ n[947];
assign t[948] = t[947] ^ n[948];
assign t[949] = t[948] ^ n[949];
assign t[950] = t[949] ^ n[950];
assign t[951] = t[950] ^ n[951];
assign t[952] = t[951] ^ n[952];
assign t[953] = t[952] ^ n[953];
assign t[954] = t[953] ^ n[954];
assign t[955] = t[954] ^ n[955];
assign t[956] = t[955] ^ n[956];
assign t[957] = t[956] ^ n[957];
assign t[958] = t[957] ^ n[958];
assign t[959] = t[958] ^ n[959];
assign t[960] = t[959] ^ n[960];
assign t[961] = t[960] ^ n[961];
assign t[962] = t[961] ^ n[962];
assign t[963] = t[962] ^ n[963];
assign t[964] = t[963] ^ n[964];
assign t[965] = t[964] ^ n[965];
assign t[966] = t[965] ^ n[966];
assign t[967] = t[966] ^ n[967];
assign t[968] = t[967] ^ n[968];
assign t[969] = t[968] ^ n[969];
assign t[970] = t[969] ^ n[970];
assign t[971] = t[970] ^ n[971];
assign t[972] = t[971] ^ n[972];
assign t[973] = t[972] ^ n[973];
assign t[974] = t[973] ^ n[974];
assign t[975] = t[974] ^ n[975];
assign t[976] = t[975] ^ n[976];
assign t[977] = t[976] ^ n[977];
assign t[978] = t[977] ^ n[978];
assign t[979] = t[978] ^ n[979];
assign t[980] = t[979] ^ n[980];
assign t[981] = t[980] ^ n[981];
assign t[982] = t[981] ^ n[982];
assign t[983] = t[982] ^ n[983];
assign t[984] = t[983] ^ n[984];
assign t[985] = t[984] ^ n[985];
assign t[986] = t[985] ^ n[986];
assign t[987] = t[986] ^ n[987];
assign t[988] = t[987] ^ n[988];
assign t[989] = t[988] ^ n[989];
assign t[990] = t[989] ^ n[990];
assign t[991] = t[990] ^ n[991];
assign t[992] = t[991] ^ n[992];
assign t[993] = t[992] ^ n[993];
assign t[994] = t[993] ^ n[994];
assign t[995] = t[994] ^ n[995];
assign t[996] = t[995] ^ n[996];
assign t[997] = t[996] ^ n[997];
assign t[998] = t[997] ^ n[998];
assign t[999] = t[998] ^ n[999];
assign t[1000] = t[999] ^ n[1000];
assign t[1001] = t[1000] ^ n[1001];
assign t[1002] = t[1001] ^ n[1002];
assign t[1003] = t[1002] ^ n[1003];
assign t[1004] = t[1003] ^ n[1004];
assign t[1005] = t[1004] ^ n[1005];
assign t[1006] = t[1005] ^ n[1006];
assign t[1007] = t[1006] ^ n[1007];
assign t[1008] = t[1007] ^ n[1008];
assign t[1009] = t[1008] ^ n[1009];
assign t[1010] = t[1009] ^ n[1010];
assign t[1011] = t[1010] ^ n[1011];

assign s[8] = ( a[8] ^ b [8] ) ^ t[1011];

//asigning bit 9
assign t[1012] = n[1012];
assign t[1013] = t[1012] ^ n[1013];
assign t[1014] = t[1013] ^ n[1014];
assign t[1015] = t[1014] ^ n[1015];
assign t[1016] = t[1015] ^ n[1016];
assign t[1017] = t[1016] ^ n[1017];
assign t[1018] = t[1017] ^ n[1018];
assign t[1019] = t[1018] ^ n[1019];
assign t[1020] = t[1019] ^ n[1020];
assign t[1021] = t[1020] ^ n[1021];
assign t[1022] = t[1021] ^ n[1022];
assign t[1023] = t[1022] ^ n[1023];
assign t[1024] = t[1023] ^ n[1024];
assign t[1025] = t[1024] ^ n[1025];
assign t[1026] = t[1025] ^ n[1026];
assign t[1027] = t[1026] ^ n[1027];
assign t[1028] = t[1027] ^ n[1028];
assign t[1029] = t[1028] ^ n[1029];
assign t[1030] = t[1029] ^ n[1030];
assign t[1031] = t[1030] ^ n[1031];
assign t[1032] = t[1031] ^ n[1032];
assign t[1033] = t[1032] ^ n[1033];
assign t[1034] = t[1033] ^ n[1034];
assign t[1035] = t[1034] ^ n[1035];
assign t[1036] = t[1035] ^ n[1036];
assign t[1037] = t[1036] ^ n[1037];
assign t[1038] = t[1037] ^ n[1038];
assign t[1039] = t[1038] ^ n[1039];
assign t[1040] = t[1039] ^ n[1040];
assign t[1041] = t[1040] ^ n[1041];
assign t[1042] = t[1041] ^ n[1042];
assign t[1043] = t[1042] ^ n[1043];
assign t[1044] = t[1043] ^ n[1044];
assign t[1045] = t[1044] ^ n[1045];
assign t[1046] = t[1045] ^ n[1046];
assign t[1047] = t[1046] ^ n[1047];
assign t[1048] = t[1047] ^ n[1048];
assign t[1049] = t[1048] ^ n[1049];
assign t[1050] = t[1049] ^ n[1050];
assign t[1051] = t[1050] ^ n[1051];
assign t[1052] = t[1051] ^ n[1052];
assign t[1053] = t[1052] ^ n[1053];
assign t[1054] = t[1053] ^ n[1054];
assign t[1055] = t[1054] ^ n[1055];
assign t[1056] = t[1055] ^ n[1056];
assign t[1057] = t[1056] ^ n[1057];
assign t[1058] = t[1057] ^ n[1058];
assign t[1059] = t[1058] ^ n[1059];
assign t[1060] = t[1059] ^ n[1060];
assign t[1061] = t[1060] ^ n[1061];
assign t[1062] = t[1061] ^ n[1062];
assign t[1063] = t[1062] ^ n[1063];
assign t[1064] = t[1063] ^ n[1064];
assign t[1065] = t[1064] ^ n[1065];
assign t[1066] = t[1065] ^ n[1066];
assign t[1067] = t[1066] ^ n[1067];
assign t[1068] = t[1067] ^ n[1068];
assign t[1069] = t[1068] ^ n[1069];
assign t[1070] = t[1069] ^ n[1070];
assign t[1071] = t[1070] ^ n[1071];
assign t[1072] = t[1071] ^ n[1072];
assign t[1073] = t[1072] ^ n[1073];
assign t[1074] = t[1073] ^ n[1074];
assign t[1075] = t[1074] ^ n[1075];
assign t[1076] = t[1075] ^ n[1076];
assign t[1077] = t[1076] ^ n[1077];
assign t[1078] = t[1077] ^ n[1078];
assign t[1079] = t[1078] ^ n[1079];
assign t[1080] = t[1079] ^ n[1080];
assign t[1081] = t[1080] ^ n[1081];
assign t[1082] = t[1081] ^ n[1082];
assign t[1083] = t[1082] ^ n[1083];
assign t[1084] = t[1083] ^ n[1084];
assign t[1085] = t[1084] ^ n[1085];
assign t[1086] = t[1085] ^ n[1086];
assign t[1087] = t[1086] ^ n[1087];
assign t[1088] = t[1087] ^ n[1088];
assign t[1089] = t[1088] ^ n[1089];
assign t[1090] = t[1089] ^ n[1090];
assign t[1091] = t[1090] ^ n[1091];
assign t[1092] = t[1091] ^ n[1092];
assign t[1093] = t[1092] ^ n[1093];
assign t[1094] = t[1093] ^ n[1094];
assign t[1095] = t[1094] ^ n[1095];
assign t[1096] = t[1095] ^ n[1096];
assign t[1097] = t[1096] ^ n[1097];
assign t[1098] = t[1097] ^ n[1098];
assign t[1099] = t[1098] ^ n[1099];
assign t[1100] = t[1099] ^ n[1100];
assign t[1101] = t[1100] ^ n[1101];
assign t[1102] = t[1101] ^ n[1102];
assign t[1103] = t[1102] ^ n[1103];
assign t[1104] = t[1103] ^ n[1104];
assign t[1105] = t[1104] ^ n[1105];
assign t[1106] = t[1105] ^ n[1106];
assign t[1107] = t[1106] ^ n[1107];
assign t[1108] = t[1107] ^ n[1108];
assign t[1109] = t[1108] ^ n[1109];
assign t[1110] = t[1109] ^ n[1110];
assign t[1111] = t[1110] ^ n[1111];
assign t[1112] = t[1111] ^ n[1112];
assign t[1113] = t[1112] ^ n[1113];
assign t[1114] = t[1113] ^ n[1114];
assign t[1115] = t[1114] ^ n[1115];
assign t[1116] = t[1115] ^ n[1116];
assign t[1117] = t[1116] ^ n[1117];
assign t[1118] = t[1117] ^ n[1118];
assign t[1119] = t[1118] ^ n[1119];
assign t[1120] = t[1119] ^ n[1120];
assign t[1121] = t[1120] ^ n[1121];
assign t[1122] = t[1121] ^ n[1122];
assign t[1123] = t[1122] ^ n[1123];
assign t[1124] = t[1123] ^ n[1124];
assign t[1125] = t[1124] ^ n[1125];
assign t[1126] = t[1125] ^ n[1126];
assign t[1127] = t[1126] ^ n[1127];
assign t[1128] = t[1127] ^ n[1128];
assign t[1129] = t[1128] ^ n[1129];
assign t[1130] = t[1129] ^ n[1130];
assign t[1131] = t[1130] ^ n[1131];
assign t[1132] = t[1131] ^ n[1132];
assign t[1133] = t[1132] ^ n[1133];
assign t[1134] = t[1133] ^ n[1134];
assign t[1135] = t[1134] ^ n[1135];
assign t[1136] = t[1135] ^ n[1136];
assign t[1137] = t[1136] ^ n[1137];
assign t[1138] = t[1137] ^ n[1138];
assign t[1139] = t[1138] ^ n[1139];
assign t[1140] = t[1139] ^ n[1140];
assign t[1141] = t[1140] ^ n[1141];
assign t[1142] = t[1141] ^ n[1142];
assign t[1143] = t[1142] ^ n[1143];
assign t[1144] = t[1143] ^ n[1144];
assign t[1145] = t[1144] ^ n[1145];
assign t[1146] = t[1145] ^ n[1146];
assign t[1147] = t[1146] ^ n[1147];
assign t[1148] = t[1147] ^ n[1148];
assign t[1149] = t[1148] ^ n[1149];
assign t[1150] = t[1149] ^ n[1150];
assign t[1151] = t[1150] ^ n[1151];
assign t[1152] = t[1151] ^ n[1152];
assign t[1153] = t[1152] ^ n[1153];
assign t[1154] = t[1153] ^ n[1154];
assign t[1155] = t[1154] ^ n[1155];
assign t[1156] = t[1155] ^ n[1156];
assign t[1157] = t[1156] ^ n[1157];
assign t[1158] = t[1157] ^ n[1158];
assign t[1159] = t[1158] ^ n[1159];
assign t[1160] = t[1159] ^ n[1160];
assign t[1161] = t[1160] ^ n[1161];
assign t[1162] = t[1161] ^ n[1162];
assign t[1163] = t[1162] ^ n[1163];
assign t[1164] = t[1163] ^ n[1164];
assign t[1165] = t[1164] ^ n[1165];
assign t[1166] = t[1165] ^ n[1166];
assign t[1167] = t[1166] ^ n[1167];
assign t[1168] = t[1167] ^ n[1168];
assign t[1169] = t[1168] ^ n[1169];
assign t[1170] = t[1169] ^ n[1170];
assign t[1171] = t[1170] ^ n[1171];
assign t[1172] = t[1171] ^ n[1172];
assign t[1173] = t[1172] ^ n[1173];
assign t[1174] = t[1173] ^ n[1174];
assign t[1175] = t[1174] ^ n[1175];
assign t[1176] = t[1175] ^ n[1176];
assign t[1177] = t[1176] ^ n[1177];
assign t[1178] = t[1177] ^ n[1178];
assign t[1179] = t[1178] ^ n[1179];
assign t[1180] = t[1179] ^ n[1180];
assign t[1181] = t[1180] ^ n[1181];
assign t[1182] = t[1181] ^ n[1182];
assign t[1183] = t[1182] ^ n[1183];
assign t[1184] = t[1183] ^ n[1184];
assign t[1185] = t[1184] ^ n[1185];
assign t[1186] = t[1185] ^ n[1186];
assign t[1187] = t[1186] ^ n[1187];
assign t[1188] = t[1187] ^ n[1188];
assign t[1189] = t[1188] ^ n[1189];
assign t[1190] = t[1189] ^ n[1190];
assign t[1191] = t[1190] ^ n[1191];
assign t[1192] = t[1191] ^ n[1192];
assign t[1193] = t[1192] ^ n[1193];
assign t[1194] = t[1193] ^ n[1194];
assign t[1195] = t[1194] ^ n[1195];
assign t[1196] = t[1195] ^ n[1196];
assign t[1197] = t[1196] ^ n[1197];
assign t[1198] = t[1197] ^ n[1198];
assign t[1199] = t[1198] ^ n[1199];
assign t[1200] = t[1199] ^ n[1200];
assign t[1201] = t[1200] ^ n[1201];
assign t[1202] = t[1201] ^ n[1202];
assign t[1203] = t[1202] ^ n[1203];
assign t[1204] = t[1203] ^ n[1204];
assign t[1205] = t[1204] ^ n[1205];
assign t[1206] = t[1205] ^ n[1206];
assign t[1207] = t[1206] ^ n[1207];
assign t[1208] = t[1207] ^ n[1208];
assign t[1209] = t[1208] ^ n[1209];
assign t[1210] = t[1209] ^ n[1210];
assign t[1211] = t[1210] ^ n[1211];
assign t[1212] = t[1211] ^ n[1212];
assign t[1213] = t[1212] ^ n[1213];
assign t[1214] = t[1213] ^ n[1214];
assign t[1215] = t[1214] ^ n[1215];
assign t[1216] = t[1215] ^ n[1216];
assign t[1217] = t[1216] ^ n[1217];
assign t[1218] = t[1217] ^ n[1218];
assign t[1219] = t[1218] ^ n[1219];
assign t[1220] = t[1219] ^ n[1220];
assign t[1221] = t[1220] ^ n[1221];
assign t[1222] = t[1221] ^ n[1222];
assign t[1223] = t[1222] ^ n[1223];
assign t[1224] = t[1223] ^ n[1224];
assign t[1225] = t[1224] ^ n[1225];
assign t[1226] = t[1225] ^ n[1226];
assign t[1227] = t[1226] ^ n[1227];
assign t[1228] = t[1227] ^ n[1228];
assign t[1229] = t[1228] ^ n[1229];
assign t[1230] = t[1229] ^ n[1230];
assign t[1231] = t[1230] ^ n[1231];
assign t[1232] = t[1231] ^ n[1232];
assign t[1233] = t[1232] ^ n[1233];
assign t[1234] = t[1233] ^ n[1234];
assign t[1235] = t[1234] ^ n[1235];
assign t[1236] = t[1235] ^ n[1236];
assign t[1237] = t[1236] ^ n[1237];
assign t[1238] = t[1237] ^ n[1238];
assign t[1239] = t[1238] ^ n[1239];
assign t[1240] = t[1239] ^ n[1240];
assign t[1241] = t[1240] ^ n[1241];
assign t[1242] = t[1241] ^ n[1242];
assign t[1243] = t[1242] ^ n[1243];
assign t[1244] = t[1243] ^ n[1244];
assign t[1245] = t[1244] ^ n[1245];
assign t[1246] = t[1245] ^ n[1246];
assign t[1247] = t[1246] ^ n[1247];
assign t[1248] = t[1247] ^ n[1248];
assign t[1249] = t[1248] ^ n[1249];
assign t[1250] = t[1249] ^ n[1250];
assign t[1251] = t[1250] ^ n[1251];
assign t[1252] = t[1251] ^ n[1252];
assign t[1253] = t[1252] ^ n[1253];
assign t[1254] = t[1253] ^ n[1254];
assign t[1255] = t[1254] ^ n[1255];
assign t[1256] = t[1255] ^ n[1256];
assign t[1257] = t[1256] ^ n[1257];
assign t[1258] = t[1257] ^ n[1258];
assign t[1259] = t[1258] ^ n[1259];
assign t[1260] = t[1259] ^ n[1260];
assign t[1261] = t[1260] ^ n[1261];
assign t[1262] = t[1261] ^ n[1262];
assign t[1263] = t[1262] ^ n[1263];
assign t[1264] = t[1263] ^ n[1264];
assign t[1265] = t[1264] ^ n[1265];
assign t[1266] = t[1265] ^ n[1266];
assign t[1267] = t[1266] ^ n[1267];
assign t[1268] = t[1267] ^ n[1268];
assign t[1269] = t[1268] ^ n[1269];
assign t[1270] = t[1269] ^ n[1270];
assign t[1271] = t[1270] ^ n[1271];
assign t[1272] = t[1271] ^ n[1272];
assign t[1273] = t[1272] ^ n[1273];
assign t[1274] = t[1273] ^ n[1274];
assign t[1275] = t[1274] ^ n[1275];
assign t[1276] = t[1275] ^ n[1276];
assign t[1277] = t[1276] ^ n[1277];
assign t[1278] = t[1277] ^ n[1278];
assign t[1279] = t[1278] ^ n[1279];
assign t[1280] = t[1279] ^ n[1280];
assign t[1281] = t[1280] ^ n[1281];
assign t[1282] = t[1281] ^ n[1282];
assign t[1283] = t[1282] ^ n[1283];
assign t[1284] = t[1283] ^ n[1284];
assign t[1285] = t[1284] ^ n[1285];
assign t[1286] = t[1285] ^ n[1286];
assign t[1287] = t[1286] ^ n[1287];
assign t[1288] = t[1287] ^ n[1288];
assign t[1289] = t[1288] ^ n[1289];
assign t[1290] = t[1289] ^ n[1290];
assign t[1291] = t[1290] ^ n[1291];
assign t[1292] = t[1291] ^ n[1292];
assign t[1293] = t[1292] ^ n[1293];
assign t[1294] = t[1293] ^ n[1294];
assign t[1295] = t[1294] ^ n[1295];
assign t[1296] = t[1295] ^ n[1296];
assign t[1297] = t[1296] ^ n[1297];
assign t[1298] = t[1297] ^ n[1298];
assign t[1299] = t[1298] ^ n[1299];
assign t[1300] = t[1299] ^ n[1300];
assign t[1301] = t[1300] ^ n[1301];
assign t[1302] = t[1301] ^ n[1302];
assign t[1303] = t[1302] ^ n[1303];
assign t[1304] = t[1303] ^ n[1304];
assign t[1305] = t[1304] ^ n[1305];
assign t[1306] = t[1305] ^ n[1306];
assign t[1307] = t[1306] ^ n[1307];
assign t[1308] = t[1307] ^ n[1308];
assign t[1309] = t[1308] ^ n[1309];
assign t[1310] = t[1309] ^ n[1310];
assign t[1311] = t[1310] ^ n[1311];
assign t[1312] = t[1311] ^ n[1312];
assign t[1313] = t[1312] ^ n[1313];
assign t[1314] = t[1313] ^ n[1314];
assign t[1315] = t[1314] ^ n[1315];
assign t[1316] = t[1315] ^ n[1316];
assign t[1317] = t[1316] ^ n[1317];
assign t[1318] = t[1317] ^ n[1318];
assign t[1319] = t[1318] ^ n[1319];
assign t[1320] = t[1319] ^ n[1320];
assign t[1321] = t[1320] ^ n[1321];
assign t[1322] = t[1321] ^ n[1322];
assign t[1323] = t[1322] ^ n[1323];
assign t[1324] = t[1323] ^ n[1324];
assign t[1325] = t[1324] ^ n[1325];
assign t[1326] = t[1325] ^ n[1326];
assign t[1327] = t[1326] ^ n[1327];
assign t[1328] = t[1327] ^ n[1328];
assign t[1329] = t[1328] ^ n[1329];
assign t[1330] = t[1329] ^ n[1330];
assign t[1331] = t[1330] ^ n[1331];
assign t[1332] = t[1331] ^ n[1332];
assign t[1333] = t[1332] ^ n[1333];
assign t[1334] = t[1333] ^ n[1334];
assign t[1335] = t[1334] ^ n[1335];
assign t[1336] = t[1335] ^ n[1336];
assign t[1337] = t[1336] ^ n[1337];
assign t[1338] = t[1337] ^ n[1338];
assign t[1339] = t[1338] ^ n[1339];
assign t[1340] = t[1339] ^ n[1340];
assign t[1341] = t[1340] ^ n[1341];
assign t[1342] = t[1341] ^ n[1342];
assign t[1343] = t[1342] ^ n[1343];
assign t[1344] = t[1343] ^ n[1344];
assign t[1345] = t[1344] ^ n[1345];
assign t[1346] = t[1345] ^ n[1346];
assign t[1347] = t[1346] ^ n[1347];
assign t[1348] = t[1347] ^ n[1348];
assign t[1349] = t[1348] ^ n[1349];
assign t[1350] = t[1349] ^ n[1350];
assign t[1351] = t[1350] ^ n[1351];
assign t[1352] = t[1351] ^ n[1352];
assign t[1353] = t[1352] ^ n[1353];
assign t[1354] = t[1353] ^ n[1354];
assign t[1355] = t[1354] ^ n[1355];
assign t[1356] = t[1355] ^ n[1356];
assign t[1357] = t[1356] ^ n[1357];
assign t[1358] = t[1357] ^ n[1358];
assign t[1359] = t[1358] ^ n[1359];
assign t[1360] = t[1359] ^ n[1360];
assign t[1361] = t[1360] ^ n[1361];
assign t[1362] = t[1361] ^ n[1362];
assign t[1363] = t[1362] ^ n[1363];
assign t[1364] = t[1363] ^ n[1364];
assign t[1365] = t[1364] ^ n[1365];
assign t[1366] = t[1365] ^ n[1366];
assign t[1367] = t[1366] ^ n[1367];
assign t[1368] = t[1367] ^ n[1368];
assign t[1369] = t[1368] ^ n[1369];
assign t[1370] = t[1369] ^ n[1370];
assign t[1371] = t[1370] ^ n[1371];
assign t[1372] = t[1371] ^ n[1372];
assign t[1373] = t[1372] ^ n[1373];
assign t[1374] = t[1373] ^ n[1374];
assign t[1375] = t[1374] ^ n[1375];
assign t[1376] = t[1375] ^ n[1376];
assign t[1377] = t[1376] ^ n[1377];
assign t[1378] = t[1377] ^ n[1378];
assign t[1379] = t[1378] ^ n[1379];
assign t[1380] = t[1379] ^ n[1380];
assign t[1381] = t[1380] ^ n[1381];
assign t[1382] = t[1381] ^ n[1382];
assign t[1383] = t[1382] ^ n[1383];
assign t[1384] = t[1383] ^ n[1384];
assign t[1385] = t[1384] ^ n[1385];
assign t[1386] = t[1385] ^ n[1386];
assign t[1387] = t[1386] ^ n[1387];
assign t[1388] = t[1387] ^ n[1388];
assign t[1389] = t[1388] ^ n[1389];
assign t[1390] = t[1389] ^ n[1390];
assign t[1391] = t[1390] ^ n[1391];
assign t[1392] = t[1391] ^ n[1392];
assign t[1393] = t[1392] ^ n[1393];
assign t[1394] = t[1393] ^ n[1394];
assign t[1395] = t[1394] ^ n[1395];
assign t[1396] = t[1395] ^ n[1396];
assign t[1397] = t[1396] ^ n[1397];
assign t[1398] = t[1397] ^ n[1398];
assign t[1399] = t[1398] ^ n[1399];
assign t[1400] = t[1399] ^ n[1400];
assign t[1401] = t[1400] ^ n[1401];
assign t[1402] = t[1401] ^ n[1402];
assign t[1403] = t[1402] ^ n[1403];
assign t[1404] = t[1403] ^ n[1404];
assign t[1405] = t[1404] ^ n[1405];
assign t[1406] = t[1405] ^ n[1406];
assign t[1407] = t[1406] ^ n[1407];
assign t[1408] = t[1407] ^ n[1408];
assign t[1409] = t[1408] ^ n[1409];
assign t[1410] = t[1409] ^ n[1410];
assign t[1411] = t[1410] ^ n[1411];
assign t[1412] = t[1411] ^ n[1412];
assign t[1413] = t[1412] ^ n[1413];
assign t[1414] = t[1413] ^ n[1414];
assign t[1415] = t[1414] ^ n[1415];
assign t[1416] = t[1415] ^ n[1416];
assign t[1417] = t[1416] ^ n[1417];
assign t[1418] = t[1417] ^ n[1418];
assign t[1419] = t[1418] ^ n[1419];
assign t[1420] = t[1419] ^ n[1420];
assign t[1421] = t[1420] ^ n[1421];
assign t[1422] = t[1421] ^ n[1422];
assign t[1423] = t[1422] ^ n[1423];
assign t[1424] = t[1423] ^ n[1424];
assign t[1425] = t[1424] ^ n[1425];
assign t[1426] = t[1425] ^ n[1426];
assign t[1427] = t[1426] ^ n[1427];
assign t[1428] = t[1427] ^ n[1428];
assign t[1429] = t[1428] ^ n[1429];
assign t[1430] = t[1429] ^ n[1430];
assign t[1431] = t[1430] ^ n[1431];
assign t[1432] = t[1431] ^ n[1432];
assign t[1433] = t[1432] ^ n[1433];
assign t[1434] = t[1433] ^ n[1434];
assign t[1435] = t[1434] ^ n[1435];
assign t[1436] = t[1435] ^ n[1436];
assign t[1437] = t[1436] ^ n[1437];
assign t[1438] = t[1437] ^ n[1438];
assign t[1439] = t[1438] ^ n[1439];
assign t[1440] = t[1439] ^ n[1440];
assign t[1441] = t[1440] ^ n[1441];
assign t[1442] = t[1441] ^ n[1442];
assign t[1443] = t[1442] ^ n[1443];
assign t[1444] = t[1443] ^ n[1444];
assign t[1445] = t[1444] ^ n[1445];
assign t[1446] = t[1445] ^ n[1446];
assign t[1447] = t[1446] ^ n[1447];
assign t[1448] = t[1447] ^ n[1448];
assign t[1449] = t[1448] ^ n[1449];
assign t[1450] = t[1449] ^ n[1450];
assign t[1451] = t[1450] ^ n[1451];
assign t[1452] = t[1451] ^ n[1452];
assign t[1453] = t[1452] ^ n[1453];
assign t[1454] = t[1453] ^ n[1454];
assign t[1455] = t[1454] ^ n[1455];
assign t[1456] = t[1455] ^ n[1456];
assign t[1457] = t[1456] ^ n[1457];
assign t[1458] = t[1457] ^ n[1458];
assign t[1459] = t[1458] ^ n[1459];
assign t[1460] = t[1459] ^ n[1460];
assign t[1461] = t[1460] ^ n[1461];
assign t[1462] = t[1461] ^ n[1462];
assign t[1463] = t[1462] ^ n[1463];
assign t[1464] = t[1463] ^ n[1464];
assign t[1465] = t[1464] ^ n[1465];
assign t[1466] = t[1465] ^ n[1466];
assign t[1467] = t[1466] ^ n[1467];
assign t[1468] = t[1467] ^ n[1468];
assign t[1469] = t[1468] ^ n[1469];
assign t[1470] = t[1469] ^ n[1470];
assign t[1471] = t[1470] ^ n[1471];
assign t[1472] = t[1471] ^ n[1472];
assign t[1473] = t[1472] ^ n[1473];
assign t[1474] = t[1473] ^ n[1474];
assign t[1475] = t[1474] ^ n[1475];
assign t[1476] = t[1475] ^ n[1476];
assign t[1477] = t[1476] ^ n[1477];
assign t[1478] = t[1477] ^ n[1478];
assign t[1479] = t[1478] ^ n[1479];
assign t[1480] = t[1479] ^ n[1480];
assign t[1481] = t[1480] ^ n[1481];
assign t[1482] = t[1481] ^ n[1482];
assign t[1483] = t[1482] ^ n[1483];
assign t[1484] = t[1483] ^ n[1484];
assign t[1485] = t[1484] ^ n[1485];
assign t[1486] = t[1485] ^ n[1486];
assign t[1487] = t[1486] ^ n[1487];
assign t[1488] = t[1487] ^ n[1488];
assign t[1489] = t[1488] ^ n[1489];
assign t[1490] = t[1489] ^ n[1490];
assign t[1491] = t[1490] ^ n[1491];
assign t[1492] = t[1491] ^ n[1492];
assign t[1493] = t[1492] ^ n[1493];
assign t[1494] = t[1493] ^ n[1494];
assign t[1495] = t[1494] ^ n[1495];
assign t[1496] = t[1495] ^ n[1496];
assign t[1497] = t[1496] ^ n[1497];
assign t[1498] = t[1497] ^ n[1498];
assign t[1499] = t[1498] ^ n[1499];
assign t[1500] = t[1499] ^ n[1500];
assign t[1501] = t[1500] ^ n[1501];
assign t[1502] = t[1501] ^ n[1502];
assign t[1503] = t[1502] ^ n[1503];
assign t[1504] = t[1503] ^ n[1504];
assign t[1505] = t[1504] ^ n[1505];
assign t[1506] = t[1505] ^ n[1506];
assign t[1507] = t[1506] ^ n[1507];
assign t[1508] = t[1507] ^ n[1508];
assign t[1509] = t[1508] ^ n[1509];
assign t[1510] = t[1509] ^ n[1510];
assign t[1511] = t[1510] ^ n[1511];
assign t[1512] = t[1511] ^ n[1512];
assign t[1513] = t[1512] ^ n[1513];
assign t[1514] = t[1513] ^ n[1514];
assign t[1515] = t[1514] ^ n[1515];
assign t[1516] = t[1515] ^ n[1516];
assign t[1517] = t[1516] ^ n[1517];
assign t[1518] = t[1517] ^ n[1518];
assign t[1519] = t[1518] ^ n[1519];
assign t[1520] = t[1519] ^ n[1520];
assign t[1521] = t[1520] ^ n[1521];
assign t[1522] = t[1521] ^ n[1522];
assign t[1523] = t[1522] ^ n[1523];
assign t[1524] = t[1523] ^ n[1524];
assign t[1525] = t[1524] ^ n[1525];
assign t[1526] = t[1525] ^ n[1526];
assign t[1527] = t[1526] ^ n[1527];
assign t[1528] = t[1527] ^ n[1528];
assign t[1529] = t[1528] ^ n[1529];
assign t[1530] = t[1529] ^ n[1530];
assign t[1531] = t[1530] ^ n[1531];
assign t[1532] = t[1531] ^ n[1532];
assign t[1533] = t[1532] ^ n[1533];
assign t[1534] = t[1533] ^ n[1534];
assign t[1535] = t[1534] ^ n[1535];
assign t[1536] = t[1535] ^ n[1536];
assign t[1537] = t[1536] ^ n[1537];
assign t[1538] = t[1537] ^ n[1538];
assign t[1539] = t[1538] ^ n[1539];
assign t[1540] = t[1539] ^ n[1540];
assign t[1541] = t[1540] ^ n[1541];
assign t[1542] = t[1541] ^ n[1542];
assign t[1543] = t[1542] ^ n[1543];
assign t[1544] = t[1543] ^ n[1544];
assign t[1545] = t[1544] ^ n[1545];
assign t[1546] = t[1545] ^ n[1546];
assign t[1547] = t[1546] ^ n[1547];
assign t[1548] = t[1547] ^ n[1548];
assign t[1549] = t[1548] ^ n[1549];
assign t[1550] = t[1549] ^ n[1550];
assign t[1551] = t[1550] ^ n[1551];
assign t[1552] = t[1551] ^ n[1552];
assign t[1553] = t[1552] ^ n[1553];
assign t[1554] = t[1553] ^ n[1554];
assign t[1555] = t[1554] ^ n[1555];
assign t[1556] = t[1555] ^ n[1556];
assign t[1557] = t[1556] ^ n[1557];
assign t[1558] = t[1557] ^ n[1558];
assign t[1559] = t[1558] ^ n[1559];
assign t[1560] = t[1559] ^ n[1560];
assign t[1561] = t[1560] ^ n[1561];
assign t[1562] = t[1561] ^ n[1562];
assign t[1563] = t[1562] ^ n[1563];
assign t[1564] = t[1563] ^ n[1564];
assign t[1565] = t[1564] ^ n[1565];
assign t[1566] = t[1565] ^ n[1566];
assign t[1567] = t[1566] ^ n[1567];
assign t[1568] = t[1567] ^ n[1568];
assign t[1569] = t[1568] ^ n[1569];
assign t[1570] = t[1569] ^ n[1570];
assign t[1571] = t[1570] ^ n[1571];
assign t[1572] = t[1571] ^ n[1572];
assign t[1573] = t[1572] ^ n[1573];
assign t[1574] = t[1573] ^ n[1574];
assign t[1575] = t[1574] ^ n[1575];
assign t[1576] = t[1575] ^ n[1576];
assign t[1577] = t[1576] ^ n[1577];
assign t[1578] = t[1577] ^ n[1578];
assign t[1579] = t[1578] ^ n[1579];
assign t[1580] = t[1579] ^ n[1580];
assign t[1581] = t[1580] ^ n[1581];
assign t[1582] = t[1581] ^ n[1582];
assign t[1583] = t[1582] ^ n[1583];
assign t[1584] = t[1583] ^ n[1584];
assign t[1585] = t[1584] ^ n[1585];
assign t[1586] = t[1585] ^ n[1586];
assign t[1587] = t[1586] ^ n[1587];
assign t[1588] = t[1587] ^ n[1588];
assign t[1589] = t[1588] ^ n[1589];
assign t[1590] = t[1589] ^ n[1590];
assign t[1591] = t[1590] ^ n[1591];
assign t[1592] = t[1591] ^ n[1592];
assign t[1593] = t[1592] ^ n[1593];
assign t[1594] = t[1593] ^ n[1594];
assign t[1595] = t[1594] ^ n[1595];
assign t[1596] = t[1595] ^ n[1596];
assign t[1597] = t[1596] ^ n[1597];
assign t[1598] = t[1597] ^ n[1598];
assign t[1599] = t[1598] ^ n[1599];
assign t[1600] = t[1599] ^ n[1600];
assign t[1601] = t[1600] ^ n[1601];
assign t[1602] = t[1601] ^ n[1602];
assign t[1603] = t[1602] ^ n[1603];
assign t[1604] = t[1603] ^ n[1604];
assign t[1605] = t[1604] ^ n[1605];
assign t[1606] = t[1605] ^ n[1606];
assign t[1607] = t[1606] ^ n[1607];
assign t[1608] = t[1607] ^ n[1608];
assign t[1609] = t[1608] ^ n[1609];
assign t[1610] = t[1609] ^ n[1610];
assign t[1611] = t[1610] ^ n[1611];
assign t[1612] = t[1611] ^ n[1612];
assign t[1613] = t[1612] ^ n[1613];
assign t[1614] = t[1613] ^ n[1614];
assign t[1615] = t[1614] ^ n[1615];
assign t[1616] = t[1615] ^ n[1616];
assign t[1617] = t[1616] ^ n[1617];
assign t[1618] = t[1617] ^ n[1618];
assign t[1619] = t[1618] ^ n[1619];
assign t[1620] = t[1619] ^ n[1620];
assign t[1621] = t[1620] ^ n[1621];
assign t[1622] = t[1621] ^ n[1622];
assign t[1623] = t[1622] ^ n[1623];
assign t[1624] = t[1623] ^ n[1624];
assign t[1625] = t[1624] ^ n[1625];
assign t[1626] = t[1625] ^ n[1626];
assign t[1627] = t[1626] ^ n[1627];
assign t[1628] = t[1627] ^ n[1628];
assign t[1629] = t[1628] ^ n[1629];
assign t[1630] = t[1629] ^ n[1630];
assign t[1631] = t[1630] ^ n[1631];
assign t[1632] = t[1631] ^ n[1632];
assign t[1633] = t[1632] ^ n[1633];
assign t[1634] = t[1633] ^ n[1634];
assign t[1635] = t[1634] ^ n[1635];
assign t[1636] = t[1635] ^ n[1636];
assign t[1637] = t[1636] ^ n[1637];
assign t[1638] = t[1637] ^ n[1638];
assign t[1639] = t[1638] ^ n[1639];
assign t[1640] = t[1639] ^ n[1640];
assign t[1641] = t[1640] ^ n[1641];
assign t[1642] = t[1641] ^ n[1642];
assign t[1643] = t[1642] ^ n[1643];
assign t[1644] = t[1643] ^ n[1644];
assign t[1645] = t[1644] ^ n[1645];
assign t[1646] = t[1645] ^ n[1646];
assign t[1647] = t[1646] ^ n[1647];
assign t[1648] = t[1647] ^ n[1648];
assign t[1649] = t[1648] ^ n[1649];
assign t[1650] = t[1649] ^ n[1650];
assign t[1651] = t[1650] ^ n[1651];
assign t[1652] = t[1651] ^ n[1652];
assign t[1653] = t[1652] ^ n[1653];
assign t[1654] = t[1653] ^ n[1654];
assign t[1655] = t[1654] ^ n[1655];
assign t[1656] = t[1655] ^ n[1656];
assign t[1657] = t[1656] ^ n[1657];
assign t[1658] = t[1657] ^ n[1658];
assign t[1659] = t[1658] ^ n[1659];
assign t[1660] = t[1659] ^ n[1660];
assign t[1661] = t[1660] ^ n[1661];
assign t[1662] = t[1661] ^ n[1662];
assign t[1663] = t[1662] ^ n[1663];
assign t[1664] = t[1663] ^ n[1664];
assign t[1665] = t[1664] ^ n[1665];
assign t[1666] = t[1665] ^ n[1666];
assign t[1667] = t[1666] ^ n[1667];
assign t[1668] = t[1667] ^ n[1668];
assign t[1669] = t[1668] ^ n[1669];
assign t[1670] = t[1669] ^ n[1670];
assign t[1671] = t[1670] ^ n[1671];
assign t[1672] = t[1671] ^ n[1672];
assign t[1673] = t[1672] ^ n[1673];
assign t[1674] = t[1673] ^ n[1674];
assign t[1675] = t[1674] ^ n[1675];
assign t[1676] = t[1675] ^ n[1676];
assign t[1677] = t[1676] ^ n[1677];
assign t[1678] = t[1677] ^ n[1678];
assign t[1679] = t[1678] ^ n[1679];
assign t[1680] = t[1679] ^ n[1680];
assign t[1681] = t[1680] ^ n[1681];
assign t[1682] = t[1681] ^ n[1682];
assign t[1683] = t[1682] ^ n[1683];
assign t[1684] = t[1683] ^ n[1684];
assign t[1685] = t[1684] ^ n[1685];
assign t[1686] = t[1685] ^ n[1686];
assign t[1687] = t[1686] ^ n[1687];
assign t[1688] = t[1687] ^ n[1688];
assign t[1689] = t[1688] ^ n[1689];
assign t[1690] = t[1689] ^ n[1690];
assign t[1691] = t[1690] ^ n[1691];
assign t[1692] = t[1691] ^ n[1692];
assign t[1693] = t[1692] ^ n[1693];
assign t[1694] = t[1693] ^ n[1694];
assign t[1695] = t[1694] ^ n[1695];
assign t[1696] = t[1695] ^ n[1696];
assign t[1697] = t[1696] ^ n[1697];
assign t[1698] = t[1697] ^ n[1698];
assign t[1699] = t[1698] ^ n[1699];
assign t[1700] = t[1699] ^ n[1700];
assign t[1701] = t[1700] ^ n[1701];
assign t[1702] = t[1701] ^ n[1702];
assign t[1703] = t[1702] ^ n[1703];
assign t[1704] = t[1703] ^ n[1704];
assign t[1705] = t[1704] ^ n[1705];
assign t[1706] = t[1705] ^ n[1706];
assign t[1707] = t[1706] ^ n[1707];
assign t[1708] = t[1707] ^ n[1708];
assign t[1709] = t[1708] ^ n[1709];
assign t[1710] = t[1709] ^ n[1710];
assign t[1711] = t[1710] ^ n[1711];
assign t[1712] = t[1711] ^ n[1712];
assign t[1713] = t[1712] ^ n[1713];
assign t[1714] = t[1713] ^ n[1714];
assign t[1715] = t[1714] ^ n[1715];
assign t[1716] = t[1715] ^ n[1716];
assign t[1717] = t[1716] ^ n[1717];
assign t[1718] = t[1717] ^ n[1718];
assign t[1719] = t[1718] ^ n[1719];
assign t[1720] = t[1719] ^ n[1720];
assign t[1721] = t[1720] ^ n[1721];
assign t[1722] = t[1721] ^ n[1722];
assign t[1723] = t[1722] ^ n[1723];
assign t[1724] = t[1723] ^ n[1724];
assign t[1725] = t[1724] ^ n[1725];
assign t[1726] = t[1725] ^ n[1726];
assign t[1727] = t[1726] ^ n[1727];
assign t[1728] = t[1727] ^ n[1728];
assign t[1729] = t[1728] ^ n[1729];
assign t[1730] = t[1729] ^ n[1730];
assign t[1731] = t[1730] ^ n[1731];
assign t[1732] = t[1731] ^ n[1732];
assign t[1733] = t[1732] ^ n[1733];
assign t[1734] = t[1733] ^ n[1734];
assign t[1735] = t[1734] ^ n[1735];
assign t[1736] = t[1735] ^ n[1736];
assign t[1737] = t[1736] ^ n[1737];
assign t[1738] = t[1737] ^ n[1738];
assign t[1739] = t[1738] ^ n[1739];
assign t[1740] = t[1739] ^ n[1740];
assign t[1741] = t[1740] ^ n[1741];
assign t[1742] = t[1741] ^ n[1742];
assign t[1743] = t[1742] ^ n[1743];
assign t[1744] = t[1743] ^ n[1744];
assign t[1745] = t[1744] ^ n[1745];
assign t[1746] = t[1745] ^ n[1746];
assign t[1747] = t[1746] ^ n[1747];
assign t[1748] = t[1747] ^ n[1748];
assign t[1749] = t[1748] ^ n[1749];
assign t[1750] = t[1749] ^ n[1750];
assign t[1751] = t[1750] ^ n[1751];
assign t[1752] = t[1751] ^ n[1752];
assign t[1753] = t[1752] ^ n[1753];
assign t[1754] = t[1753] ^ n[1754];
assign t[1755] = t[1754] ^ n[1755];
assign t[1756] = t[1755] ^ n[1756];
assign t[1757] = t[1756] ^ n[1757];
assign t[1758] = t[1757] ^ n[1758];
assign t[1759] = t[1758] ^ n[1759];
assign t[1760] = t[1759] ^ n[1760];
assign t[1761] = t[1760] ^ n[1761];
assign t[1762] = t[1761] ^ n[1762];
assign t[1763] = t[1762] ^ n[1763];
assign t[1764] = t[1763] ^ n[1764];
assign t[1765] = t[1764] ^ n[1765];
assign t[1766] = t[1765] ^ n[1766];
assign t[1767] = t[1766] ^ n[1767];
assign t[1768] = t[1767] ^ n[1768];
assign t[1769] = t[1768] ^ n[1769];
assign t[1770] = t[1769] ^ n[1770];
assign t[1771] = t[1770] ^ n[1771];
assign t[1772] = t[1771] ^ n[1772];
assign t[1773] = t[1772] ^ n[1773];
assign t[1774] = t[1773] ^ n[1774];
assign t[1775] = t[1774] ^ n[1775];
assign t[1776] = t[1775] ^ n[1776];
assign t[1777] = t[1776] ^ n[1777];
assign t[1778] = t[1777] ^ n[1778];
assign t[1779] = t[1778] ^ n[1779];
assign t[1780] = t[1779] ^ n[1780];
assign t[1781] = t[1780] ^ n[1781];
assign t[1782] = t[1781] ^ n[1782];
assign t[1783] = t[1782] ^ n[1783];
assign t[1784] = t[1783] ^ n[1784];
assign t[1785] = t[1784] ^ n[1785];
assign t[1786] = t[1785] ^ n[1786];
assign t[1787] = t[1786] ^ n[1787];
assign t[1788] = t[1787] ^ n[1788];
assign t[1789] = t[1788] ^ n[1789];
assign t[1790] = t[1789] ^ n[1790];
assign t[1791] = t[1790] ^ n[1791];
assign t[1792] = t[1791] ^ n[1792];
assign t[1793] = t[1792] ^ n[1793];
assign t[1794] = t[1793] ^ n[1794];
assign t[1795] = t[1794] ^ n[1795];
assign t[1796] = t[1795] ^ n[1796];
assign t[1797] = t[1796] ^ n[1797];
assign t[1798] = t[1797] ^ n[1798];
assign t[1799] = t[1798] ^ n[1799];
assign t[1800] = t[1799] ^ n[1800];
assign t[1801] = t[1800] ^ n[1801];
assign t[1802] = t[1801] ^ n[1802];
assign t[1803] = t[1802] ^ n[1803];
assign t[1804] = t[1803] ^ n[1804];
assign t[1805] = t[1804] ^ n[1805];
assign t[1806] = t[1805] ^ n[1806];
assign t[1807] = t[1806] ^ n[1807];
assign t[1808] = t[1807] ^ n[1808];
assign t[1809] = t[1808] ^ n[1809];
assign t[1810] = t[1809] ^ n[1810];
assign t[1811] = t[1810] ^ n[1811];
assign t[1812] = t[1811] ^ n[1812];
assign t[1813] = t[1812] ^ n[1813];
assign t[1814] = t[1813] ^ n[1814];
assign t[1815] = t[1814] ^ n[1815];
assign t[1816] = t[1815] ^ n[1816];
assign t[1817] = t[1816] ^ n[1817];
assign t[1818] = t[1817] ^ n[1818];
assign t[1819] = t[1818] ^ n[1819];
assign t[1820] = t[1819] ^ n[1820];
assign t[1821] = t[1820] ^ n[1821];
assign t[1822] = t[1821] ^ n[1822];
assign t[1823] = t[1822] ^ n[1823];
assign t[1824] = t[1823] ^ n[1824];
assign t[1825] = t[1824] ^ n[1825];
assign t[1826] = t[1825] ^ n[1826];
assign t[1827] = t[1826] ^ n[1827];
assign t[1828] = t[1827] ^ n[1828];
assign t[1829] = t[1828] ^ n[1829];
assign t[1830] = t[1829] ^ n[1830];
assign t[1831] = t[1830] ^ n[1831];
assign t[1832] = t[1831] ^ n[1832];
assign t[1833] = t[1832] ^ n[1833];
assign t[1834] = t[1833] ^ n[1834];
assign t[1835] = t[1834] ^ n[1835];
assign t[1836] = t[1835] ^ n[1836];
assign t[1837] = t[1836] ^ n[1837];
assign t[1838] = t[1837] ^ n[1838];
assign t[1839] = t[1838] ^ n[1839];
assign t[1840] = t[1839] ^ n[1840];
assign t[1841] = t[1840] ^ n[1841];
assign t[1842] = t[1841] ^ n[1842];
assign t[1843] = t[1842] ^ n[1843];
assign t[1844] = t[1843] ^ n[1844];
assign t[1845] = t[1844] ^ n[1845];
assign t[1846] = t[1845] ^ n[1846];
assign t[1847] = t[1846] ^ n[1847];
assign t[1848] = t[1847] ^ n[1848];
assign t[1849] = t[1848] ^ n[1849];
assign t[1850] = t[1849] ^ n[1850];
assign t[1851] = t[1850] ^ n[1851];
assign t[1852] = t[1851] ^ n[1852];
assign t[1853] = t[1852] ^ n[1853];
assign t[1854] = t[1853] ^ n[1854];
assign t[1855] = t[1854] ^ n[1855];
assign t[1856] = t[1855] ^ n[1856];
assign t[1857] = t[1856] ^ n[1857];
assign t[1858] = t[1857] ^ n[1858];
assign t[1859] = t[1858] ^ n[1859];
assign t[1860] = t[1859] ^ n[1860];
assign t[1861] = t[1860] ^ n[1861];
assign t[1862] = t[1861] ^ n[1862];
assign t[1863] = t[1862] ^ n[1863];
assign t[1864] = t[1863] ^ n[1864];
assign t[1865] = t[1864] ^ n[1865];
assign t[1866] = t[1865] ^ n[1866];
assign t[1867] = t[1866] ^ n[1867];
assign t[1868] = t[1867] ^ n[1868];
assign t[1869] = t[1868] ^ n[1869];
assign t[1870] = t[1869] ^ n[1870];
assign t[1871] = t[1870] ^ n[1871];
assign t[1872] = t[1871] ^ n[1872];
assign t[1873] = t[1872] ^ n[1873];
assign t[1874] = t[1873] ^ n[1874];
assign t[1875] = t[1874] ^ n[1875];
assign t[1876] = t[1875] ^ n[1876];
assign t[1877] = t[1876] ^ n[1877];
assign t[1878] = t[1877] ^ n[1878];
assign t[1879] = t[1878] ^ n[1879];
assign t[1880] = t[1879] ^ n[1880];
assign t[1881] = t[1880] ^ n[1881];
assign t[1882] = t[1881] ^ n[1882];
assign t[1883] = t[1882] ^ n[1883];
assign t[1884] = t[1883] ^ n[1884];
assign t[1885] = t[1884] ^ n[1885];
assign t[1886] = t[1885] ^ n[1886];
assign t[1887] = t[1886] ^ n[1887];
assign t[1888] = t[1887] ^ n[1888];
assign t[1889] = t[1888] ^ n[1889];
assign t[1890] = t[1889] ^ n[1890];
assign t[1891] = t[1890] ^ n[1891];
assign t[1892] = t[1891] ^ n[1892];
assign t[1893] = t[1892] ^ n[1893];
assign t[1894] = t[1893] ^ n[1894];
assign t[1895] = t[1894] ^ n[1895];
assign t[1896] = t[1895] ^ n[1896];
assign t[1897] = t[1896] ^ n[1897];
assign t[1898] = t[1897] ^ n[1898];
assign t[1899] = t[1898] ^ n[1899];
assign t[1900] = t[1899] ^ n[1900];
assign t[1901] = t[1900] ^ n[1901];
assign t[1902] = t[1901] ^ n[1902];
assign t[1903] = t[1902] ^ n[1903];
assign t[1904] = t[1903] ^ n[1904];
assign t[1905] = t[1904] ^ n[1905];
assign t[1906] = t[1905] ^ n[1906];
assign t[1907] = t[1906] ^ n[1907];
assign t[1908] = t[1907] ^ n[1908];
assign t[1909] = t[1908] ^ n[1909];
assign t[1910] = t[1909] ^ n[1910];
assign t[1911] = t[1910] ^ n[1911];
assign t[1912] = t[1911] ^ n[1912];
assign t[1913] = t[1912] ^ n[1913];
assign t[1914] = t[1913] ^ n[1914];
assign t[1915] = t[1914] ^ n[1915];
assign t[1916] = t[1915] ^ n[1916];
assign t[1917] = t[1916] ^ n[1917];
assign t[1918] = t[1917] ^ n[1918];
assign t[1919] = t[1918] ^ n[1919];
assign t[1920] = t[1919] ^ n[1920];
assign t[1921] = t[1920] ^ n[1921];
assign t[1922] = t[1921] ^ n[1922];
assign t[1923] = t[1922] ^ n[1923];
assign t[1924] = t[1923] ^ n[1924];
assign t[1925] = t[1924] ^ n[1925];
assign t[1926] = t[1925] ^ n[1926];
assign t[1927] = t[1926] ^ n[1927];
assign t[1928] = t[1927] ^ n[1928];
assign t[1929] = t[1928] ^ n[1929];
assign t[1930] = t[1929] ^ n[1930];
assign t[1931] = t[1930] ^ n[1931];
assign t[1932] = t[1931] ^ n[1932];
assign t[1933] = t[1932] ^ n[1933];
assign t[1934] = t[1933] ^ n[1934];
assign t[1935] = t[1934] ^ n[1935];
assign t[1936] = t[1935] ^ n[1936];
assign t[1937] = t[1936] ^ n[1937];
assign t[1938] = t[1937] ^ n[1938];
assign t[1939] = t[1938] ^ n[1939];
assign t[1940] = t[1939] ^ n[1940];
assign t[1941] = t[1940] ^ n[1941];
assign t[1942] = t[1941] ^ n[1942];
assign t[1943] = t[1942] ^ n[1943];
assign t[1944] = t[1943] ^ n[1944];
assign t[1945] = t[1944] ^ n[1945];
assign t[1946] = t[1945] ^ n[1946];
assign t[1947] = t[1946] ^ n[1947];
assign t[1948] = t[1947] ^ n[1948];
assign t[1949] = t[1948] ^ n[1949];
assign t[1950] = t[1949] ^ n[1950];
assign t[1951] = t[1950] ^ n[1951];
assign t[1952] = t[1951] ^ n[1952];
assign t[1953] = t[1952] ^ n[1953];
assign t[1954] = t[1953] ^ n[1954];
assign t[1955] = t[1954] ^ n[1955];
assign t[1956] = t[1955] ^ n[1956];
assign t[1957] = t[1956] ^ n[1957];
assign t[1958] = t[1957] ^ n[1958];
assign t[1959] = t[1958] ^ n[1959];
assign t[1960] = t[1959] ^ n[1960];
assign t[1961] = t[1960] ^ n[1961];
assign t[1962] = t[1961] ^ n[1962];
assign t[1963] = t[1962] ^ n[1963];
assign t[1964] = t[1963] ^ n[1964];
assign t[1965] = t[1964] ^ n[1965];
assign t[1966] = t[1965] ^ n[1966];
assign t[1967] = t[1966] ^ n[1967];
assign t[1968] = t[1967] ^ n[1968];
assign t[1969] = t[1968] ^ n[1969];
assign t[1970] = t[1969] ^ n[1970];
assign t[1971] = t[1970] ^ n[1971];
assign t[1972] = t[1971] ^ n[1972];
assign t[1973] = t[1972] ^ n[1973];
assign t[1974] = t[1973] ^ n[1974];
assign t[1975] = t[1974] ^ n[1975];
assign t[1976] = t[1975] ^ n[1976];
assign t[1977] = t[1976] ^ n[1977];
assign t[1978] = t[1977] ^ n[1978];
assign t[1979] = t[1978] ^ n[1979];
assign t[1980] = t[1979] ^ n[1980];
assign t[1981] = t[1980] ^ n[1981];
assign t[1982] = t[1981] ^ n[1982];
assign t[1983] = t[1982] ^ n[1983];
assign t[1984] = t[1983] ^ n[1984];
assign t[1985] = t[1984] ^ n[1985];
assign t[1986] = t[1985] ^ n[1986];
assign t[1987] = t[1986] ^ n[1987];
assign t[1988] = t[1987] ^ n[1988];
assign t[1989] = t[1988] ^ n[1989];
assign t[1990] = t[1989] ^ n[1990];
assign t[1991] = t[1990] ^ n[1991];
assign t[1992] = t[1991] ^ n[1992];
assign t[1993] = t[1992] ^ n[1993];
assign t[1994] = t[1993] ^ n[1994];
assign t[1995] = t[1994] ^ n[1995];
assign t[1996] = t[1995] ^ n[1996];
assign t[1997] = t[1996] ^ n[1997];
assign t[1998] = t[1997] ^ n[1998];
assign t[1999] = t[1998] ^ n[1999];
assign t[2000] = t[1999] ^ n[2000];
assign t[2001] = t[2000] ^ n[2001];
assign t[2002] = t[2001] ^ n[2002];
assign t[2003] = t[2002] ^ n[2003];
assign t[2004] = t[2003] ^ n[2004];
assign t[2005] = t[2004] ^ n[2005];
assign t[2006] = t[2005] ^ n[2006];
assign t[2007] = t[2006] ^ n[2007];
assign t[2008] = t[2007] ^ n[2008];
assign t[2009] = t[2008] ^ n[2009];
assign t[2010] = t[2009] ^ n[2010];
assign t[2011] = t[2010] ^ n[2011];
assign t[2012] = t[2011] ^ n[2012];
assign t[2013] = t[2012] ^ n[2013];
assign t[2014] = t[2013] ^ n[2014];
assign t[2015] = t[2014] ^ n[2015];
assign t[2016] = t[2015] ^ n[2016];
assign t[2017] = t[2016] ^ n[2017];
assign t[2018] = t[2017] ^ n[2018];
assign t[2019] = t[2018] ^ n[2019];
assign t[2020] = t[2019] ^ n[2020];
assign t[2021] = t[2020] ^ n[2021];
assign t[2022] = t[2021] ^ n[2022];
assign t[2023] = t[2022] ^ n[2023];
assign t[2024] = t[2023] ^ n[2024];
assign t[2025] = t[2024] ^ n[2025];
assign t[2026] = t[2025] ^ n[2026];
assign t[2027] = t[2026] ^ n[2027];
assign t[2028] = t[2027] ^ n[2028];
assign t[2029] = t[2028] ^ n[2029];
assign t[2030] = t[2029] ^ n[2030];
assign t[2031] = t[2030] ^ n[2031];
assign t[2032] = t[2031] ^ n[2032];
assign t[2033] = t[2032] ^ n[2033];
assign t[2034] = t[2033] ^ n[2034];

assign s[9] = ( a[9] ^ b [9] ) ^ t[2034];

//asigning bit 10
assign t[2035] = n[2035];
assign t[2036] = t[2035] ^ n[2036];
assign t[2037] = t[2036] ^ n[2037];
assign t[2038] = t[2037] ^ n[2038];
assign t[2039] = t[2038] ^ n[2039];
assign t[2040] = t[2039] ^ n[2040];
assign t[2041] = t[2040] ^ n[2041];
assign t[2042] = t[2041] ^ n[2042];
assign t[2043] = t[2042] ^ n[2043];
assign t[2044] = t[2043] ^ n[2044];
assign t[2045] = t[2044] ^ n[2045];
assign t[2046] = t[2045] ^ n[2046];
assign t[2047] = t[2046] ^ n[2047];
assign t[2048] = t[2047] ^ n[2048];
assign t[2049] = t[2048] ^ n[2049];
assign t[2050] = t[2049] ^ n[2050];
assign t[2051] = t[2050] ^ n[2051];
assign t[2052] = t[2051] ^ n[2052];
assign t[2053] = t[2052] ^ n[2053];
assign t[2054] = t[2053] ^ n[2054];
assign t[2055] = t[2054] ^ n[2055];
assign t[2056] = t[2055] ^ n[2056];
assign t[2057] = t[2056] ^ n[2057];
assign t[2058] = t[2057] ^ n[2058];
assign t[2059] = t[2058] ^ n[2059];
assign t[2060] = t[2059] ^ n[2060];
assign t[2061] = t[2060] ^ n[2061];
assign t[2062] = t[2061] ^ n[2062];
assign t[2063] = t[2062] ^ n[2063];
assign t[2064] = t[2063] ^ n[2064];
assign t[2065] = t[2064] ^ n[2065];
assign t[2066] = t[2065] ^ n[2066];
assign t[2067] = t[2066] ^ n[2067];
assign t[2068] = t[2067] ^ n[2068];
assign t[2069] = t[2068] ^ n[2069];
assign t[2070] = t[2069] ^ n[2070];
assign t[2071] = t[2070] ^ n[2071];
assign t[2072] = t[2071] ^ n[2072];
assign t[2073] = t[2072] ^ n[2073];
assign t[2074] = t[2073] ^ n[2074];
assign t[2075] = t[2074] ^ n[2075];
assign t[2076] = t[2075] ^ n[2076];
assign t[2077] = t[2076] ^ n[2077];
assign t[2078] = t[2077] ^ n[2078];
assign t[2079] = t[2078] ^ n[2079];
assign t[2080] = t[2079] ^ n[2080];
assign t[2081] = t[2080] ^ n[2081];
assign t[2082] = t[2081] ^ n[2082];
assign t[2083] = t[2082] ^ n[2083];
assign t[2084] = t[2083] ^ n[2084];
assign t[2085] = t[2084] ^ n[2085];
assign t[2086] = t[2085] ^ n[2086];
assign t[2087] = t[2086] ^ n[2087];
assign t[2088] = t[2087] ^ n[2088];
assign t[2089] = t[2088] ^ n[2089];
assign t[2090] = t[2089] ^ n[2090];
assign t[2091] = t[2090] ^ n[2091];
assign t[2092] = t[2091] ^ n[2092];
assign t[2093] = t[2092] ^ n[2093];
assign t[2094] = t[2093] ^ n[2094];
assign t[2095] = t[2094] ^ n[2095];
assign t[2096] = t[2095] ^ n[2096];
assign t[2097] = t[2096] ^ n[2097];
assign t[2098] = t[2097] ^ n[2098];
assign t[2099] = t[2098] ^ n[2099];
assign t[2100] = t[2099] ^ n[2100];
assign t[2101] = t[2100] ^ n[2101];
assign t[2102] = t[2101] ^ n[2102];
assign t[2103] = t[2102] ^ n[2103];
assign t[2104] = t[2103] ^ n[2104];
assign t[2105] = t[2104] ^ n[2105];
assign t[2106] = t[2105] ^ n[2106];
assign t[2107] = t[2106] ^ n[2107];
assign t[2108] = t[2107] ^ n[2108];
assign t[2109] = t[2108] ^ n[2109];
assign t[2110] = t[2109] ^ n[2110];
assign t[2111] = t[2110] ^ n[2111];
assign t[2112] = t[2111] ^ n[2112];
assign t[2113] = t[2112] ^ n[2113];
assign t[2114] = t[2113] ^ n[2114];
assign t[2115] = t[2114] ^ n[2115];
assign t[2116] = t[2115] ^ n[2116];
assign t[2117] = t[2116] ^ n[2117];
assign t[2118] = t[2117] ^ n[2118];
assign t[2119] = t[2118] ^ n[2119];
assign t[2120] = t[2119] ^ n[2120];
assign t[2121] = t[2120] ^ n[2121];
assign t[2122] = t[2121] ^ n[2122];
assign t[2123] = t[2122] ^ n[2123];
assign t[2124] = t[2123] ^ n[2124];
assign t[2125] = t[2124] ^ n[2125];
assign t[2126] = t[2125] ^ n[2126];
assign t[2127] = t[2126] ^ n[2127];
assign t[2128] = t[2127] ^ n[2128];
assign t[2129] = t[2128] ^ n[2129];
assign t[2130] = t[2129] ^ n[2130];
assign t[2131] = t[2130] ^ n[2131];
assign t[2132] = t[2131] ^ n[2132];
assign t[2133] = t[2132] ^ n[2133];
assign t[2134] = t[2133] ^ n[2134];
assign t[2135] = t[2134] ^ n[2135];
assign t[2136] = t[2135] ^ n[2136];
assign t[2137] = t[2136] ^ n[2137];
assign t[2138] = t[2137] ^ n[2138];
assign t[2139] = t[2138] ^ n[2139];
assign t[2140] = t[2139] ^ n[2140];
assign t[2141] = t[2140] ^ n[2141];
assign t[2142] = t[2141] ^ n[2142];
assign t[2143] = t[2142] ^ n[2143];
assign t[2144] = t[2143] ^ n[2144];
assign t[2145] = t[2144] ^ n[2145];
assign t[2146] = t[2145] ^ n[2146];
assign t[2147] = t[2146] ^ n[2147];
assign t[2148] = t[2147] ^ n[2148];
assign t[2149] = t[2148] ^ n[2149];
assign t[2150] = t[2149] ^ n[2150];
assign t[2151] = t[2150] ^ n[2151];
assign t[2152] = t[2151] ^ n[2152];
assign t[2153] = t[2152] ^ n[2153];
assign t[2154] = t[2153] ^ n[2154];
assign t[2155] = t[2154] ^ n[2155];
assign t[2156] = t[2155] ^ n[2156];
assign t[2157] = t[2156] ^ n[2157];
assign t[2158] = t[2157] ^ n[2158];
assign t[2159] = t[2158] ^ n[2159];
assign t[2160] = t[2159] ^ n[2160];
assign t[2161] = t[2160] ^ n[2161];
assign t[2162] = t[2161] ^ n[2162];
assign t[2163] = t[2162] ^ n[2163];
assign t[2164] = t[2163] ^ n[2164];
assign t[2165] = t[2164] ^ n[2165];
assign t[2166] = t[2165] ^ n[2166];
assign t[2167] = t[2166] ^ n[2167];
assign t[2168] = t[2167] ^ n[2168];
assign t[2169] = t[2168] ^ n[2169];
assign t[2170] = t[2169] ^ n[2170];
assign t[2171] = t[2170] ^ n[2171];
assign t[2172] = t[2171] ^ n[2172];
assign t[2173] = t[2172] ^ n[2173];
assign t[2174] = t[2173] ^ n[2174];
assign t[2175] = t[2174] ^ n[2175];
assign t[2176] = t[2175] ^ n[2176];
assign t[2177] = t[2176] ^ n[2177];
assign t[2178] = t[2177] ^ n[2178];
assign t[2179] = t[2178] ^ n[2179];
assign t[2180] = t[2179] ^ n[2180];
assign t[2181] = t[2180] ^ n[2181];
assign t[2182] = t[2181] ^ n[2182];
assign t[2183] = t[2182] ^ n[2183];
assign t[2184] = t[2183] ^ n[2184];
assign t[2185] = t[2184] ^ n[2185];
assign t[2186] = t[2185] ^ n[2186];
assign t[2187] = t[2186] ^ n[2187];
assign t[2188] = t[2187] ^ n[2188];
assign t[2189] = t[2188] ^ n[2189];
assign t[2190] = t[2189] ^ n[2190];
assign t[2191] = t[2190] ^ n[2191];
assign t[2192] = t[2191] ^ n[2192];
assign t[2193] = t[2192] ^ n[2193];
assign t[2194] = t[2193] ^ n[2194];
assign t[2195] = t[2194] ^ n[2195];
assign t[2196] = t[2195] ^ n[2196];
assign t[2197] = t[2196] ^ n[2197];
assign t[2198] = t[2197] ^ n[2198];
assign t[2199] = t[2198] ^ n[2199];
assign t[2200] = t[2199] ^ n[2200];
assign t[2201] = t[2200] ^ n[2201];
assign t[2202] = t[2201] ^ n[2202];
assign t[2203] = t[2202] ^ n[2203];
assign t[2204] = t[2203] ^ n[2204];
assign t[2205] = t[2204] ^ n[2205];
assign t[2206] = t[2205] ^ n[2206];
assign t[2207] = t[2206] ^ n[2207];
assign t[2208] = t[2207] ^ n[2208];
assign t[2209] = t[2208] ^ n[2209];
assign t[2210] = t[2209] ^ n[2210];
assign t[2211] = t[2210] ^ n[2211];
assign t[2212] = t[2211] ^ n[2212];
assign t[2213] = t[2212] ^ n[2213];
assign t[2214] = t[2213] ^ n[2214];
assign t[2215] = t[2214] ^ n[2215];
assign t[2216] = t[2215] ^ n[2216];
assign t[2217] = t[2216] ^ n[2217];
assign t[2218] = t[2217] ^ n[2218];
assign t[2219] = t[2218] ^ n[2219];
assign t[2220] = t[2219] ^ n[2220];
assign t[2221] = t[2220] ^ n[2221];
assign t[2222] = t[2221] ^ n[2222];
assign t[2223] = t[2222] ^ n[2223];
assign t[2224] = t[2223] ^ n[2224];
assign t[2225] = t[2224] ^ n[2225];
assign t[2226] = t[2225] ^ n[2226];
assign t[2227] = t[2226] ^ n[2227];
assign t[2228] = t[2227] ^ n[2228];
assign t[2229] = t[2228] ^ n[2229];
assign t[2230] = t[2229] ^ n[2230];
assign t[2231] = t[2230] ^ n[2231];
assign t[2232] = t[2231] ^ n[2232];
assign t[2233] = t[2232] ^ n[2233];
assign t[2234] = t[2233] ^ n[2234];
assign t[2235] = t[2234] ^ n[2235];
assign t[2236] = t[2235] ^ n[2236];
assign t[2237] = t[2236] ^ n[2237];
assign t[2238] = t[2237] ^ n[2238];
assign t[2239] = t[2238] ^ n[2239];
assign t[2240] = t[2239] ^ n[2240];
assign t[2241] = t[2240] ^ n[2241];
assign t[2242] = t[2241] ^ n[2242];
assign t[2243] = t[2242] ^ n[2243];
assign t[2244] = t[2243] ^ n[2244];
assign t[2245] = t[2244] ^ n[2245];
assign t[2246] = t[2245] ^ n[2246];
assign t[2247] = t[2246] ^ n[2247];
assign t[2248] = t[2247] ^ n[2248];
assign t[2249] = t[2248] ^ n[2249];
assign t[2250] = t[2249] ^ n[2250];
assign t[2251] = t[2250] ^ n[2251];
assign t[2252] = t[2251] ^ n[2252];
assign t[2253] = t[2252] ^ n[2253];
assign t[2254] = t[2253] ^ n[2254];
assign t[2255] = t[2254] ^ n[2255];
assign t[2256] = t[2255] ^ n[2256];
assign t[2257] = t[2256] ^ n[2257];
assign t[2258] = t[2257] ^ n[2258];
assign t[2259] = t[2258] ^ n[2259];
assign t[2260] = t[2259] ^ n[2260];
assign t[2261] = t[2260] ^ n[2261];
assign t[2262] = t[2261] ^ n[2262];
assign t[2263] = t[2262] ^ n[2263];
assign t[2264] = t[2263] ^ n[2264];
assign t[2265] = t[2264] ^ n[2265];
assign t[2266] = t[2265] ^ n[2266];
assign t[2267] = t[2266] ^ n[2267];
assign t[2268] = t[2267] ^ n[2268];
assign t[2269] = t[2268] ^ n[2269];
assign t[2270] = t[2269] ^ n[2270];
assign t[2271] = t[2270] ^ n[2271];
assign t[2272] = t[2271] ^ n[2272];
assign t[2273] = t[2272] ^ n[2273];
assign t[2274] = t[2273] ^ n[2274];
assign t[2275] = t[2274] ^ n[2275];
assign t[2276] = t[2275] ^ n[2276];
assign t[2277] = t[2276] ^ n[2277];
assign t[2278] = t[2277] ^ n[2278];
assign t[2279] = t[2278] ^ n[2279];
assign t[2280] = t[2279] ^ n[2280];
assign t[2281] = t[2280] ^ n[2281];
assign t[2282] = t[2281] ^ n[2282];
assign t[2283] = t[2282] ^ n[2283];
assign t[2284] = t[2283] ^ n[2284];
assign t[2285] = t[2284] ^ n[2285];
assign t[2286] = t[2285] ^ n[2286];
assign t[2287] = t[2286] ^ n[2287];
assign t[2288] = t[2287] ^ n[2288];
assign t[2289] = t[2288] ^ n[2289];
assign t[2290] = t[2289] ^ n[2290];
assign t[2291] = t[2290] ^ n[2291];
assign t[2292] = t[2291] ^ n[2292];
assign t[2293] = t[2292] ^ n[2293];
assign t[2294] = t[2293] ^ n[2294];
assign t[2295] = t[2294] ^ n[2295];
assign t[2296] = t[2295] ^ n[2296];
assign t[2297] = t[2296] ^ n[2297];
assign t[2298] = t[2297] ^ n[2298];
assign t[2299] = t[2298] ^ n[2299];
assign t[2300] = t[2299] ^ n[2300];
assign t[2301] = t[2300] ^ n[2301];
assign t[2302] = t[2301] ^ n[2302];
assign t[2303] = t[2302] ^ n[2303];
assign t[2304] = t[2303] ^ n[2304];
assign t[2305] = t[2304] ^ n[2305];
assign t[2306] = t[2305] ^ n[2306];
assign t[2307] = t[2306] ^ n[2307];
assign t[2308] = t[2307] ^ n[2308];
assign t[2309] = t[2308] ^ n[2309];
assign t[2310] = t[2309] ^ n[2310];
assign t[2311] = t[2310] ^ n[2311];
assign t[2312] = t[2311] ^ n[2312];
assign t[2313] = t[2312] ^ n[2313];
assign t[2314] = t[2313] ^ n[2314];
assign t[2315] = t[2314] ^ n[2315];
assign t[2316] = t[2315] ^ n[2316];
assign t[2317] = t[2316] ^ n[2317];
assign t[2318] = t[2317] ^ n[2318];
assign t[2319] = t[2318] ^ n[2319];
assign t[2320] = t[2319] ^ n[2320];
assign t[2321] = t[2320] ^ n[2321];
assign t[2322] = t[2321] ^ n[2322];
assign t[2323] = t[2322] ^ n[2323];
assign t[2324] = t[2323] ^ n[2324];
assign t[2325] = t[2324] ^ n[2325];
assign t[2326] = t[2325] ^ n[2326];
assign t[2327] = t[2326] ^ n[2327];
assign t[2328] = t[2327] ^ n[2328];
assign t[2329] = t[2328] ^ n[2329];
assign t[2330] = t[2329] ^ n[2330];
assign t[2331] = t[2330] ^ n[2331];
assign t[2332] = t[2331] ^ n[2332];
assign t[2333] = t[2332] ^ n[2333];
assign t[2334] = t[2333] ^ n[2334];
assign t[2335] = t[2334] ^ n[2335];
assign t[2336] = t[2335] ^ n[2336];
assign t[2337] = t[2336] ^ n[2337];
assign t[2338] = t[2337] ^ n[2338];
assign t[2339] = t[2338] ^ n[2339];
assign t[2340] = t[2339] ^ n[2340];
assign t[2341] = t[2340] ^ n[2341];
assign t[2342] = t[2341] ^ n[2342];
assign t[2343] = t[2342] ^ n[2343];
assign t[2344] = t[2343] ^ n[2344];
assign t[2345] = t[2344] ^ n[2345];
assign t[2346] = t[2345] ^ n[2346];
assign t[2347] = t[2346] ^ n[2347];
assign t[2348] = t[2347] ^ n[2348];
assign t[2349] = t[2348] ^ n[2349];
assign t[2350] = t[2349] ^ n[2350];
assign t[2351] = t[2350] ^ n[2351];
assign t[2352] = t[2351] ^ n[2352];
assign t[2353] = t[2352] ^ n[2353];
assign t[2354] = t[2353] ^ n[2354];
assign t[2355] = t[2354] ^ n[2355];
assign t[2356] = t[2355] ^ n[2356];
assign t[2357] = t[2356] ^ n[2357];
assign t[2358] = t[2357] ^ n[2358];
assign t[2359] = t[2358] ^ n[2359];
assign t[2360] = t[2359] ^ n[2360];
assign t[2361] = t[2360] ^ n[2361];
assign t[2362] = t[2361] ^ n[2362];
assign t[2363] = t[2362] ^ n[2363];
assign t[2364] = t[2363] ^ n[2364];
assign t[2365] = t[2364] ^ n[2365];
assign t[2366] = t[2365] ^ n[2366];
assign t[2367] = t[2366] ^ n[2367];
assign t[2368] = t[2367] ^ n[2368];
assign t[2369] = t[2368] ^ n[2369];
assign t[2370] = t[2369] ^ n[2370];
assign t[2371] = t[2370] ^ n[2371];
assign t[2372] = t[2371] ^ n[2372];
assign t[2373] = t[2372] ^ n[2373];
assign t[2374] = t[2373] ^ n[2374];
assign t[2375] = t[2374] ^ n[2375];
assign t[2376] = t[2375] ^ n[2376];
assign t[2377] = t[2376] ^ n[2377];
assign t[2378] = t[2377] ^ n[2378];
assign t[2379] = t[2378] ^ n[2379];
assign t[2380] = t[2379] ^ n[2380];
assign t[2381] = t[2380] ^ n[2381];
assign t[2382] = t[2381] ^ n[2382];
assign t[2383] = t[2382] ^ n[2383];
assign t[2384] = t[2383] ^ n[2384];
assign t[2385] = t[2384] ^ n[2385];
assign t[2386] = t[2385] ^ n[2386];
assign t[2387] = t[2386] ^ n[2387];
assign t[2388] = t[2387] ^ n[2388];
assign t[2389] = t[2388] ^ n[2389];
assign t[2390] = t[2389] ^ n[2390];
assign t[2391] = t[2390] ^ n[2391];
assign t[2392] = t[2391] ^ n[2392];
assign t[2393] = t[2392] ^ n[2393];
assign t[2394] = t[2393] ^ n[2394];
assign t[2395] = t[2394] ^ n[2395];
assign t[2396] = t[2395] ^ n[2396];
assign t[2397] = t[2396] ^ n[2397];
assign t[2398] = t[2397] ^ n[2398];
assign t[2399] = t[2398] ^ n[2399];
assign t[2400] = t[2399] ^ n[2400];
assign t[2401] = t[2400] ^ n[2401];
assign t[2402] = t[2401] ^ n[2402];
assign t[2403] = t[2402] ^ n[2403];
assign t[2404] = t[2403] ^ n[2404];
assign t[2405] = t[2404] ^ n[2405];
assign t[2406] = t[2405] ^ n[2406];
assign t[2407] = t[2406] ^ n[2407];
assign t[2408] = t[2407] ^ n[2408];
assign t[2409] = t[2408] ^ n[2409];
assign t[2410] = t[2409] ^ n[2410];
assign t[2411] = t[2410] ^ n[2411];
assign t[2412] = t[2411] ^ n[2412];
assign t[2413] = t[2412] ^ n[2413];
assign t[2414] = t[2413] ^ n[2414];
assign t[2415] = t[2414] ^ n[2415];
assign t[2416] = t[2415] ^ n[2416];
assign t[2417] = t[2416] ^ n[2417];
assign t[2418] = t[2417] ^ n[2418];
assign t[2419] = t[2418] ^ n[2419];
assign t[2420] = t[2419] ^ n[2420];
assign t[2421] = t[2420] ^ n[2421];
assign t[2422] = t[2421] ^ n[2422];
assign t[2423] = t[2422] ^ n[2423];
assign t[2424] = t[2423] ^ n[2424];
assign t[2425] = t[2424] ^ n[2425];
assign t[2426] = t[2425] ^ n[2426];
assign t[2427] = t[2426] ^ n[2427];
assign t[2428] = t[2427] ^ n[2428];
assign t[2429] = t[2428] ^ n[2429];
assign t[2430] = t[2429] ^ n[2430];
assign t[2431] = t[2430] ^ n[2431];
assign t[2432] = t[2431] ^ n[2432];
assign t[2433] = t[2432] ^ n[2433];
assign t[2434] = t[2433] ^ n[2434];
assign t[2435] = t[2434] ^ n[2435];
assign t[2436] = t[2435] ^ n[2436];
assign t[2437] = t[2436] ^ n[2437];
assign t[2438] = t[2437] ^ n[2438];
assign t[2439] = t[2438] ^ n[2439];
assign t[2440] = t[2439] ^ n[2440];
assign t[2441] = t[2440] ^ n[2441];
assign t[2442] = t[2441] ^ n[2442];
assign t[2443] = t[2442] ^ n[2443];
assign t[2444] = t[2443] ^ n[2444];
assign t[2445] = t[2444] ^ n[2445];
assign t[2446] = t[2445] ^ n[2446];
assign t[2447] = t[2446] ^ n[2447];
assign t[2448] = t[2447] ^ n[2448];
assign t[2449] = t[2448] ^ n[2449];
assign t[2450] = t[2449] ^ n[2450];
assign t[2451] = t[2450] ^ n[2451];
assign t[2452] = t[2451] ^ n[2452];
assign t[2453] = t[2452] ^ n[2453];
assign t[2454] = t[2453] ^ n[2454];
assign t[2455] = t[2454] ^ n[2455];
assign t[2456] = t[2455] ^ n[2456];
assign t[2457] = t[2456] ^ n[2457];
assign t[2458] = t[2457] ^ n[2458];
assign t[2459] = t[2458] ^ n[2459];
assign t[2460] = t[2459] ^ n[2460];
assign t[2461] = t[2460] ^ n[2461];
assign t[2462] = t[2461] ^ n[2462];
assign t[2463] = t[2462] ^ n[2463];
assign t[2464] = t[2463] ^ n[2464];
assign t[2465] = t[2464] ^ n[2465];
assign t[2466] = t[2465] ^ n[2466];
assign t[2467] = t[2466] ^ n[2467];
assign t[2468] = t[2467] ^ n[2468];
assign t[2469] = t[2468] ^ n[2469];
assign t[2470] = t[2469] ^ n[2470];
assign t[2471] = t[2470] ^ n[2471];
assign t[2472] = t[2471] ^ n[2472];
assign t[2473] = t[2472] ^ n[2473];
assign t[2474] = t[2473] ^ n[2474];
assign t[2475] = t[2474] ^ n[2475];
assign t[2476] = t[2475] ^ n[2476];
assign t[2477] = t[2476] ^ n[2477];
assign t[2478] = t[2477] ^ n[2478];
assign t[2479] = t[2478] ^ n[2479];
assign t[2480] = t[2479] ^ n[2480];
assign t[2481] = t[2480] ^ n[2481];
assign t[2482] = t[2481] ^ n[2482];
assign t[2483] = t[2482] ^ n[2483];
assign t[2484] = t[2483] ^ n[2484];
assign t[2485] = t[2484] ^ n[2485];
assign t[2486] = t[2485] ^ n[2486];
assign t[2487] = t[2486] ^ n[2487];
assign t[2488] = t[2487] ^ n[2488];
assign t[2489] = t[2488] ^ n[2489];
assign t[2490] = t[2489] ^ n[2490];
assign t[2491] = t[2490] ^ n[2491];
assign t[2492] = t[2491] ^ n[2492];
assign t[2493] = t[2492] ^ n[2493];
assign t[2494] = t[2493] ^ n[2494];
assign t[2495] = t[2494] ^ n[2495];
assign t[2496] = t[2495] ^ n[2496];
assign t[2497] = t[2496] ^ n[2497];
assign t[2498] = t[2497] ^ n[2498];
assign t[2499] = t[2498] ^ n[2499];
assign t[2500] = t[2499] ^ n[2500];
assign t[2501] = t[2500] ^ n[2501];
assign t[2502] = t[2501] ^ n[2502];
assign t[2503] = t[2502] ^ n[2503];
assign t[2504] = t[2503] ^ n[2504];
assign t[2505] = t[2504] ^ n[2505];
assign t[2506] = t[2505] ^ n[2506];
assign t[2507] = t[2506] ^ n[2507];
assign t[2508] = t[2507] ^ n[2508];
assign t[2509] = t[2508] ^ n[2509];
assign t[2510] = t[2509] ^ n[2510];
assign t[2511] = t[2510] ^ n[2511];
assign t[2512] = t[2511] ^ n[2512];
assign t[2513] = t[2512] ^ n[2513];
assign t[2514] = t[2513] ^ n[2514];
assign t[2515] = t[2514] ^ n[2515];
assign t[2516] = t[2515] ^ n[2516];
assign t[2517] = t[2516] ^ n[2517];
assign t[2518] = t[2517] ^ n[2518];
assign t[2519] = t[2518] ^ n[2519];
assign t[2520] = t[2519] ^ n[2520];
assign t[2521] = t[2520] ^ n[2521];
assign t[2522] = t[2521] ^ n[2522];
assign t[2523] = t[2522] ^ n[2523];
assign t[2524] = t[2523] ^ n[2524];
assign t[2525] = t[2524] ^ n[2525];
assign t[2526] = t[2525] ^ n[2526];
assign t[2527] = t[2526] ^ n[2527];
assign t[2528] = t[2527] ^ n[2528];
assign t[2529] = t[2528] ^ n[2529];
assign t[2530] = t[2529] ^ n[2530];
assign t[2531] = t[2530] ^ n[2531];
assign t[2532] = t[2531] ^ n[2532];
assign t[2533] = t[2532] ^ n[2533];
assign t[2534] = t[2533] ^ n[2534];
assign t[2535] = t[2534] ^ n[2535];
assign t[2536] = t[2535] ^ n[2536];
assign t[2537] = t[2536] ^ n[2537];
assign t[2538] = t[2537] ^ n[2538];
assign t[2539] = t[2538] ^ n[2539];
assign t[2540] = t[2539] ^ n[2540];
assign t[2541] = t[2540] ^ n[2541];
assign t[2542] = t[2541] ^ n[2542];
assign t[2543] = t[2542] ^ n[2543];
assign t[2544] = t[2543] ^ n[2544];
assign t[2545] = t[2544] ^ n[2545];
assign t[2546] = t[2545] ^ n[2546];
assign t[2547] = t[2546] ^ n[2547];
assign t[2548] = t[2547] ^ n[2548];
assign t[2549] = t[2548] ^ n[2549];
assign t[2550] = t[2549] ^ n[2550];
assign t[2551] = t[2550] ^ n[2551];
assign t[2552] = t[2551] ^ n[2552];
assign t[2553] = t[2552] ^ n[2553];
assign t[2554] = t[2553] ^ n[2554];
assign t[2555] = t[2554] ^ n[2555];
assign t[2556] = t[2555] ^ n[2556];
assign t[2557] = t[2556] ^ n[2557];
assign t[2558] = t[2557] ^ n[2558];
assign t[2559] = t[2558] ^ n[2559];
assign t[2560] = t[2559] ^ n[2560];
assign t[2561] = t[2560] ^ n[2561];
assign t[2562] = t[2561] ^ n[2562];
assign t[2563] = t[2562] ^ n[2563];
assign t[2564] = t[2563] ^ n[2564];
assign t[2565] = t[2564] ^ n[2565];
assign t[2566] = t[2565] ^ n[2566];
assign t[2567] = t[2566] ^ n[2567];
assign t[2568] = t[2567] ^ n[2568];
assign t[2569] = t[2568] ^ n[2569];
assign t[2570] = t[2569] ^ n[2570];
assign t[2571] = t[2570] ^ n[2571];
assign t[2572] = t[2571] ^ n[2572];
assign t[2573] = t[2572] ^ n[2573];
assign t[2574] = t[2573] ^ n[2574];
assign t[2575] = t[2574] ^ n[2575];
assign t[2576] = t[2575] ^ n[2576];
assign t[2577] = t[2576] ^ n[2577];
assign t[2578] = t[2577] ^ n[2578];
assign t[2579] = t[2578] ^ n[2579];
assign t[2580] = t[2579] ^ n[2580];
assign t[2581] = t[2580] ^ n[2581];
assign t[2582] = t[2581] ^ n[2582];
assign t[2583] = t[2582] ^ n[2583];
assign t[2584] = t[2583] ^ n[2584];
assign t[2585] = t[2584] ^ n[2585];
assign t[2586] = t[2585] ^ n[2586];
assign t[2587] = t[2586] ^ n[2587];
assign t[2588] = t[2587] ^ n[2588];
assign t[2589] = t[2588] ^ n[2589];
assign t[2590] = t[2589] ^ n[2590];
assign t[2591] = t[2590] ^ n[2591];
assign t[2592] = t[2591] ^ n[2592];
assign t[2593] = t[2592] ^ n[2593];
assign t[2594] = t[2593] ^ n[2594];
assign t[2595] = t[2594] ^ n[2595];
assign t[2596] = t[2595] ^ n[2596];
assign t[2597] = t[2596] ^ n[2597];
assign t[2598] = t[2597] ^ n[2598];
assign t[2599] = t[2598] ^ n[2599];
assign t[2600] = t[2599] ^ n[2600];
assign t[2601] = t[2600] ^ n[2601];
assign t[2602] = t[2601] ^ n[2602];
assign t[2603] = t[2602] ^ n[2603];
assign t[2604] = t[2603] ^ n[2604];
assign t[2605] = t[2604] ^ n[2605];
assign t[2606] = t[2605] ^ n[2606];
assign t[2607] = t[2606] ^ n[2607];
assign t[2608] = t[2607] ^ n[2608];
assign t[2609] = t[2608] ^ n[2609];
assign t[2610] = t[2609] ^ n[2610];
assign t[2611] = t[2610] ^ n[2611];
assign t[2612] = t[2611] ^ n[2612];
assign t[2613] = t[2612] ^ n[2613];
assign t[2614] = t[2613] ^ n[2614];
assign t[2615] = t[2614] ^ n[2615];
assign t[2616] = t[2615] ^ n[2616];
assign t[2617] = t[2616] ^ n[2617];
assign t[2618] = t[2617] ^ n[2618];
assign t[2619] = t[2618] ^ n[2619];
assign t[2620] = t[2619] ^ n[2620];
assign t[2621] = t[2620] ^ n[2621];
assign t[2622] = t[2621] ^ n[2622];
assign t[2623] = t[2622] ^ n[2623];
assign t[2624] = t[2623] ^ n[2624];
assign t[2625] = t[2624] ^ n[2625];
assign t[2626] = t[2625] ^ n[2626];
assign t[2627] = t[2626] ^ n[2627];
assign t[2628] = t[2627] ^ n[2628];
assign t[2629] = t[2628] ^ n[2629];
assign t[2630] = t[2629] ^ n[2630];
assign t[2631] = t[2630] ^ n[2631];
assign t[2632] = t[2631] ^ n[2632];
assign t[2633] = t[2632] ^ n[2633];
assign t[2634] = t[2633] ^ n[2634];
assign t[2635] = t[2634] ^ n[2635];
assign t[2636] = t[2635] ^ n[2636];
assign t[2637] = t[2636] ^ n[2637];
assign t[2638] = t[2637] ^ n[2638];
assign t[2639] = t[2638] ^ n[2639];
assign t[2640] = t[2639] ^ n[2640];
assign t[2641] = t[2640] ^ n[2641];
assign t[2642] = t[2641] ^ n[2642];
assign t[2643] = t[2642] ^ n[2643];
assign t[2644] = t[2643] ^ n[2644];
assign t[2645] = t[2644] ^ n[2645];
assign t[2646] = t[2645] ^ n[2646];
assign t[2647] = t[2646] ^ n[2647];
assign t[2648] = t[2647] ^ n[2648];
assign t[2649] = t[2648] ^ n[2649];
assign t[2650] = t[2649] ^ n[2650];
assign t[2651] = t[2650] ^ n[2651];
assign t[2652] = t[2651] ^ n[2652];
assign t[2653] = t[2652] ^ n[2653];
assign t[2654] = t[2653] ^ n[2654];
assign t[2655] = t[2654] ^ n[2655];
assign t[2656] = t[2655] ^ n[2656];
assign t[2657] = t[2656] ^ n[2657];
assign t[2658] = t[2657] ^ n[2658];
assign t[2659] = t[2658] ^ n[2659];
assign t[2660] = t[2659] ^ n[2660];
assign t[2661] = t[2660] ^ n[2661];
assign t[2662] = t[2661] ^ n[2662];
assign t[2663] = t[2662] ^ n[2663];
assign t[2664] = t[2663] ^ n[2664];
assign t[2665] = t[2664] ^ n[2665];
assign t[2666] = t[2665] ^ n[2666];
assign t[2667] = t[2666] ^ n[2667];
assign t[2668] = t[2667] ^ n[2668];
assign t[2669] = t[2668] ^ n[2669];
assign t[2670] = t[2669] ^ n[2670];
assign t[2671] = t[2670] ^ n[2671];
assign t[2672] = t[2671] ^ n[2672];
assign t[2673] = t[2672] ^ n[2673];
assign t[2674] = t[2673] ^ n[2674];
assign t[2675] = t[2674] ^ n[2675];
assign t[2676] = t[2675] ^ n[2676];
assign t[2677] = t[2676] ^ n[2677];
assign t[2678] = t[2677] ^ n[2678];
assign t[2679] = t[2678] ^ n[2679];
assign t[2680] = t[2679] ^ n[2680];
assign t[2681] = t[2680] ^ n[2681];
assign t[2682] = t[2681] ^ n[2682];
assign t[2683] = t[2682] ^ n[2683];
assign t[2684] = t[2683] ^ n[2684];
assign t[2685] = t[2684] ^ n[2685];
assign t[2686] = t[2685] ^ n[2686];
assign t[2687] = t[2686] ^ n[2687];
assign t[2688] = t[2687] ^ n[2688];
assign t[2689] = t[2688] ^ n[2689];
assign t[2690] = t[2689] ^ n[2690];
assign t[2691] = t[2690] ^ n[2691];
assign t[2692] = t[2691] ^ n[2692];
assign t[2693] = t[2692] ^ n[2693];
assign t[2694] = t[2693] ^ n[2694];
assign t[2695] = t[2694] ^ n[2695];
assign t[2696] = t[2695] ^ n[2696];
assign t[2697] = t[2696] ^ n[2697];
assign t[2698] = t[2697] ^ n[2698];
assign t[2699] = t[2698] ^ n[2699];
assign t[2700] = t[2699] ^ n[2700];
assign t[2701] = t[2700] ^ n[2701];
assign t[2702] = t[2701] ^ n[2702];
assign t[2703] = t[2702] ^ n[2703];
assign t[2704] = t[2703] ^ n[2704];
assign t[2705] = t[2704] ^ n[2705];
assign t[2706] = t[2705] ^ n[2706];
assign t[2707] = t[2706] ^ n[2707];
assign t[2708] = t[2707] ^ n[2708];
assign t[2709] = t[2708] ^ n[2709];
assign t[2710] = t[2709] ^ n[2710];
assign t[2711] = t[2710] ^ n[2711];
assign t[2712] = t[2711] ^ n[2712];
assign t[2713] = t[2712] ^ n[2713];
assign t[2714] = t[2713] ^ n[2714];
assign t[2715] = t[2714] ^ n[2715];
assign t[2716] = t[2715] ^ n[2716];
assign t[2717] = t[2716] ^ n[2717];
assign t[2718] = t[2717] ^ n[2718];
assign t[2719] = t[2718] ^ n[2719];
assign t[2720] = t[2719] ^ n[2720];
assign t[2721] = t[2720] ^ n[2721];
assign t[2722] = t[2721] ^ n[2722];
assign t[2723] = t[2722] ^ n[2723];
assign t[2724] = t[2723] ^ n[2724];
assign t[2725] = t[2724] ^ n[2725];
assign t[2726] = t[2725] ^ n[2726];
assign t[2727] = t[2726] ^ n[2727];
assign t[2728] = t[2727] ^ n[2728];
assign t[2729] = t[2728] ^ n[2729];
assign t[2730] = t[2729] ^ n[2730];
assign t[2731] = t[2730] ^ n[2731];
assign t[2732] = t[2731] ^ n[2732];
assign t[2733] = t[2732] ^ n[2733];
assign t[2734] = t[2733] ^ n[2734];
assign t[2735] = t[2734] ^ n[2735];
assign t[2736] = t[2735] ^ n[2736];
assign t[2737] = t[2736] ^ n[2737];
assign t[2738] = t[2737] ^ n[2738];
assign t[2739] = t[2738] ^ n[2739];
assign t[2740] = t[2739] ^ n[2740];
assign t[2741] = t[2740] ^ n[2741];
assign t[2742] = t[2741] ^ n[2742];
assign t[2743] = t[2742] ^ n[2743];
assign t[2744] = t[2743] ^ n[2744];
assign t[2745] = t[2744] ^ n[2745];
assign t[2746] = t[2745] ^ n[2746];
assign t[2747] = t[2746] ^ n[2747];
assign t[2748] = t[2747] ^ n[2748];
assign t[2749] = t[2748] ^ n[2749];
assign t[2750] = t[2749] ^ n[2750];
assign t[2751] = t[2750] ^ n[2751];
assign t[2752] = t[2751] ^ n[2752];
assign t[2753] = t[2752] ^ n[2753];
assign t[2754] = t[2753] ^ n[2754];
assign t[2755] = t[2754] ^ n[2755];
assign t[2756] = t[2755] ^ n[2756];
assign t[2757] = t[2756] ^ n[2757];
assign t[2758] = t[2757] ^ n[2758];
assign t[2759] = t[2758] ^ n[2759];
assign t[2760] = t[2759] ^ n[2760];
assign t[2761] = t[2760] ^ n[2761];
assign t[2762] = t[2761] ^ n[2762];
assign t[2763] = t[2762] ^ n[2763];
assign t[2764] = t[2763] ^ n[2764];
assign t[2765] = t[2764] ^ n[2765];
assign t[2766] = t[2765] ^ n[2766];
assign t[2767] = t[2766] ^ n[2767];
assign t[2768] = t[2767] ^ n[2768];
assign t[2769] = t[2768] ^ n[2769];
assign t[2770] = t[2769] ^ n[2770];
assign t[2771] = t[2770] ^ n[2771];
assign t[2772] = t[2771] ^ n[2772];
assign t[2773] = t[2772] ^ n[2773];
assign t[2774] = t[2773] ^ n[2774];
assign t[2775] = t[2774] ^ n[2775];
assign t[2776] = t[2775] ^ n[2776];
assign t[2777] = t[2776] ^ n[2777];
assign t[2778] = t[2777] ^ n[2778];
assign t[2779] = t[2778] ^ n[2779];
assign t[2780] = t[2779] ^ n[2780];
assign t[2781] = t[2780] ^ n[2781];
assign t[2782] = t[2781] ^ n[2782];
assign t[2783] = t[2782] ^ n[2783];
assign t[2784] = t[2783] ^ n[2784];
assign t[2785] = t[2784] ^ n[2785];
assign t[2786] = t[2785] ^ n[2786];
assign t[2787] = t[2786] ^ n[2787];
assign t[2788] = t[2787] ^ n[2788];
assign t[2789] = t[2788] ^ n[2789];
assign t[2790] = t[2789] ^ n[2790];
assign t[2791] = t[2790] ^ n[2791];
assign t[2792] = t[2791] ^ n[2792];
assign t[2793] = t[2792] ^ n[2793];
assign t[2794] = t[2793] ^ n[2794];
assign t[2795] = t[2794] ^ n[2795];
assign t[2796] = t[2795] ^ n[2796];
assign t[2797] = t[2796] ^ n[2797];
assign t[2798] = t[2797] ^ n[2798];
assign t[2799] = t[2798] ^ n[2799];
assign t[2800] = t[2799] ^ n[2800];
assign t[2801] = t[2800] ^ n[2801];
assign t[2802] = t[2801] ^ n[2802];
assign t[2803] = t[2802] ^ n[2803];
assign t[2804] = t[2803] ^ n[2804];
assign t[2805] = t[2804] ^ n[2805];
assign t[2806] = t[2805] ^ n[2806];
assign t[2807] = t[2806] ^ n[2807];
assign t[2808] = t[2807] ^ n[2808];
assign t[2809] = t[2808] ^ n[2809];
assign t[2810] = t[2809] ^ n[2810];
assign t[2811] = t[2810] ^ n[2811];
assign t[2812] = t[2811] ^ n[2812];
assign t[2813] = t[2812] ^ n[2813];
assign t[2814] = t[2813] ^ n[2814];
assign t[2815] = t[2814] ^ n[2815];
assign t[2816] = t[2815] ^ n[2816];
assign t[2817] = t[2816] ^ n[2817];
assign t[2818] = t[2817] ^ n[2818];
assign t[2819] = t[2818] ^ n[2819];
assign t[2820] = t[2819] ^ n[2820];
assign t[2821] = t[2820] ^ n[2821];
assign t[2822] = t[2821] ^ n[2822];
assign t[2823] = t[2822] ^ n[2823];
assign t[2824] = t[2823] ^ n[2824];
assign t[2825] = t[2824] ^ n[2825];
assign t[2826] = t[2825] ^ n[2826];
assign t[2827] = t[2826] ^ n[2827];
assign t[2828] = t[2827] ^ n[2828];
assign t[2829] = t[2828] ^ n[2829];
assign t[2830] = t[2829] ^ n[2830];
assign t[2831] = t[2830] ^ n[2831];
assign t[2832] = t[2831] ^ n[2832];
assign t[2833] = t[2832] ^ n[2833];
assign t[2834] = t[2833] ^ n[2834];
assign t[2835] = t[2834] ^ n[2835];
assign t[2836] = t[2835] ^ n[2836];
assign t[2837] = t[2836] ^ n[2837];
assign t[2838] = t[2837] ^ n[2838];
assign t[2839] = t[2838] ^ n[2839];
assign t[2840] = t[2839] ^ n[2840];
assign t[2841] = t[2840] ^ n[2841];
assign t[2842] = t[2841] ^ n[2842];
assign t[2843] = t[2842] ^ n[2843];
assign t[2844] = t[2843] ^ n[2844];
assign t[2845] = t[2844] ^ n[2845];
assign t[2846] = t[2845] ^ n[2846];
assign t[2847] = t[2846] ^ n[2847];
assign t[2848] = t[2847] ^ n[2848];
assign t[2849] = t[2848] ^ n[2849];
assign t[2850] = t[2849] ^ n[2850];
assign t[2851] = t[2850] ^ n[2851];
assign t[2852] = t[2851] ^ n[2852];
assign t[2853] = t[2852] ^ n[2853];
assign t[2854] = t[2853] ^ n[2854];
assign t[2855] = t[2854] ^ n[2855];
assign t[2856] = t[2855] ^ n[2856];
assign t[2857] = t[2856] ^ n[2857];
assign t[2858] = t[2857] ^ n[2858];
assign t[2859] = t[2858] ^ n[2859];
assign t[2860] = t[2859] ^ n[2860];
assign t[2861] = t[2860] ^ n[2861];
assign t[2862] = t[2861] ^ n[2862];
assign t[2863] = t[2862] ^ n[2863];
assign t[2864] = t[2863] ^ n[2864];
assign t[2865] = t[2864] ^ n[2865];
assign t[2866] = t[2865] ^ n[2866];
assign t[2867] = t[2866] ^ n[2867];
assign t[2868] = t[2867] ^ n[2868];
assign t[2869] = t[2868] ^ n[2869];
assign t[2870] = t[2869] ^ n[2870];
assign t[2871] = t[2870] ^ n[2871];
assign t[2872] = t[2871] ^ n[2872];
assign t[2873] = t[2872] ^ n[2873];
assign t[2874] = t[2873] ^ n[2874];
assign t[2875] = t[2874] ^ n[2875];
assign t[2876] = t[2875] ^ n[2876];
assign t[2877] = t[2876] ^ n[2877];
assign t[2878] = t[2877] ^ n[2878];
assign t[2879] = t[2878] ^ n[2879];
assign t[2880] = t[2879] ^ n[2880];
assign t[2881] = t[2880] ^ n[2881];
assign t[2882] = t[2881] ^ n[2882];
assign t[2883] = t[2882] ^ n[2883];
assign t[2884] = t[2883] ^ n[2884];
assign t[2885] = t[2884] ^ n[2885];
assign t[2886] = t[2885] ^ n[2886];
assign t[2887] = t[2886] ^ n[2887];
assign t[2888] = t[2887] ^ n[2888];
assign t[2889] = t[2888] ^ n[2889];
assign t[2890] = t[2889] ^ n[2890];
assign t[2891] = t[2890] ^ n[2891];
assign t[2892] = t[2891] ^ n[2892];
assign t[2893] = t[2892] ^ n[2893];
assign t[2894] = t[2893] ^ n[2894];
assign t[2895] = t[2894] ^ n[2895];
assign t[2896] = t[2895] ^ n[2896];
assign t[2897] = t[2896] ^ n[2897];
assign t[2898] = t[2897] ^ n[2898];
assign t[2899] = t[2898] ^ n[2899];
assign t[2900] = t[2899] ^ n[2900];
assign t[2901] = t[2900] ^ n[2901];
assign t[2902] = t[2901] ^ n[2902];
assign t[2903] = t[2902] ^ n[2903];
assign t[2904] = t[2903] ^ n[2904];
assign t[2905] = t[2904] ^ n[2905];
assign t[2906] = t[2905] ^ n[2906];
assign t[2907] = t[2906] ^ n[2907];
assign t[2908] = t[2907] ^ n[2908];
assign t[2909] = t[2908] ^ n[2909];
assign t[2910] = t[2909] ^ n[2910];
assign t[2911] = t[2910] ^ n[2911];
assign t[2912] = t[2911] ^ n[2912];
assign t[2913] = t[2912] ^ n[2913];
assign t[2914] = t[2913] ^ n[2914];
assign t[2915] = t[2914] ^ n[2915];
assign t[2916] = t[2915] ^ n[2916];
assign t[2917] = t[2916] ^ n[2917];
assign t[2918] = t[2917] ^ n[2918];
assign t[2919] = t[2918] ^ n[2919];
assign t[2920] = t[2919] ^ n[2920];
assign t[2921] = t[2920] ^ n[2921];
assign t[2922] = t[2921] ^ n[2922];
assign t[2923] = t[2922] ^ n[2923];
assign t[2924] = t[2923] ^ n[2924];
assign t[2925] = t[2924] ^ n[2925];
assign t[2926] = t[2925] ^ n[2926];
assign t[2927] = t[2926] ^ n[2927];
assign t[2928] = t[2927] ^ n[2928];
assign t[2929] = t[2928] ^ n[2929];
assign t[2930] = t[2929] ^ n[2930];
assign t[2931] = t[2930] ^ n[2931];
assign t[2932] = t[2931] ^ n[2932];
assign t[2933] = t[2932] ^ n[2933];
assign t[2934] = t[2933] ^ n[2934];
assign t[2935] = t[2934] ^ n[2935];
assign t[2936] = t[2935] ^ n[2936];
assign t[2937] = t[2936] ^ n[2937];
assign t[2938] = t[2937] ^ n[2938];
assign t[2939] = t[2938] ^ n[2939];
assign t[2940] = t[2939] ^ n[2940];
assign t[2941] = t[2940] ^ n[2941];
assign t[2942] = t[2941] ^ n[2942];
assign t[2943] = t[2942] ^ n[2943];
assign t[2944] = t[2943] ^ n[2944];
assign t[2945] = t[2944] ^ n[2945];
assign t[2946] = t[2945] ^ n[2946];
assign t[2947] = t[2946] ^ n[2947];
assign t[2948] = t[2947] ^ n[2948];
assign t[2949] = t[2948] ^ n[2949];
assign t[2950] = t[2949] ^ n[2950];
assign t[2951] = t[2950] ^ n[2951];
assign t[2952] = t[2951] ^ n[2952];
assign t[2953] = t[2952] ^ n[2953];
assign t[2954] = t[2953] ^ n[2954];
assign t[2955] = t[2954] ^ n[2955];
assign t[2956] = t[2955] ^ n[2956];
assign t[2957] = t[2956] ^ n[2957];
assign t[2958] = t[2957] ^ n[2958];
assign t[2959] = t[2958] ^ n[2959];
assign t[2960] = t[2959] ^ n[2960];
assign t[2961] = t[2960] ^ n[2961];
assign t[2962] = t[2961] ^ n[2962];
assign t[2963] = t[2962] ^ n[2963];
assign t[2964] = t[2963] ^ n[2964];
assign t[2965] = t[2964] ^ n[2965];
assign t[2966] = t[2965] ^ n[2966];
assign t[2967] = t[2966] ^ n[2967];
assign t[2968] = t[2967] ^ n[2968];
assign t[2969] = t[2968] ^ n[2969];
assign t[2970] = t[2969] ^ n[2970];
assign t[2971] = t[2970] ^ n[2971];
assign t[2972] = t[2971] ^ n[2972];
assign t[2973] = t[2972] ^ n[2973];
assign t[2974] = t[2973] ^ n[2974];
assign t[2975] = t[2974] ^ n[2975];
assign t[2976] = t[2975] ^ n[2976];
assign t[2977] = t[2976] ^ n[2977];
assign t[2978] = t[2977] ^ n[2978];
assign t[2979] = t[2978] ^ n[2979];
assign t[2980] = t[2979] ^ n[2980];
assign t[2981] = t[2980] ^ n[2981];
assign t[2982] = t[2981] ^ n[2982];
assign t[2983] = t[2982] ^ n[2983];
assign t[2984] = t[2983] ^ n[2984];
assign t[2985] = t[2984] ^ n[2985];
assign t[2986] = t[2985] ^ n[2986];
assign t[2987] = t[2986] ^ n[2987];
assign t[2988] = t[2987] ^ n[2988];
assign t[2989] = t[2988] ^ n[2989];
assign t[2990] = t[2989] ^ n[2990];
assign t[2991] = t[2990] ^ n[2991];
assign t[2992] = t[2991] ^ n[2992];
assign t[2993] = t[2992] ^ n[2993];
assign t[2994] = t[2993] ^ n[2994];
assign t[2995] = t[2994] ^ n[2995];
assign t[2996] = t[2995] ^ n[2996];
assign t[2997] = t[2996] ^ n[2997];
assign t[2998] = t[2997] ^ n[2998];
assign t[2999] = t[2998] ^ n[2999];
assign t[3000] = t[2999] ^ n[3000];
assign t[3001] = t[3000] ^ n[3001];
assign t[3002] = t[3001] ^ n[3002];
assign t[3003] = t[3002] ^ n[3003];
assign t[3004] = t[3003] ^ n[3004];
assign t[3005] = t[3004] ^ n[3005];
assign t[3006] = t[3005] ^ n[3006];
assign t[3007] = t[3006] ^ n[3007];
assign t[3008] = t[3007] ^ n[3008];
assign t[3009] = t[3008] ^ n[3009];
assign t[3010] = t[3009] ^ n[3010];
assign t[3011] = t[3010] ^ n[3011];
assign t[3012] = t[3011] ^ n[3012];
assign t[3013] = t[3012] ^ n[3013];
assign t[3014] = t[3013] ^ n[3014];
assign t[3015] = t[3014] ^ n[3015];
assign t[3016] = t[3015] ^ n[3016];
assign t[3017] = t[3016] ^ n[3017];
assign t[3018] = t[3017] ^ n[3018];
assign t[3019] = t[3018] ^ n[3019];
assign t[3020] = t[3019] ^ n[3020];
assign t[3021] = t[3020] ^ n[3021];
assign t[3022] = t[3021] ^ n[3022];
assign t[3023] = t[3022] ^ n[3023];
assign t[3024] = t[3023] ^ n[3024];
assign t[3025] = t[3024] ^ n[3025];
assign t[3026] = t[3025] ^ n[3026];
assign t[3027] = t[3026] ^ n[3027];
assign t[3028] = t[3027] ^ n[3028];
assign t[3029] = t[3028] ^ n[3029];
assign t[3030] = t[3029] ^ n[3030];
assign t[3031] = t[3030] ^ n[3031];
assign t[3032] = t[3031] ^ n[3032];
assign t[3033] = t[3032] ^ n[3033];
assign t[3034] = t[3033] ^ n[3034];
assign t[3035] = t[3034] ^ n[3035];
assign t[3036] = t[3035] ^ n[3036];
assign t[3037] = t[3036] ^ n[3037];
assign t[3038] = t[3037] ^ n[3038];
assign t[3039] = t[3038] ^ n[3039];
assign t[3040] = t[3039] ^ n[3040];
assign t[3041] = t[3040] ^ n[3041];
assign t[3042] = t[3041] ^ n[3042];
assign t[3043] = t[3042] ^ n[3043];
assign t[3044] = t[3043] ^ n[3044];
assign t[3045] = t[3044] ^ n[3045];
assign t[3046] = t[3045] ^ n[3046];
assign t[3047] = t[3046] ^ n[3047];
assign t[3048] = t[3047] ^ n[3048];
assign t[3049] = t[3048] ^ n[3049];
assign t[3050] = t[3049] ^ n[3050];
assign t[3051] = t[3050] ^ n[3051];
assign t[3052] = t[3051] ^ n[3052];
assign t[3053] = t[3052] ^ n[3053];
assign t[3054] = t[3053] ^ n[3054];
assign t[3055] = t[3054] ^ n[3055];
assign t[3056] = t[3055] ^ n[3056];
assign t[3057] = t[3056] ^ n[3057];
assign t[3058] = t[3057] ^ n[3058];
assign t[3059] = t[3058] ^ n[3059];
assign t[3060] = t[3059] ^ n[3060];
assign t[3061] = t[3060] ^ n[3061];
assign t[3062] = t[3061] ^ n[3062];
assign t[3063] = t[3062] ^ n[3063];
assign t[3064] = t[3063] ^ n[3064];
assign t[3065] = t[3064] ^ n[3065];
assign t[3066] = t[3065] ^ n[3066];
assign t[3067] = t[3066] ^ n[3067];
assign t[3068] = t[3067] ^ n[3068];
assign t[3069] = t[3068] ^ n[3069];
assign t[3070] = t[3069] ^ n[3070];
assign t[3071] = t[3070] ^ n[3071];
assign t[3072] = t[3071] ^ n[3072];
assign t[3073] = t[3072] ^ n[3073];
assign t[3074] = t[3073] ^ n[3074];
assign t[3075] = t[3074] ^ n[3075];
assign t[3076] = t[3075] ^ n[3076];
assign t[3077] = t[3076] ^ n[3077];
assign t[3078] = t[3077] ^ n[3078];
assign t[3079] = t[3078] ^ n[3079];
assign t[3080] = t[3079] ^ n[3080];
assign t[3081] = t[3080] ^ n[3081];
assign t[3082] = t[3081] ^ n[3082];
assign t[3083] = t[3082] ^ n[3083];
assign t[3084] = t[3083] ^ n[3084];
assign t[3085] = t[3084] ^ n[3085];
assign t[3086] = t[3085] ^ n[3086];
assign t[3087] = t[3086] ^ n[3087];
assign t[3088] = t[3087] ^ n[3088];
assign t[3089] = t[3088] ^ n[3089];
assign t[3090] = t[3089] ^ n[3090];
assign t[3091] = t[3090] ^ n[3091];
assign t[3092] = t[3091] ^ n[3092];
assign t[3093] = t[3092] ^ n[3093];
assign t[3094] = t[3093] ^ n[3094];
assign t[3095] = t[3094] ^ n[3095];
assign t[3096] = t[3095] ^ n[3096];
assign t[3097] = t[3096] ^ n[3097];
assign t[3098] = t[3097] ^ n[3098];
assign t[3099] = t[3098] ^ n[3099];
assign t[3100] = t[3099] ^ n[3100];
assign t[3101] = t[3100] ^ n[3101];
assign t[3102] = t[3101] ^ n[3102];
assign t[3103] = t[3102] ^ n[3103];
assign t[3104] = t[3103] ^ n[3104];
assign t[3105] = t[3104] ^ n[3105];
assign t[3106] = t[3105] ^ n[3106];
assign t[3107] = t[3106] ^ n[3107];
assign t[3108] = t[3107] ^ n[3108];
assign t[3109] = t[3108] ^ n[3109];
assign t[3110] = t[3109] ^ n[3110];
assign t[3111] = t[3110] ^ n[3111];
assign t[3112] = t[3111] ^ n[3112];
assign t[3113] = t[3112] ^ n[3113];
assign t[3114] = t[3113] ^ n[3114];
assign t[3115] = t[3114] ^ n[3115];
assign t[3116] = t[3115] ^ n[3116];
assign t[3117] = t[3116] ^ n[3117];
assign t[3118] = t[3117] ^ n[3118];
assign t[3119] = t[3118] ^ n[3119];
assign t[3120] = t[3119] ^ n[3120];
assign t[3121] = t[3120] ^ n[3121];
assign t[3122] = t[3121] ^ n[3122];
assign t[3123] = t[3122] ^ n[3123];
assign t[3124] = t[3123] ^ n[3124];
assign t[3125] = t[3124] ^ n[3125];
assign t[3126] = t[3125] ^ n[3126];
assign t[3127] = t[3126] ^ n[3127];
assign t[3128] = t[3127] ^ n[3128];
assign t[3129] = t[3128] ^ n[3129];
assign t[3130] = t[3129] ^ n[3130];
assign t[3131] = t[3130] ^ n[3131];
assign t[3132] = t[3131] ^ n[3132];
assign t[3133] = t[3132] ^ n[3133];
assign t[3134] = t[3133] ^ n[3134];
assign t[3135] = t[3134] ^ n[3135];
assign t[3136] = t[3135] ^ n[3136];
assign t[3137] = t[3136] ^ n[3137];
assign t[3138] = t[3137] ^ n[3138];
assign t[3139] = t[3138] ^ n[3139];
assign t[3140] = t[3139] ^ n[3140];
assign t[3141] = t[3140] ^ n[3141];
assign t[3142] = t[3141] ^ n[3142];
assign t[3143] = t[3142] ^ n[3143];
assign t[3144] = t[3143] ^ n[3144];
assign t[3145] = t[3144] ^ n[3145];
assign t[3146] = t[3145] ^ n[3146];
assign t[3147] = t[3146] ^ n[3147];
assign t[3148] = t[3147] ^ n[3148];
assign t[3149] = t[3148] ^ n[3149];
assign t[3150] = t[3149] ^ n[3150];
assign t[3151] = t[3150] ^ n[3151];
assign t[3152] = t[3151] ^ n[3152];
assign t[3153] = t[3152] ^ n[3153];
assign t[3154] = t[3153] ^ n[3154];
assign t[3155] = t[3154] ^ n[3155];
assign t[3156] = t[3155] ^ n[3156];
assign t[3157] = t[3156] ^ n[3157];
assign t[3158] = t[3157] ^ n[3158];
assign t[3159] = t[3158] ^ n[3159];
assign t[3160] = t[3159] ^ n[3160];
assign t[3161] = t[3160] ^ n[3161];
assign t[3162] = t[3161] ^ n[3162];
assign t[3163] = t[3162] ^ n[3163];
assign t[3164] = t[3163] ^ n[3164];
assign t[3165] = t[3164] ^ n[3165];
assign t[3166] = t[3165] ^ n[3166];
assign t[3167] = t[3166] ^ n[3167];
assign t[3168] = t[3167] ^ n[3168];
assign t[3169] = t[3168] ^ n[3169];
assign t[3170] = t[3169] ^ n[3170];
assign t[3171] = t[3170] ^ n[3171];
assign t[3172] = t[3171] ^ n[3172];
assign t[3173] = t[3172] ^ n[3173];
assign t[3174] = t[3173] ^ n[3174];
assign t[3175] = t[3174] ^ n[3175];
assign t[3176] = t[3175] ^ n[3176];
assign t[3177] = t[3176] ^ n[3177];
assign t[3178] = t[3177] ^ n[3178];
assign t[3179] = t[3178] ^ n[3179];
assign t[3180] = t[3179] ^ n[3180];
assign t[3181] = t[3180] ^ n[3181];
assign t[3182] = t[3181] ^ n[3182];
assign t[3183] = t[3182] ^ n[3183];
assign t[3184] = t[3183] ^ n[3184];
assign t[3185] = t[3184] ^ n[3185];
assign t[3186] = t[3185] ^ n[3186];
assign t[3187] = t[3186] ^ n[3187];
assign t[3188] = t[3187] ^ n[3188];
assign t[3189] = t[3188] ^ n[3189];
assign t[3190] = t[3189] ^ n[3190];
assign t[3191] = t[3190] ^ n[3191];
assign t[3192] = t[3191] ^ n[3192];
assign t[3193] = t[3192] ^ n[3193];
assign t[3194] = t[3193] ^ n[3194];
assign t[3195] = t[3194] ^ n[3195];
assign t[3196] = t[3195] ^ n[3196];
assign t[3197] = t[3196] ^ n[3197];
assign t[3198] = t[3197] ^ n[3198];
assign t[3199] = t[3198] ^ n[3199];
assign t[3200] = t[3199] ^ n[3200];
assign t[3201] = t[3200] ^ n[3201];
assign t[3202] = t[3201] ^ n[3202];
assign t[3203] = t[3202] ^ n[3203];
assign t[3204] = t[3203] ^ n[3204];
assign t[3205] = t[3204] ^ n[3205];
assign t[3206] = t[3205] ^ n[3206];
assign t[3207] = t[3206] ^ n[3207];
assign t[3208] = t[3207] ^ n[3208];
assign t[3209] = t[3208] ^ n[3209];
assign t[3210] = t[3209] ^ n[3210];
assign t[3211] = t[3210] ^ n[3211];
assign t[3212] = t[3211] ^ n[3212];
assign t[3213] = t[3212] ^ n[3213];
assign t[3214] = t[3213] ^ n[3214];
assign t[3215] = t[3214] ^ n[3215];
assign t[3216] = t[3215] ^ n[3216];
assign t[3217] = t[3216] ^ n[3217];
assign t[3218] = t[3217] ^ n[3218];
assign t[3219] = t[3218] ^ n[3219];
assign t[3220] = t[3219] ^ n[3220];
assign t[3221] = t[3220] ^ n[3221];
assign t[3222] = t[3221] ^ n[3222];
assign t[3223] = t[3222] ^ n[3223];
assign t[3224] = t[3223] ^ n[3224];
assign t[3225] = t[3224] ^ n[3225];
assign t[3226] = t[3225] ^ n[3226];
assign t[3227] = t[3226] ^ n[3227];
assign t[3228] = t[3227] ^ n[3228];
assign t[3229] = t[3228] ^ n[3229];
assign t[3230] = t[3229] ^ n[3230];
assign t[3231] = t[3230] ^ n[3231];
assign t[3232] = t[3231] ^ n[3232];
assign t[3233] = t[3232] ^ n[3233];
assign t[3234] = t[3233] ^ n[3234];
assign t[3235] = t[3234] ^ n[3235];
assign t[3236] = t[3235] ^ n[3236];
assign t[3237] = t[3236] ^ n[3237];
assign t[3238] = t[3237] ^ n[3238];
assign t[3239] = t[3238] ^ n[3239];
assign t[3240] = t[3239] ^ n[3240];
assign t[3241] = t[3240] ^ n[3241];
assign t[3242] = t[3241] ^ n[3242];
assign t[3243] = t[3242] ^ n[3243];
assign t[3244] = t[3243] ^ n[3244];
assign t[3245] = t[3244] ^ n[3245];
assign t[3246] = t[3245] ^ n[3246];
assign t[3247] = t[3246] ^ n[3247];
assign t[3248] = t[3247] ^ n[3248];
assign t[3249] = t[3248] ^ n[3249];
assign t[3250] = t[3249] ^ n[3250];
assign t[3251] = t[3250] ^ n[3251];
assign t[3252] = t[3251] ^ n[3252];
assign t[3253] = t[3252] ^ n[3253];
assign t[3254] = t[3253] ^ n[3254];
assign t[3255] = t[3254] ^ n[3255];
assign t[3256] = t[3255] ^ n[3256];
assign t[3257] = t[3256] ^ n[3257];
assign t[3258] = t[3257] ^ n[3258];
assign t[3259] = t[3258] ^ n[3259];
assign t[3260] = t[3259] ^ n[3260];
assign t[3261] = t[3260] ^ n[3261];
assign t[3262] = t[3261] ^ n[3262];
assign t[3263] = t[3262] ^ n[3263];
assign t[3264] = t[3263] ^ n[3264];
assign t[3265] = t[3264] ^ n[3265];
assign t[3266] = t[3265] ^ n[3266];
assign t[3267] = t[3266] ^ n[3267];
assign t[3268] = t[3267] ^ n[3268];
assign t[3269] = t[3268] ^ n[3269];
assign t[3270] = t[3269] ^ n[3270];
assign t[3271] = t[3270] ^ n[3271];
assign t[3272] = t[3271] ^ n[3272];
assign t[3273] = t[3272] ^ n[3273];
assign t[3274] = t[3273] ^ n[3274];
assign t[3275] = t[3274] ^ n[3275];
assign t[3276] = t[3275] ^ n[3276];
assign t[3277] = t[3276] ^ n[3277];
assign t[3278] = t[3277] ^ n[3278];
assign t[3279] = t[3278] ^ n[3279];
assign t[3280] = t[3279] ^ n[3280];
assign t[3281] = t[3280] ^ n[3281];
assign t[3282] = t[3281] ^ n[3282];
assign t[3283] = t[3282] ^ n[3283];
assign t[3284] = t[3283] ^ n[3284];
assign t[3285] = t[3284] ^ n[3285];
assign t[3286] = t[3285] ^ n[3286];
assign t[3287] = t[3286] ^ n[3287];
assign t[3288] = t[3287] ^ n[3288];
assign t[3289] = t[3288] ^ n[3289];
assign t[3290] = t[3289] ^ n[3290];
assign t[3291] = t[3290] ^ n[3291];
assign t[3292] = t[3291] ^ n[3292];
assign t[3293] = t[3292] ^ n[3293];
assign t[3294] = t[3293] ^ n[3294];
assign t[3295] = t[3294] ^ n[3295];
assign t[3296] = t[3295] ^ n[3296];
assign t[3297] = t[3296] ^ n[3297];
assign t[3298] = t[3297] ^ n[3298];
assign t[3299] = t[3298] ^ n[3299];
assign t[3300] = t[3299] ^ n[3300];
assign t[3301] = t[3300] ^ n[3301];
assign t[3302] = t[3301] ^ n[3302];
assign t[3303] = t[3302] ^ n[3303];
assign t[3304] = t[3303] ^ n[3304];
assign t[3305] = t[3304] ^ n[3305];
assign t[3306] = t[3305] ^ n[3306];
assign t[3307] = t[3306] ^ n[3307];
assign t[3308] = t[3307] ^ n[3308];
assign t[3309] = t[3308] ^ n[3309];
assign t[3310] = t[3309] ^ n[3310];
assign t[3311] = t[3310] ^ n[3311];
assign t[3312] = t[3311] ^ n[3312];
assign t[3313] = t[3312] ^ n[3313];
assign t[3314] = t[3313] ^ n[3314];
assign t[3315] = t[3314] ^ n[3315];
assign t[3316] = t[3315] ^ n[3316];
assign t[3317] = t[3316] ^ n[3317];
assign t[3318] = t[3317] ^ n[3318];
assign t[3319] = t[3318] ^ n[3319];
assign t[3320] = t[3319] ^ n[3320];
assign t[3321] = t[3320] ^ n[3321];
assign t[3322] = t[3321] ^ n[3322];
assign t[3323] = t[3322] ^ n[3323];
assign t[3324] = t[3323] ^ n[3324];
assign t[3325] = t[3324] ^ n[3325];
assign t[3326] = t[3325] ^ n[3326];
assign t[3327] = t[3326] ^ n[3327];
assign t[3328] = t[3327] ^ n[3328];
assign t[3329] = t[3328] ^ n[3329];
assign t[3330] = t[3329] ^ n[3330];
assign t[3331] = t[3330] ^ n[3331];
assign t[3332] = t[3331] ^ n[3332];
assign t[3333] = t[3332] ^ n[3333];
assign t[3334] = t[3333] ^ n[3334];
assign t[3335] = t[3334] ^ n[3335];
assign t[3336] = t[3335] ^ n[3336];
assign t[3337] = t[3336] ^ n[3337];
assign t[3338] = t[3337] ^ n[3338];
assign t[3339] = t[3338] ^ n[3339];
assign t[3340] = t[3339] ^ n[3340];
assign t[3341] = t[3340] ^ n[3341];
assign t[3342] = t[3341] ^ n[3342];
assign t[3343] = t[3342] ^ n[3343];
assign t[3344] = t[3343] ^ n[3344];
assign t[3345] = t[3344] ^ n[3345];
assign t[3346] = t[3345] ^ n[3346];
assign t[3347] = t[3346] ^ n[3347];
assign t[3348] = t[3347] ^ n[3348];
assign t[3349] = t[3348] ^ n[3349];
assign t[3350] = t[3349] ^ n[3350];
assign t[3351] = t[3350] ^ n[3351];
assign t[3352] = t[3351] ^ n[3352];
assign t[3353] = t[3352] ^ n[3353];
assign t[3354] = t[3353] ^ n[3354];
assign t[3355] = t[3354] ^ n[3355];
assign t[3356] = t[3355] ^ n[3356];
assign t[3357] = t[3356] ^ n[3357];
assign t[3358] = t[3357] ^ n[3358];
assign t[3359] = t[3358] ^ n[3359];
assign t[3360] = t[3359] ^ n[3360];
assign t[3361] = t[3360] ^ n[3361];
assign t[3362] = t[3361] ^ n[3362];
assign t[3363] = t[3362] ^ n[3363];
assign t[3364] = t[3363] ^ n[3364];
assign t[3365] = t[3364] ^ n[3365];
assign t[3366] = t[3365] ^ n[3366];
assign t[3367] = t[3366] ^ n[3367];
assign t[3368] = t[3367] ^ n[3368];
assign t[3369] = t[3368] ^ n[3369];
assign t[3370] = t[3369] ^ n[3370];
assign t[3371] = t[3370] ^ n[3371];
assign t[3372] = t[3371] ^ n[3372];
assign t[3373] = t[3372] ^ n[3373];
assign t[3374] = t[3373] ^ n[3374];
assign t[3375] = t[3374] ^ n[3375];
assign t[3376] = t[3375] ^ n[3376];
assign t[3377] = t[3376] ^ n[3377];
assign t[3378] = t[3377] ^ n[3378];
assign t[3379] = t[3378] ^ n[3379];
assign t[3380] = t[3379] ^ n[3380];
assign t[3381] = t[3380] ^ n[3381];
assign t[3382] = t[3381] ^ n[3382];
assign t[3383] = t[3382] ^ n[3383];
assign t[3384] = t[3383] ^ n[3384];
assign t[3385] = t[3384] ^ n[3385];
assign t[3386] = t[3385] ^ n[3386];
assign t[3387] = t[3386] ^ n[3387];
assign t[3388] = t[3387] ^ n[3388];
assign t[3389] = t[3388] ^ n[3389];
assign t[3390] = t[3389] ^ n[3390];
assign t[3391] = t[3390] ^ n[3391];
assign t[3392] = t[3391] ^ n[3392];
assign t[3393] = t[3392] ^ n[3393];
assign t[3394] = t[3393] ^ n[3394];
assign t[3395] = t[3394] ^ n[3395];
assign t[3396] = t[3395] ^ n[3396];
assign t[3397] = t[3396] ^ n[3397];
assign t[3398] = t[3397] ^ n[3398];
assign t[3399] = t[3398] ^ n[3399];
assign t[3400] = t[3399] ^ n[3400];
assign t[3401] = t[3400] ^ n[3401];
assign t[3402] = t[3401] ^ n[3402];
assign t[3403] = t[3402] ^ n[3403];
assign t[3404] = t[3403] ^ n[3404];
assign t[3405] = t[3404] ^ n[3405];
assign t[3406] = t[3405] ^ n[3406];
assign t[3407] = t[3406] ^ n[3407];
assign t[3408] = t[3407] ^ n[3408];
assign t[3409] = t[3408] ^ n[3409];
assign t[3410] = t[3409] ^ n[3410];
assign t[3411] = t[3410] ^ n[3411];
assign t[3412] = t[3411] ^ n[3412];
assign t[3413] = t[3412] ^ n[3413];
assign t[3414] = t[3413] ^ n[3414];
assign t[3415] = t[3414] ^ n[3415];
assign t[3416] = t[3415] ^ n[3416];
assign t[3417] = t[3416] ^ n[3417];
assign t[3418] = t[3417] ^ n[3418];
assign t[3419] = t[3418] ^ n[3419];
assign t[3420] = t[3419] ^ n[3420];
assign t[3421] = t[3420] ^ n[3421];
assign t[3422] = t[3421] ^ n[3422];
assign t[3423] = t[3422] ^ n[3423];
assign t[3424] = t[3423] ^ n[3424];
assign t[3425] = t[3424] ^ n[3425];
assign t[3426] = t[3425] ^ n[3426];
assign t[3427] = t[3426] ^ n[3427];
assign t[3428] = t[3427] ^ n[3428];
assign t[3429] = t[3428] ^ n[3429];
assign t[3430] = t[3429] ^ n[3430];
assign t[3431] = t[3430] ^ n[3431];
assign t[3432] = t[3431] ^ n[3432];
assign t[3433] = t[3432] ^ n[3433];
assign t[3434] = t[3433] ^ n[3434];
assign t[3435] = t[3434] ^ n[3435];
assign t[3436] = t[3435] ^ n[3436];
assign t[3437] = t[3436] ^ n[3437];
assign t[3438] = t[3437] ^ n[3438];
assign t[3439] = t[3438] ^ n[3439];
assign t[3440] = t[3439] ^ n[3440];
assign t[3441] = t[3440] ^ n[3441];
assign t[3442] = t[3441] ^ n[3442];
assign t[3443] = t[3442] ^ n[3443];
assign t[3444] = t[3443] ^ n[3444];
assign t[3445] = t[3444] ^ n[3445];
assign t[3446] = t[3445] ^ n[3446];
assign t[3447] = t[3446] ^ n[3447];
assign t[3448] = t[3447] ^ n[3448];
assign t[3449] = t[3448] ^ n[3449];
assign t[3450] = t[3449] ^ n[3450];
assign t[3451] = t[3450] ^ n[3451];
assign t[3452] = t[3451] ^ n[3452];
assign t[3453] = t[3452] ^ n[3453];
assign t[3454] = t[3453] ^ n[3454];
assign t[3455] = t[3454] ^ n[3455];
assign t[3456] = t[3455] ^ n[3456];
assign t[3457] = t[3456] ^ n[3457];
assign t[3458] = t[3457] ^ n[3458];
assign t[3459] = t[3458] ^ n[3459];
assign t[3460] = t[3459] ^ n[3460];
assign t[3461] = t[3460] ^ n[3461];
assign t[3462] = t[3461] ^ n[3462];
assign t[3463] = t[3462] ^ n[3463];
assign t[3464] = t[3463] ^ n[3464];
assign t[3465] = t[3464] ^ n[3465];
assign t[3466] = t[3465] ^ n[3466];
assign t[3467] = t[3466] ^ n[3467];
assign t[3468] = t[3467] ^ n[3468];
assign t[3469] = t[3468] ^ n[3469];
assign t[3470] = t[3469] ^ n[3470];
assign t[3471] = t[3470] ^ n[3471];
assign t[3472] = t[3471] ^ n[3472];
assign t[3473] = t[3472] ^ n[3473];
assign t[3474] = t[3473] ^ n[3474];
assign t[3475] = t[3474] ^ n[3475];
assign t[3476] = t[3475] ^ n[3476];
assign t[3477] = t[3476] ^ n[3477];
assign t[3478] = t[3477] ^ n[3478];
assign t[3479] = t[3478] ^ n[3479];
assign t[3480] = t[3479] ^ n[3480];
assign t[3481] = t[3480] ^ n[3481];
assign t[3482] = t[3481] ^ n[3482];
assign t[3483] = t[3482] ^ n[3483];
assign t[3484] = t[3483] ^ n[3484];
assign t[3485] = t[3484] ^ n[3485];
assign t[3486] = t[3485] ^ n[3486];
assign t[3487] = t[3486] ^ n[3487];
assign t[3488] = t[3487] ^ n[3488];
assign t[3489] = t[3488] ^ n[3489];
assign t[3490] = t[3489] ^ n[3490];
assign t[3491] = t[3490] ^ n[3491];
assign t[3492] = t[3491] ^ n[3492];
assign t[3493] = t[3492] ^ n[3493];
assign t[3494] = t[3493] ^ n[3494];
assign t[3495] = t[3494] ^ n[3495];
assign t[3496] = t[3495] ^ n[3496];
assign t[3497] = t[3496] ^ n[3497];
assign t[3498] = t[3497] ^ n[3498];
assign t[3499] = t[3498] ^ n[3499];
assign t[3500] = t[3499] ^ n[3500];
assign t[3501] = t[3500] ^ n[3501];
assign t[3502] = t[3501] ^ n[3502];
assign t[3503] = t[3502] ^ n[3503];
assign t[3504] = t[3503] ^ n[3504];
assign t[3505] = t[3504] ^ n[3505];
assign t[3506] = t[3505] ^ n[3506];
assign t[3507] = t[3506] ^ n[3507];
assign t[3508] = t[3507] ^ n[3508];
assign t[3509] = t[3508] ^ n[3509];
assign t[3510] = t[3509] ^ n[3510];
assign t[3511] = t[3510] ^ n[3511];
assign t[3512] = t[3511] ^ n[3512];
assign t[3513] = t[3512] ^ n[3513];
assign t[3514] = t[3513] ^ n[3514];
assign t[3515] = t[3514] ^ n[3515];
assign t[3516] = t[3515] ^ n[3516];
assign t[3517] = t[3516] ^ n[3517];
assign t[3518] = t[3517] ^ n[3518];
assign t[3519] = t[3518] ^ n[3519];
assign t[3520] = t[3519] ^ n[3520];
assign t[3521] = t[3520] ^ n[3521];
assign t[3522] = t[3521] ^ n[3522];
assign t[3523] = t[3522] ^ n[3523];
assign t[3524] = t[3523] ^ n[3524];
assign t[3525] = t[3524] ^ n[3525];
assign t[3526] = t[3525] ^ n[3526];
assign t[3527] = t[3526] ^ n[3527];
assign t[3528] = t[3527] ^ n[3528];
assign t[3529] = t[3528] ^ n[3529];
assign t[3530] = t[3529] ^ n[3530];
assign t[3531] = t[3530] ^ n[3531];
assign t[3532] = t[3531] ^ n[3532];
assign t[3533] = t[3532] ^ n[3533];
assign t[3534] = t[3533] ^ n[3534];
assign t[3535] = t[3534] ^ n[3535];
assign t[3536] = t[3535] ^ n[3536];
assign t[3537] = t[3536] ^ n[3537];
assign t[3538] = t[3537] ^ n[3538];
assign t[3539] = t[3538] ^ n[3539];
assign t[3540] = t[3539] ^ n[3540];
assign t[3541] = t[3540] ^ n[3541];
assign t[3542] = t[3541] ^ n[3542];
assign t[3543] = t[3542] ^ n[3543];
assign t[3544] = t[3543] ^ n[3544];
assign t[3545] = t[3544] ^ n[3545];
assign t[3546] = t[3545] ^ n[3546];
assign t[3547] = t[3546] ^ n[3547];
assign t[3548] = t[3547] ^ n[3548];
assign t[3549] = t[3548] ^ n[3549];
assign t[3550] = t[3549] ^ n[3550];
assign t[3551] = t[3550] ^ n[3551];
assign t[3552] = t[3551] ^ n[3552];
assign t[3553] = t[3552] ^ n[3553];
assign t[3554] = t[3553] ^ n[3554];
assign t[3555] = t[3554] ^ n[3555];
assign t[3556] = t[3555] ^ n[3556];
assign t[3557] = t[3556] ^ n[3557];
assign t[3558] = t[3557] ^ n[3558];
assign t[3559] = t[3558] ^ n[3559];
assign t[3560] = t[3559] ^ n[3560];
assign t[3561] = t[3560] ^ n[3561];
assign t[3562] = t[3561] ^ n[3562];
assign t[3563] = t[3562] ^ n[3563];
assign t[3564] = t[3563] ^ n[3564];
assign t[3565] = t[3564] ^ n[3565];
assign t[3566] = t[3565] ^ n[3566];
assign t[3567] = t[3566] ^ n[3567];
assign t[3568] = t[3567] ^ n[3568];
assign t[3569] = t[3568] ^ n[3569];
assign t[3570] = t[3569] ^ n[3570];
assign t[3571] = t[3570] ^ n[3571];
assign t[3572] = t[3571] ^ n[3572];
assign t[3573] = t[3572] ^ n[3573];
assign t[3574] = t[3573] ^ n[3574];
assign t[3575] = t[3574] ^ n[3575];
assign t[3576] = t[3575] ^ n[3576];
assign t[3577] = t[3576] ^ n[3577];
assign t[3578] = t[3577] ^ n[3578];
assign t[3579] = t[3578] ^ n[3579];
assign t[3580] = t[3579] ^ n[3580];
assign t[3581] = t[3580] ^ n[3581];
assign t[3582] = t[3581] ^ n[3582];
assign t[3583] = t[3582] ^ n[3583];
assign t[3584] = t[3583] ^ n[3584];
assign t[3585] = t[3584] ^ n[3585];
assign t[3586] = t[3585] ^ n[3586];
assign t[3587] = t[3586] ^ n[3587];
assign t[3588] = t[3587] ^ n[3588];
assign t[3589] = t[3588] ^ n[3589];
assign t[3590] = t[3589] ^ n[3590];
assign t[3591] = t[3590] ^ n[3591];
assign t[3592] = t[3591] ^ n[3592];
assign t[3593] = t[3592] ^ n[3593];
assign t[3594] = t[3593] ^ n[3594];
assign t[3595] = t[3594] ^ n[3595];
assign t[3596] = t[3595] ^ n[3596];
assign t[3597] = t[3596] ^ n[3597];
assign t[3598] = t[3597] ^ n[3598];
assign t[3599] = t[3598] ^ n[3599];
assign t[3600] = t[3599] ^ n[3600];
assign t[3601] = t[3600] ^ n[3601];
assign t[3602] = t[3601] ^ n[3602];
assign t[3603] = t[3602] ^ n[3603];
assign t[3604] = t[3603] ^ n[3604];
assign t[3605] = t[3604] ^ n[3605];
assign t[3606] = t[3605] ^ n[3606];
assign t[3607] = t[3606] ^ n[3607];
assign t[3608] = t[3607] ^ n[3608];
assign t[3609] = t[3608] ^ n[3609];
assign t[3610] = t[3609] ^ n[3610];
assign t[3611] = t[3610] ^ n[3611];
assign t[3612] = t[3611] ^ n[3612];
assign t[3613] = t[3612] ^ n[3613];
assign t[3614] = t[3613] ^ n[3614];
assign t[3615] = t[3614] ^ n[3615];
assign t[3616] = t[3615] ^ n[3616];
assign t[3617] = t[3616] ^ n[3617];
assign t[3618] = t[3617] ^ n[3618];
assign t[3619] = t[3618] ^ n[3619];
assign t[3620] = t[3619] ^ n[3620];
assign t[3621] = t[3620] ^ n[3621];
assign t[3622] = t[3621] ^ n[3622];
assign t[3623] = t[3622] ^ n[3623];
assign t[3624] = t[3623] ^ n[3624];
assign t[3625] = t[3624] ^ n[3625];
assign t[3626] = t[3625] ^ n[3626];
assign t[3627] = t[3626] ^ n[3627];
assign t[3628] = t[3627] ^ n[3628];
assign t[3629] = t[3628] ^ n[3629];
assign t[3630] = t[3629] ^ n[3630];
assign t[3631] = t[3630] ^ n[3631];
assign t[3632] = t[3631] ^ n[3632];
assign t[3633] = t[3632] ^ n[3633];
assign t[3634] = t[3633] ^ n[3634];
assign t[3635] = t[3634] ^ n[3635];
assign t[3636] = t[3635] ^ n[3636];
assign t[3637] = t[3636] ^ n[3637];
assign t[3638] = t[3637] ^ n[3638];
assign t[3639] = t[3638] ^ n[3639];
assign t[3640] = t[3639] ^ n[3640];
assign t[3641] = t[3640] ^ n[3641];
assign t[3642] = t[3641] ^ n[3642];
assign t[3643] = t[3642] ^ n[3643];
assign t[3644] = t[3643] ^ n[3644];
assign t[3645] = t[3644] ^ n[3645];
assign t[3646] = t[3645] ^ n[3646];
assign t[3647] = t[3646] ^ n[3647];
assign t[3648] = t[3647] ^ n[3648];
assign t[3649] = t[3648] ^ n[3649];
assign t[3650] = t[3649] ^ n[3650];
assign t[3651] = t[3650] ^ n[3651];
assign t[3652] = t[3651] ^ n[3652];
assign t[3653] = t[3652] ^ n[3653];
assign t[3654] = t[3653] ^ n[3654];
assign t[3655] = t[3654] ^ n[3655];
assign t[3656] = t[3655] ^ n[3656];
assign t[3657] = t[3656] ^ n[3657];
assign t[3658] = t[3657] ^ n[3658];
assign t[3659] = t[3658] ^ n[3659];
assign t[3660] = t[3659] ^ n[3660];
assign t[3661] = t[3660] ^ n[3661];
assign t[3662] = t[3661] ^ n[3662];
assign t[3663] = t[3662] ^ n[3663];
assign t[3664] = t[3663] ^ n[3664];
assign t[3665] = t[3664] ^ n[3665];
assign t[3666] = t[3665] ^ n[3666];
assign t[3667] = t[3666] ^ n[3667];
assign t[3668] = t[3667] ^ n[3668];
assign t[3669] = t[3668] ^ n[3669];
assign t[3670] = t[3669] ^ n[3670];
assign t[3671] = t[3670] ^ n[3671];
assign t[3672] = t[3671] ^ n[3672];
assign t[3673] = t[3672] ^ n[3673];
assign t[3674] = t[3673] ^ n[3674];
assign t[3675] = t[3674] ^ n[3675];
assign t[3676] = t[3675] ^ n[3676];
assign t[3677] = t[3676] ^ n[3677];
assign t[3678] = t[3677] ^ n[3678];
assign t[3679] = t[3678] ^ n[3679];
assign t[3680] = t[3679] ^ n[3680];
assign t[3681] = t[3680] ^ n[3681];
assign t[3682] = t[3681] ^ n[3682];
assign t[3683] = t[3682] ^ n[3683];
assign t[3684] = t[3683] ^ n[3684];
assign t[3685] = t[3684] ^ n[3685];
assign t[3686] = t[3685] ^ n[3686];
assign t[3687] = t[3686] ^ n[3687];
assign t[3688] = t[3687] ^ n[3688];
assign t[3689] = t[3688] ^ n[3689];
assign t[3690] = t[3689] ^ n[3690];
assign t[3691] = t[3690] ^ n[3691];
assign t[3692] = t[3691] ^ n[3692];
assign t[3693] = t[3692] ^ n[3693];
assign t[3694] = t[3693] ^ n[3694];
assign t[3695] = t[3694] ^ n[3695];
assign t[3696] = t[3695] ^ n[3696];
assign t[3697] = t[3696] ^ n[3697];
assign t[3698] = t[3697] ^ n[3698];
assign t[3699] = t[3698] ^ n[3699];
assign t[3700] = t[3699] ^ n[3700];
assign t[3701] = t[3700] ^ n[3701];
assign t[3702] = t[3701] ^ n[3702];
assign t[3703] = t[3702] ^ n[3703];
assign t[3704] = t[3703] ^ n[3704];
assign t[3705] = t[3704] ^ n[3705];
assign t[3706] = t[3705] ^ n[3706];
assign t[3707] = t[3706] ^ n[3707];
assign t[3708] = t[3707] ^ n[3708];
assign t[3709] = t[3708] ^ n[3709];
assign t[3710] = t[3709] ^ n[3710];
assign t[3711] = t[3710] ^ n[3711];
assign t[3712] = t[3711] ^ n[3712];
assign t[3713] = t[3712] ^ n[3713];
assign t[3714] = t[3713] ^ n[3714];
assign t[3715] = t[3714] ^ n[3715];
assign t[3716] = t[3715] ^ n[3716];
assign t[3717] = t[3716] ^ n[3717];
assign t[3718] = t[3717] ^ n[3718];
assign t[3719] = t[3718] ^ n[3719];
assign t[3720] = t[3719] ^ n[3720];
assign t[3721] = t[3720] ^ n[3721];
assign t[3722] = t[3721] ^ n[3722];
assign t[3723] = t[3722] ^ n[3723];
assign t[3724] = t[3723] ^ n[3724];
assign t[3725] = t[3724] ^ n[3725];
assign t[3726] = t[3725] ^ n[3726];
assign t[3727] = t[3726] ^ n[3727];
assign t[3728] = t[3727] ^ n[3728];
assign t[3729] = t[3728] ^ n[3729];
assign t[3730] = t[3729] ^ n[3730];
assign t[3731] = t[3730] ^ n[3731];
assign t[3732] = t[3731] ^ n[3732];
assign t[3733] = t[3732] ^ n[3733];
assign t[3734] = t[3733] ^ n[3734];
assign t[3735] = t[3734] ^ n[3735];
assign t[3736] = t[3735] ^ n[3736];
assign t[3737] = t[3736] ^ n[3737];
assign t[3738] = t[3737] ^ n[3738];
assign t[3739] = t[3738] ^ n[3739];
assign t[3740] = t[3739] ^ n[3740];
assign t[3741] = t[3740] ^ n[3741];
assign t[3742] = t[3741] ^ n[3742];
assign t[3743] = t[3742] ^ n[3743];
assign t[3744] = t[3743] ^ n[3744];
assign t[3745] = t[3744] ^ n[3745];
assign t[3746] = t[3745] ^ n[3746];
assign t[3747] = t[3746] ^ n[3747];
assign t[3748] = t[3747] ^ n[3748];
assign t[3749] = t[3748] ^ n[3749];
assign t[3750] = t[3749] ^ n[3750];
assign t[3751] = t[3750] ^ n[3751];
assign t[3752] = t[3751] ^ n[3752];
assign t[3753] = t[3752] ^ n[3753];
assign t[3754] = t[3753] ^ n[3754];
assign t[3755] = t[3754] ^ n[3755];
assign t[3756] = t[3755] ^ n[3756];
assign t[3757] = t[3756] ^ n[3757];
assign t[3758] = t[3757] ^ n[3758];
assign t[3759] = t[3758] ^ n[3759];
assign t[3760] = t[3759] ^ n[3760];
assign t[3761] = t[3760] ^ n[3761];
assign t[3762] = t[3761] ^ n[3762];
assign t[3763] = t[3762] ^ n[3763];
assign t[3764] = t[3763] ^ n[3764];
assign t[3765] = t[3764] ^ n[3765];
assign t[3766] = t[3765] ^ n[3766];
assign t[3767] = t[3766] ^ n[3767];
assign t[3768] = t[3767] ^ n[3768];
assign t[3769] = t[3768] ^ n[3769];
assign t[3770] = t[3769] ^ n[3770];
assign t[3771] = t[3770] ^ n[3771];
assign t[3772] = t[3771] ^ n[3772];
assign t[3773] = t[3772] ^ n[3773];
assign t[3774] = t[3773] ^ n[3774];
assign t[3775] = t[3774] ^ n[3775];
assign t[3776] = t[3775] ^ n[3776];
assign t[3777] = t[3776] ^ n[3777];
assign t[3778] = t[3777] ^ n[3778];
assign t[3779] = t[3778] ^ n[3779];
assign t[3780] = t[3779] ^ n[3780];
assign t[3781] = t[3780] ^ n[3781];
assign t[3782] = t[3781] ^ n[3782];
assign t[3783] = t[3782] ^ n[3783];
assign t[3784] = t[3783] ^ n[3784];
assign t[3785] = t[3784] ^ n[3785];
assign t[3786] = t[3785] ^ n[3786];
assign t[3787] = t[3786] ^ n[3787];
assign t[3788] = t[3787] ^ n[3788];
assign t[3789] = t[3788] ^ n[3789];
assign t[3790] = t[3789] ^ n[3790];
assign t[3791] = t[3790] ^ n[3791];
assign t[3792] = t[3791] ^ n[3792];
assign t[3793] = t[3792] ^ n[3793];
assign t[3794] = t[3793] ^ n[3794];
assign t[3795] = t[3794] ^ n[3795];
assign t[3796] = t[3795] ^ n[3796];
assign t[3797] = t[3796] ^ n[3797];
assign t[3798] = t[3797] ^ n[3798];
assign t[3799] = t[3798] ^ n[3799];
assign t[3800] = t[3799] ^ n[3800];
assign t[3801] = t[3800] ^ n[3801];
assign t[3802] = t[3801] ^ n[3802];
assign t[3803] = t[3802] ^ n[3803];
assign t[3804] = t[3803] ^ n[3804];
assign t[3805] = t[3804] ^ n[3805];
assign t[3806] = t[3805] ^ n[3806];
assign t[3807] = t[3806] ^ n[3807];
assign t[3808] = t[3807] ^ n[3808];
assign t[3809] = t[3808] ^ n[3809];
assign t[3810] = t[3809] ^ n[3810];
assign t[3811] = t[3810] ^ n[3811];
assign t[3812] = t[3811] ^ n[3812];
assign t[3813] = t[3812] ^ n[3813];
assign t[3814] = t[3813] ^ n[3814];
assign t[3815] = t[3814] ^ n[3815];
assign t[3816] = t[3815] ^ n[3816];
assign t[3817] = t[3816] ^ n[3817];
assign t[3818] = t[3817] ^ n[3818];
assign t[3819] = t[3818] ^ n[3819];
assign t[3820] = t[3819] ^ n[3820];
assign t[3821] = t[3820] ^ n[3821];
assign t[3822] = t[3821] ^ n[3822];
assign t[3823] = t[3822] ^ n[3823];
assign t[3824] = t[3823] ^ n[3824];
assign t[3825] = t[3824] ^ n[3825];
assign t[3826] = t[3825] ^ n[3826];
assign t[3827] = t[3826] ^ n[3827];
assign t[3828] = t[3827] ^ n[3828];
assign t[3829] = t[3828] ^ n[3829];
assign t[3830] = t[3829] ^ n[3830];
assign t[3831] = t[3830] ^ n[3831];
assign t[3832] = t[3831] ^ n[3832];
assign t[3833] = t[3832] ^ n[3833];
assign t[3834] = t[3833] ^ n[3834];
assign t[3835] = t[3834] ^ n[3835];
assign t[3836] = t[3835] ^ n[3836];
assign t[3837] = t[3836] ^ n[3837];
assign t[3838] = t[3837] ^ n[3838];
assign t[3839] = t[3838] ^ n[3839];
assign t[3840] = t[3839] ^ n[3840];
assign t[3841] = t[3840] ^ n[3841];
assign t[3842] = t[3841] ^ n[3842];
assign t[3843] = t[3842] ^ n[3843];
assign t[3844] = t[3843] ^ n[3844];
assign t[3845] = t[3844] ^ n[3845];
assign t[3846] = t[3845] ^ n[3846];
assign t[3847] = t[3846] ^ n[3847];
assign t[3848] = t[3847] ^ n[3848];
assign t[3849] = t[3848] ^ n[3849];
assign t[3850] = t[3849] ^ n[3850];
assign t[3851] = t[3850] ^ n[3851];
assign t[3852] = t[3851] ^ n[3852];
assign t[3853] = t[3852] ^ n[3853];
assign t[3854] = t[3853] ^ n[3854];
assign t[3855] = t[3854] ^ n[3855];
assign t[3856] = t[3855] ^ n[3856];
assign t[3857] = t[3856] ^ n[3857];
assign t[3858] = t[3857] ^ n[3858];
assign t[3859] = t[3858] ^ n[3859];
assign t[3860] = t[3859] ^ n[3860];
assign t[3861] = t[3860] ^ n[3861];
assign t[3862] = t[3861] ^ n[3862];
assign t[3863] = t[3862] ^ n[3863];
assign t[3864] = t[3863] ^ n[3864];
assign t[3865] = t[3864] ^ n[3865];
assign t[3866] = t[3865] ^ n[3866];
assign t[3867] = t[3866] ^ n[3867];
assign t[3868] = t[3867] ^ n[3868];
assign t[3869] = t[3868] ^ n[3869];
assign t[3870] = t[3869] ^ n[3870];
assign t[3871] = t[3870] ^ n[3871];
assign t[3872] = t[3871] ^ n[3872];
assign t[3873] = t[3872] ^ n[3873];
assign t[3874] = t[3873] ^ n[3874];
assign t[3875] = t[3874] ^ n[3875];
assign t[3876] = t[3875] ^ n[3876];
assign t[3877] = t[3876] ^ n[3877];
assign t[3878] = t[3877] ^ n[3878];
assign t[3879] = t[3878] ^ n[3879];
assign t[3880] = t[3879] ^ n[3880];
assign t[3881] = t[3880] ^ n[3881];
assign t[3882] = t[3881] ^ n[3882];
assign t[3883] = t[3882] ^ n[3883];
assign t[3884] = t[3883] ^ n[3884];
assign t[3885] = t[3884] ^ n[3885];
assign t[3886] = t[3885] ^ n[3886];
assign t[3887] = t[3886] ^ n[3887];
assign t[3888] = t[3887] ^ n[3888];
assign t[3889] = t[3888] ^ n[3889];
assign t[3890] = t[3889] ^ n[3890];
assign t[3891] = t[3890] ^ n[3891];
assign t[3892] = t[3891] ^ n[3892];
assign t[3893] = t[3892] ^ n[3893];
assign t[3894] = t[3893] ^ n[3894];
assign t[3895] = t[3894] ^ n[3895];
assign t[3896] = t[3895] ^ n[3896];
assign t[3897] = t[3896] ^ n[3897];
assign t[3898] = t[3897] ^ n[3898];
assign t[3899] = t[3898] ^ n[3899];
assign t[3900] = t[3899] ^ n[3900];
assign t[3901] = t[3900] ^ n[3901];
assign t[3902] = t[3901] ^ n[3902];
assign t[3903] = t[3902] ^ n[3903];
assign t[3904] = t[3903] ^ n[3904];
assign t[3905] = t[3904] ^ n[3905];
assign t[3906] = t[3905] ^ n[3906];
assign t[3907] = t[3906] ^ n[3907];
assign t[3908] = t[3907] ^ n[3908];
assign t[3909] = t[3908] ^ n[3909];
assign t[3910] = t[3909] ^ n[3910];
assign t[3911] = t[3910] ^ n[3911];
assign t[3912] = t[3911] ^ n[3912];
assign t[3913] = t[3912] ^ n[3913];
assign t[3914] = t[3913] ^ n[3914];
assign t[3915] = t[3914] ^ n[3915];
assign t[3916] = t[3915] ^ n[3916];
assign t[3917] = t[3916] ^ n[3917];
assign t[3918] = t[3917] ^ n[3918];
assign t[3919] = t[3918] ^ n[3919];
assign t[3920] = t[3919] ^ n[3920];
assign t[3921] = t[3920] ^ n[3921];
assign t[3922] = t[3921] ^ n[3922];
assign t[3923] = t[3922] ^ n[3923];
assign t[3924] = t[3923] ^ n[3924];
assign t[3925] = t[3924] ^ n[3925];
assign t[3926] = t[3925] ^ n[3926];
assign t[3927] = t[3926] ^ n[3927];
assign t[3928] = t[3927] ^ n[3928];
assign t[3929] = t[3928] ^ n[3929];
assign t[3930] = t[3929] ^ n[3930];
assign t[3931] = t[3930] ^ n[3931];
assign t[3932] = t[3931] ^ n[3932];
assign t[3933] = t[3932] ^ n[3933];
assign t[3934] = t[3933] ^ n[3934];
assign t[3935] = t[3934] ^ n[3935];
assign t[3936] = t[3935] ^ n[3936];
assign t[3937] = t[3936] ^ n[3937];
assign t[3938] = t[3937] ^ n[3938];
assign t[3939] = t[3938] ^ n[3939];
assign t[3940] = t[3939] ^ n[3940];
assign t[3941] = t[3940] ^ n[3941];
assign t[3942] = t[3941] ^ n[3942];
assign t[3943] = t[3942] ^ n[3943];
assign t[3944] = t[3943] ^ n[3944];
assign t[3945] = t[3944] ^ n[3945];
assign t[3946] = t[3945] ^ n[3946];
assign t[3947] = t[3946] ^ n[3947];
assign t[3948] = t[3947] ^ n[3948];
assign t[3949] = t[3948] ^ n[3949];
assign t[3950] = t[3949] ^ n[3950];
assign t[3951] = t[3950] ^ n[3951];
assign t[3952] = t[3951] ^ n[3952];
assign t[3953] = t[3952] ^ n[3953];
assign t[3954] = t[3953] ^ n[3954];
assign t[3955] = t[3954] ^ n[3955];
assign t[3956] = t[3955] ^ n[3956];
assign t[3957] = t[3956] ^ n[3957];
assign t[3958] = t[3957] ^ n[3958];
assign t[3959] = t[3958] ^ n[3959];
assign t[3960] = t[3959] ^ n[3960];
assign t[3961] = t[3960] ^ n[3961];
assign t[3962] = t[3961] ^ n[3962];
assign t[3963] = t[3962] ^ n[3963];
assign t[3964] = t[3963] ^ n[3964];
assign t[3965] = t[3964] ^ n[3965];
assign t[3966] = t[3965] ^ n[3966];
assign t[3967] = t[3966] ^ n[3967];
assign t[3968] = t[3967] ^ n[3968];
assign t[3969] = t[3968] ^ n[3969];
assign t[3970] = t[3969] ^ n[3970];
assign t[3971] = t[3970] ^ n[3971];
assign t[3972] = t[3971] ^ n[3972];
assign t[3973] = t[3972] ^ n[3973];
assign t[3974] = t[3973] ^ n[3974];
assign t[3975] = t[3974] ^ n[3975];
assign t[3976] = t[3975] ^ n[3976];
assign t[3977] = t[3976] ^ n[3977];
assign t[3978] = t[3977] ^ n[3978];
assign t[3979] = t[3978] ^ n[3979];
assign t[3980] = t[3979] ^ n[3980];
assign t[3981] = t[3980] ^ n[3981];
assign t[3982] = t[3981] ^ n[3982];
assign t[3983] = t[3982] ^ n[3983];
assign t[3984] = t[3983] ^ n[3984];
assign t[3985] = t[3984] ^ n[3985];
assign t[3986] = t[3985] ^ n[3986];
assign t[3987] = t[3986] ^ n[3987];
assign t[3988] = t[3987] ^ n[3988];
assign t[3989] = t[3988] ^ n[3989];
assign t[3990] = t[3989] ^ n[3990];
assign t[3991] = t[3990] ^ n[3991];
assign t[3992] = t[3991] ^ n[3992];
assign t[3993] = t[3992] ^ n[3993];
assign t[3994] = t[3993] ^ n[3994];
assign t[3995] = t[3994] ^ n[3995];
assign t[3996] = t[3995] ^ n[3996];
assign t[3997] = t[3996] ^ n[3997];
assign t[3998] = t[3997] ^ n[3998];
assign t[3999] = t[3998] ^ n[3999];
assign t[4000] = t[3999] ^ n[4000];
assign t[4001] = t[4000] ^ n[4001];
assign t[4002] = t[4001] ^ n[4002];
assign t[4003] = t[4002] ^ n[4003];
assign t[4004] = t[4003] ^ n[4004];
assign t[4005] = t[4004] ^ n[4005];
assign t[4006] = t[4005] ^ n[4006];
assign t[4007] = t[4006] ^ n[4007];
assign t[4008] = t[4007] ^ n[4008];
assign t[4009] = t[4008] ^ n[4009];
assign t[4010] = t[4009] ^ n[4010];
assign t[4011] = t[4010] ^ n[4011];
assign t[4012] = t[4011] ^ n[4012];
assign t[4013] = t[4012] ^ n[4013];
assign t[4014] = t[4013] ^ n[4014];
assign t[4015] = t[4014] ^ n[4015];
assign t[4016] = t[4015] ^ n[4016];
assign t[4017] = t[4016] ^ n[4017];
assign t[4018] = t[4017] ^ n[4018];
assign t[4019] = t[4018] ^ n[4019];
assign t[4020] = t[4019] ^ n[4020];
assign t[4021] = t[4020] ^ n[4021];
assign t[4022] = t[4021] ^ n[4022];
assign t[4023] = t[4022] ^ n[4023];
assign t[4024] = t[4023] ^ n[4024];
assign t[4025] = t[4024] ^ n[4025];
assign t[4026] = t[4025] ^ n[4026];
assign t[4027] = t[4026] ^ n[4027];
assign t[4028] = t[4027] ^ n[4028];
assign t[4029] = t[4028] ^ n[4029];
assign t[4030] = t[4029] ^ n[4030];
assign t[4031] = t[4030] ^ n[4031];
assign t[4032] = t[4031] ^ n[4032];
assign t[4033] = t[4032] ^ n[4033];
assign t[4034] = t[4033] ^ n[4034];
assign t[4035] = t[4034] ^ n[4035];
assign t[4036] = t[4035] ^ n[4036];
assign t[4037] = t[4036] ^ n[4037];
assign t[4038] = t[4037] ^ n[4038];
assign t[4039] = t[4038] ^ n[4039];
assign t[4040] = t[4039] ^ n[4040];
assign t[4041] = t[4040] ^ n[4041];
assign t[4042] = t[4041] ^ n[4042];
assign t[4043] = t[4042] ^ n[4043];
assign t[4044] = t[4043] ^ n[4044];
assign t[4045] = t[4044] ^ n[4045];
assign t[4046] = t[4045] ^ n[4046];
assign t[4047] = t[4046] ^ n[4047];
assign t[4048] = t[4047] ^ n[4048];
assign t[4049] = t[4048] ^ n[4049];
assign t[4050] = t[4049] ^ n[4050];
assign t[4051] = t[4050] ^ n[4051];
assign t[4052] = t[4051] ^ n[4052];
assign t[4053] = t[4052] ^ n[4053];
assign t[4054] = t[4053] ^ n[4054];
assign t[4055] = t[4054] ^ n[4055];
assign t[4056] = t[4055] ^ n[4056];
assign t[4057] = t[4056] ^ n[4057];
assign t[4058] = t[4057] ^ n[4058];
assign t[4059] = t[4058] ^ n[4059];
assign t[4060] = t[4059] ^ n[4060];
assign t[4061] = t[4060] ^ n[4061];
assign t[4062] = t[4061] ^ n[4062];
assign t[4063] = t[4062] ^ n[4063];
assign t[4064] = t[4063] ^ n[4064];
assign t[4065] = t[4064] ^ n[4065];
assign t[4066] = t[4065] ^ n[4066];
assign t[4067] = t[4066] ^ n[4067];
assign t[4068] = t[4067] ^ n[4068];
assign t[4069] = t[4068] ^ n[4069];
assign t[4070] = t[4069] ^ n[4070];
assign t[4071] = t[4070] ^ n[4071];
assign t[4072] = t[4071] ^ n[4072];
assign t[4073] = t[4072] ^ n[4073];
assign t[4074] = t[4073] ^ n[4074];
assign t[4075] = t[4074] ^ n[4075];
assign t[4076] = t[4075] ^ n[4076];
assign t[4077] = t[4076] ^ n[4077];
assign t[4078] = t[4077] ^ n[4078];
assign t[4079] = t[4078] ^ n[4079];
assign t[4080] = t[4079] ^ n[4080];
assign t[4081] = t[4080] ^ n[4081];

assign s[10] = ( a[10] ^ b [10] ) ^ t[4081];

//asigning bit 11
assign t[4082] = n[4082];
assign t[4083] = t[4082] ^ n[4083];
assign t[4084] = t[4083] ^ n[4084];
assign t[4085] = t[4084] ^ n[4085];
assign t[4086] = t[4085] ^ n[4086];
assign t[4087] = t[4086] ^ n[4087];
assign t[4088] = t[4087] ^ n[4088];
assign t[4089] = t[4088] ^ n[4089];
assign t[4090] = t[4089] ^ n[4090];
assign t[4091] = t[4090] ^ n[4091];
assign t[4092] = t[4091] ^ n[4092];
assign t[4093] = t[4092] ^ n[4093];
assign t[4094] = t[4093] ^ n[4094];
assign t[4095] = t[4094] ^ n[4095];
assign t[4096] = t[4095] ^ n[4096];
assign t[4097] = t[4096] ^ n[4097];
assign t[4098] = t[4097] ^ n[4098];
assign t[4099] = t[4098] ^ n[4099];
assign t[4100] = t[4099] ^ n[4100];
assign t[4101] = t[4100] ^ n[4101];
assign t[4102] = t[4101] ^ n[4102];
assign t[4103] = t[4102] ^ n[4103];
assign t[4104] = t[4103] ^ n[4104];
assign t[4105] = t[4104] ^ n[4105];
assign t[4106] = t[4105] ^ n[4106];
assign t[4107] = t[4106] ^ n[4107];
assign t[4108] = t[4107] ^ n[4108];
assign t[4109] = t[4108] ^ n[4109];
assign t[4110] = t[4109] ^ n[4110];
assign t[4111] = t[4110] ^ n[4111];
assign t[4112] = t[4111] ^ n[4112];
assign t[4113] = t[4112] ^ n[4113];
assign t[4114] = t[4113] ^ n[4114];
assign t[4115] = t[4114] ^ n[4115];
assign t[4116] = t[4115] ^ n[4116];
assign t[4117] = t[4116] ^ n[4117];
assign t[4118] = t[4117] ^ n[4118];
assign t[4119] = t[4118] ^ n[4119];
assign t[4120] = t[4119] ^ n[4120];
assign t[4121] = t[4120] ^ n[4121];
assign t[4122] = t[4121] ^ n[4122];
assign t[4123] = t[4122] ^ n[4123];
assign t[4124] = t[4123] ^ n[4124];
assign t[4125] = t[4124] ^ n[4125];
assign t[4126] = t[4125] ^ n[4126];
assign t[4127] = t[4126] ^ n[4127];
assign t[4128] = t[4127] ^ n[4128];
assign t[4129] = t[4128] ^ n[4129];
assign t[4130] = t[4129] ^ n[4130];
assign t[4131] = t[4130] ^ n[4131];
assign t[4132] = t[4131] ^ n[4132];
assign t[4133] = t[4132] ^ n[4133];
assign t[4134] = t[4133] ^ n[4134];
assign t[4135] = t[4134] ^ n[4135];
assign t[4136] = t[4135] ^ n[4136];
assign t[4137] = t[4136] ^ n[4137];
assign t[4138] = t[4137] ^ n[4138];
assign t[4139] = t[4138] ^ n[4139];
assign t[4140] = t[4139] ^ n[4140];
assign t[4141] = t[4140] ^ n[4141];
assign t[4142] = t[4141] ^ n[4142];
assign t[4143] = t[4142] ^ n[4143];
assign t[4144] = t[4143] ^ n[4144];
assign t[4145] = t[4144] ^ n[4145];
assign t[4146] = t[4145] ^ n[4146];
assign t[4147] = t[4146] ^ n[4147];
assign t[4148] = t[4147] ^ n[4148];
assign t[4149] = t[4148] ^ n[4149];
assign t[4150] = t[4149] ^ n[4150];
assign t[4151] = t[4150] ^ n[4151];
assign t[4152] = t[4151] ^ n[4152];
assign t[4153] = t[4152] ^ n[4153];
assign t[4154] = t[4153] ^ n[4154];
assign t[4155] = t[4154] ^ n[4155];
assign t[4156] = t[4155] ^ n[4156];
assign t[4157] = t[4156] ^ n[4157];
assign t[4158] = t[4157] ^ n[4158];
assign t[4159] = t[4158] ^ n[4159];
assign t[4160] = t[4159] ^ n[4160];
assign t[4161] = t[4160] ^ n[4161];
assign t[4162] = t[4161] ^ n[4162];
assign t[4163] = t[4162] ^ n[4163];
assign t[4164] = t[4163] ^ n[4164];
assign t[4165] = t[4164] ^ n[4165];
assign t[4166] = t[4165] ^ n[4166];
assign t[4167] = t[4166] ^ n[4167];
assign t[4168] = t[4167] ^ n[4168];
assign t[4169] = t[4168] ^ n[4169];
assign t[4170] = t[4169] ^ n[4170];
assign t[4171] = t[4170] ^ n[4171];
assign t[4172] = t[4171] ^ n[4172];
assign t[4173] = t[4172] ^ n[4173];
assign t[4174] = t[4173] ^ n[4174];
assign t[4175] = t[4174] ^ n[4175];
assign t[4176] = t[4175] ^ n[4176];
assign t[4177] = t[4176] ^ n[4177];
assign t[4178] = t[4177] ^ n[4178];
assign t[4179] = t[4178] ^ n[4179];
assign t[4180] = t[4179] ^ n[4180];
assign t[4181] = t[4180] ^ n[4181];
assign t[4182] = t[4181] ^ n[4182];
assign t[4183] = t[4182] ^ n[4183];
assign t[4184] = t[4183] ^ n[4184];
assign t[4185] = t[4184] ^ n[4185];
assign t[4186] = t[4185] ^ n[4186];
assign t[4187] = t[4186] ^ n[4187];
assign t[4188] = t[4187] ^ n[4188];
assign t[4189] = t[4188] ^ n[4189];
assign t[4190] = t[4189] ^ n[4190];
assign t[4191] = t[4190] ^ n[4191];
assign t[4192] = t[4191] ^ n[4192];
assign t[4193] = t[4192] ^ n[4193];
assign t[4194] = t[4193] ^ n[4194];
assign t[4195] = t[4194] ^ n[4195];
assign t[4196] = t[4195] ^ n[4196];
assign t[4197] = t[4196] ^ n[4197];
assign t[4198] = t[4197] ^ n[4198];
assign t[4199] = t[4198] ^ n[4199];
assign t[4200] = t[4199] ^ n[4200];
assign t[4201] = t[4200] ^ n[4201];
assign t[4202] = t[4201] ^ n[4202];
assign t[4203] = t[4202] ^ n[4203];
assign t[4204] = t[4203] ^ n[4204];
assign t[4205] = t[4204] ^ n[4205];
assign t[4206] = t[4205] ^ n[4206];
assign t[4207] = t[4206] ^ n[4207];
assign t[4208] = t[4207] ^ n[4208];
assign t[4209] = t[4208] ^ n[4209];
assign t[4210] = t[4209] ^ n[4210];
assign t[4211] = t[4210] ^ n[4211];
assign t[4212] = t[4211] ^ n[4212];
assign t[4213] = t[4212] ^ n[4213];
assign t[4214] = t[4213] ^ n[4214];
assign t[4215] = t[4214] ^ n[4215];
assign t[4216] = t[4215] ^ n[4216];
assign t[4217] = t[4216] ^ n[4217];
assign t[4218] = t[4217] ^ n[4218];
assign t[4219] = t[4218] ^ n[4219];
assign t[4220] = t[4219] ^ n[4220];
assign t[4221] = t[4220] ^ n[4221];
assign t[4222] = t[4221] ^ n[4222];
assign t[4223] = t[4222] ^ n[4223];
assign t[4224] = t[4223] ^ n[4224];
assign t[4225] = t[4224] ^ n[4225];
assign t[4226] = t[4225] ^ n[4226];
assign t[4227] = t[4226] ^ n[4227];
assign t[4228] = t[4227] ^ n[4228];
assign t[4229] = t[4228] ^ n[4229];
assign t[4230] = t[4229] ^ n[4230];
assign t[4231] = t[4230] ^ n[4231];
assign t[4232] = t[4231] ^ n[4232];
assign t[4233] = t[4232] ^ n[4233];
assign t[4234] = t[4233] ^ n[4234];
assign t[4235] = t[4234] ^ n[4235];
assign t[4236] = t[4235] ^ n[4236];
assign t[4237] = t[4236] ^ n[4237];
assign t[4238] = t[4237] ^ n[4238];
assign t[4239] = t[4238] ^ n[4239];
assign t[4240] = t[4239] ^ n[4240];
assign t[4241] = t[4240] ^ n[4241];
assign t[4242] = t[4241] ^ n[4242];
assign t[4243] = t[4242] ^ n[4243];
assign t[4244] = t[4243] ^ n[4244];
assign t[4245] = t[4244] ^ n[4245];
assign t[4246] = t[4245] ^ n[4246];
assign t[4247] = t[4246] ^ n[4247];
assign t[4248] = t[4247] ^ n[4248];
assign t[4249] = t[4248] ^ n[4249];
assign t[4250] = t[4249] ^ n[4250];
assign t[4251] = t[4250] ^ n[4251];
assign t[4252] = t[4251] ^ n[4252];
assign t[4253] = t[4252] ^ n[4253];
assign t[4254] = t[4253] ^ n[4254];
assign t[4255] = t[4254] ^ n[4255];
assign t[4256] = t[4255] ^ n[4256];
assign t[4257] = t[4256] ^ n[4257];
assign t[4258] = t[4257] ^ n[4258];
assign t[4259] = t[4258] ^ n[4259];
assign t[4260] = t[4259] ^ n[4260];
assign t[4261] = t[4260] ^ n[4261];
assign t[4262] = t[4261] ^ n[4262];
assign t[4263] = t[4262] ^ n[4263];
assign t[4264] = t[4263] ^ n[4264];
assign t[4265] = t[4264] ^ n[4265];
assign t[4266] = t[4265] ^ n[4266];
assign t[4267] = t[4266] ^ n[4267];
assign t[4268] = t[4267] ^ n[4268];
assign t[4269] = t[4268] ^ n[4269];
assign t[4270] = t[4269] ^ n[4270];
assign t[4271] = t[4270] ^ n[4271];
assign t[4272] = t[4271] ^ n[4272];
assign t[4273] = t[4272] ^ n[4273];
assign t[4274] = t[4273] ^ n[4274];
assign t[4275] = t[4274] ^ n[4275];
assign t[4276] = t[4275] ^ n[4276];
assign t[4277] = t[4276] ^ n[4277];
assign t[4278] = t[4277] ^ n[4278];
assign t[4279] = t[4278] ^ n[4279];
assign t[4280] = t[4279] ^ n[4280];
assign t[4281] = t[4280] ^ n[4281];
assign t[4282] = t[4281] ^ n[4282];
assign t[4283] = t[4282] ^ n[4283];
assign t[4284] = t[4283] ^ n[4284];
assign t[4285] = t[4284] ^ n[4285];
assign t[4286] = t[4285] ^ n[4286];
assign t[4287] = t[4286] ^ n[4287];
assign t[4288] = t[4287] ^ n[4288];
assign t[4289] = t[4288] ^ n[4289];
assign t[4290] = t[4289] ^ n[4290];
assign t[4291] = t[4290] ^ n[4291];
assign t[4292] = t[4291] ^ n[4292];
assign t[4293] = t[4292] ^ n[4293];
assign t[4294] = t[4293] ^ n[4294];
assign t[4295] = t[4294] ^ n[4295];
assign t[4296] = t[4295] ^ n[4296];
assign t[4297] = t[4296] ^ n[4297];
assign t[4298] = t[4297] ^ n[4298];
assign t[4299] = t[4298] ^ n[4299];
assign t[4300] = t[4299] ^ n[4300];
assign t[4301] = t[4300] ^ n[4301];
assign t[4302] = t[4301] ^ n[4302];
assign t[4303] = t[4302] ^ n[4303];
assign t[4304] = t[4303] ^ n[4304];
assign t[4305] = t[4304] ^ n[4305];
assign t[4306] = t[4305] ^ n[4306];
assign t[4307] = t[4306] ^ n[4307];
assign t[4308] = t[4307] ^ n[4308];
assign t[4309] = t[4308] ^ n[4309];
assign t[4310] = t[4309] ^ n[4310];
assign t[4311] = t[4310] ^ n[4311];
assign t[4312] = t[4311] ^ n[4312];
assign t[4313] = t[4312] ^ n[4313];
assign t[4314] = t[4313] ^ n[4314];
assign t[4315] = t[4314] ^ n[4315];
assign t[4316] = t[4315] ^ n[4316];
assign t[4317] = t[4316] ^ n[4317];
assign t[4318] = t[4317] ^ n[4318];
assign t[4319] = t[4318] ^ n[4319];
assign t[4320] = t[4319] ^ n[4320];
assign t[4321] = t[4320] ^ n[4321];
assign t[4322] = t[4321] ^ n[4322];
assign t[4323] = t[4322] ^ n[4323];
assign t[4324] = t[4323] ^ n[4324];
assign t[4325] = t[4324] ^ n[4325];
assign t[4326] = t[4325] ^ n[4326];
assign t[4327] = t[4326] ^ n[4327];
assign t[4328] = t[4327] ^ n[4328];
assign t[4329] = t[4328] ^ n[4329];
assign t[4330] = t[4329] ^ n[4330];
assign t[4331] = t[4330] ^ n[4331];
assign t[4332] = t[4331] ^ n[4332];
assign t[4333] = t[4332] ^ n[4333];
assign t[4334] = t[4333] ^ n[4334];
assign t[4335] = t[4334] ^ n[4335];
assign t[4336] = t[4335] ^ n[4336];
assign t[4337] = t[4336] ^ n[4337];
assign t[4338] = t[4337] ^ n[4338];
assign t[4339] = t[4338] ^ n[4339];
assign t[4340] = t[4339] ^ n[4340];
assign t[4341] = t[4340] ^ n[4341];
assign t[4342] = t[4341] ^ n[4342];
assign t[4343] = t[4342] ^ n[4343];
assign t[4344] = t[4343] ^ n[4344];
assign t[4345] = t[4344] ^ n[4345];
assign t[4346] = t[4345] ^ n[4346];
assign t[4347] = t[4346] ^ n[4347];
assign t[4348] = t[4347] ^ n[4348];
assign t[4349] = t[4348] ^ n[4349];
assign t[4350] = t[4349] ^ n[4350];
assign t[4351] = t[4350] ^ n[4351];
assign t[4352] = t[4351] ^ n[4352];
assign t[4353] = t[4352] ^ n[4353];
assign t[4354] = t[4353] ^ n[4354];
assign t[4355] = t[4354] ^ n[4355];
assign t[4356] = t[4355] ^ n[4356];
assign t[4357] = t[4356] ^ n[4357];
assign t[4358] = t[4357] ^ n[4358];
assign t[4359] = t[4358] ^ n[4359];
assign t[4360] = t[4359] ^ n[4360];
assign t[4361] = t[4360] ^ n[4361];
assign t[4362] = t[4361] ^ n[4362];
assign t[4363] = t[4362] ^ n[4363];
assign t[4364] = t[4363] ^ n[4364];
assign t[4365] = t[4364] ^ n[4365];
assign t[4366] = t[4365] ^ n[4366];
assign t[4367] = t[4366] ^ n[4367];
assign t[4368] = t[4367] ^ n[4368];
assign t[4369] = t[4368] ^ n[4369];
assign t[4370] = t[4369] ^ n[4370];
assign t[4371] = t[4370] ^ n[4371];
assign t[4372] = t[4371] ^ n[4372];
assign t[4373] = t[4372] ^ n[4373];
assign t[4374] = t[4373] ^ n[4374];
assign t[4375] = t[4374] ^ n[4375];
assign t[4376] = t[4375] ^ n[4376];
assign t[4377] = t[4376] ^ n[4377];
assign t[4378] = t[4377] ^ n[4378];
assign t[4379] = t[4378] ^ n[4379];
assign t[4380] = t[4379] ^ n[4380];
assign t[4381] = t[4380] ^ n[4381];
assign t[4382] = t[4381] ^ n[4382];
assign t[4383] = t[4382] ^ n[4383];
assign t[4384] = t[4383] ^ n[4384];
assign t[4385] = t[4384] ^ n[4385];
assign t[4386] = t[4385] ^ n[4386];
assign t[4387] = t[4386] ^ n[4387];
assign t[4388] = t[4387] ^ n[4388];
assign t[4389] = t[4388] ^ n[4389];
assign t[4390] = t[4389] ^ n[4390];
assign t[4391] = t[4390] ^ n[4391];
assign t[4392] = t[4391] ^ n[4392];
assign t[4393] = t[4392] ^ n[4393];
assign t[4394] = t[4393] ^ n[4394];
assign t[4395] = t[4394] ^ n[4395];
assign t[4396] = t[4395] ^ n[4396];
assign t[4397] = t[4396] ^ n[4397];
assign t[4398] = t[4397] ^ n[4398];
assign t[4399] = t[4398] ^ n[4399];
assign t[4400] = t[4399] ^ n[4400];
assign t[4401] = t[4400] ^ n[4401];
assign t[4402] = t[4401] ^ n[4402];
assign t[4403] = t[4402] ^ n[4403];
assign t[4404] = t[4403] ^ n[4404];
assign t[4405] = t[4404] ^ n[4405];
assign t[4406] = t[4405] ^ n[4406];
assign t[4407] = t[4406] ^ n[4407];
assign t[4408] = t[4407] ^ n[4408];
assign t[4409] = t[4408] ^ n[4409];
assign t[4410] = t[4409] ^ n[4410];
assign t[4411] = t[4410] ^ n[4411];
assign t[4412] = t[4411] ^ n[4412];
assign t[4413] = t[4412] ^ n[4413];
assign t[4414] = t[4413] ^ n[4414];
assign t[4415] = t[4414] ^ n[4415];
assign t[4416] = t[4415] ^ n[4416];
assign t[4417] = t[4416] ^ n[4417];
assign t[4418] = t[4417] ^ n[4418];
assign t[4419] = t[4418] ^ n[4419];
assign t[4420] = t[4419] ^ n[4420];
assign t[4421] = t[4420] ^ n[4421];
assign t[4422] = t[4421] ^ n[4422];
assign t[4423] = t[4422] ^ n[4423];
assign t[4424] = t[4423] ^ n[4424];
assign t[4425] = t[4424] ^ n[4425];
assign t[4426] = t[4425] ^ n[4426];
assign t[4427] = t[4426] ^ n[4427];
assign t[4428] = t[4427] ^ n[4428];
assign t[4429] = t[4428] ^ n[4429];
assign t[4430] = t[4429] ^ n[4430];
assign t[4431] = t[4430] ^ n[4431];
assign t[4432] = t[4431] ^ n[4432];
assign t[4433] = t[4432] ^ n[4433];
assign t[4434] = t[4433] ^ n[4434];
assign t[4435] = t[4434] ^ n[4435];
assign t[4436] = t[4435] ^ n[4436];
assign t[4437] = t[4436] ^ n[4437];
assign t[4438] = t[4437] ^ n[4438];
assign t[4439] = t[4438] ^ n[4439];
assign t[4440] = t[4439] ^ n[4440];
assign t[4441] = t[4440] ^ n[4441];
assign t[4442] = t[4441] ^ n[4442];
assign t[4443] = t[4442] ^ n[4443];
assign t[4444] = t[4443] ^ n[4444];
assign t[4445] = t[4444] ^ n[4445];
assign t[4446] = t[4445] ^ n[4446];
assign t[4447] = t[4446] ^ n[4447];
assign t[4448] = t[4447] ^ n[4448];
assign t[4449] = t[4448] ^ n[4449];
assign t[4450] = t[4449] ^ n[4450];
assign t[4451] = t[4450] ^ n[4451];
assign t[4452] = t[4451] ^ n[4452];
assign t[4453] = t[4452] ^ n[4453];
assign t[4454] = t[4453] ^ n[4454];
assign t[4455] = t[4454] ^ n[4455];
assign t[4456] = t[4455] ^ n[4456];
assign t[4457] = t[4456] ^ n[4457];
assign t[4458] = t[4457] ^ n[4458];
assign t[4459] = t[4458] ^ n[4459];
assign t[4460] = t[4459] ^ n[4460];
assign t[4461] = t[4460] ^ n[4461];
assign t[4462] = t[4461] ^ n[4462];
assign t[4463] = t[4462] ^ n[4463];
assign t[4464] = t[4463] ^ n[4464];
assign t[4465] = t[4464] ^ n[4465];
assign t[4466] = t[4465] ^ n[4466];
assign t[4467] = t[4466] ^ n[4467];
assign t[4468] = t[4467] ^ n[4468];
assign t[4469] = t[4468] ^ n[4469];
assign t[4470] = t[4469] ^ n[4470];
assign t[4471] = t[4470] ^ n[4471];
assign t[4472] = t[4471] ^ n[4472];
assign t[4473] = t[4472] ^ n[4473];
assign t[4474] = t[4473] ^ n[4474];
assign t[4475] = t[4474] ^ n[4475];
assign t[4476] = t[4475] ^ n[4476];
assign t[4477] = t[4476] ^ n[4477];
assign t[4478] = t[4477] ^ n[4478];
assign t[4479] = t[4478] ^ n[4479];
assign t[4480] = t[4479] ^ n[4480];
assign t[4481] = t[4480] ^ n[4481];
assign t[4482] = t[4481] ^ n[4482];
assign t[4483] = t[4482] ^ n[4483];
assign t[4484] = t[4483] ^ n[4484];
assign t[4485] = t[4484] ^ n[4485];
assign t[4486] = t[4485] ^ n[4486];
assign t[4487] = t[4486] ^ n[4487];
assign t[4488] = t[4487] ^ n[4488];
assign t[4489] = t[4488] ^ n[4489];
assign t[4490] = t[4489] ^ n[4490];
assign t[4491] = t[4490] ^ n[4491];
assign t[4492] = t[4491] ^ n[4492];
assign t[4493] = t[4492] ^ n[4493];
assign t[4494] = t[4493] ^ n[4494];
assign t[4495] = t[4494] ^ n[4495];
assign t[4496] = t[4495] ^ n[4496];
assign t[4497] = t[4496] ^ n[4497];
assign t[4498] = t[4497] ^ n[4498];
assign t[4499] = t[4498] ^ n[4499];
assign t[4500] = t[4499] ^ n[4500];
assign t[4501] = t[4500] ^ n[4501];
assign t[4502] = t[4501] ^ n[4502];
assign t[4503] = t[4502] ^ n[4503];
assign t[4504] = t[4503] ^ n[4504];
assign t[4505] = t[4504] ^ n[4505];
assign t[4506] = t[4505] ^ n[4506];
assign t[4507] = t[4506] ^ n[4507];
assign t[4508] = t[4507] ^ n[4508];
assign t[4509] = t[4508] ^ n[4509];
assign t[4510] = t[4509] ^ n[4510];
assign t[4511] = t[4510] ^ n[4511];
assign t[4512] = t[4511] ^ n[4512];
assign t[4513] = t[4512] ^ n[4513];
assign t[4514] = t[4513] ^ n[4514];
assign t[4515] = t[4514] ^ n[4515];
assign t[4516] = t[4515] ^ n[4516];
assign t[4517] = t[4516] ^ n[4517];
assign t[4518] = t[4517] ^ n[4518];
assign t[4519] = t[4518] ^ n[4519];
assign t[4520] = t[4519] ^ n[4520];
assign t[4521] = t[4520] ^ n[4521];
assign t[4522] = t[4521] ^ n[4522];
assign t[4523] = t[4522] ^ n[4523];
assign t[4524] = t[4523] ^ n[4524];
assign t[4525] = t[4524] ^ n[4525];
assign t[4526] = t[4525] ^ n[4526];
assign t[4527] = t[4526] ^ n[4527];
assign t[4528] = t[4527] ^ n[4528];
assign t[4529] = t[4528] ^ n[4529];
assign t[4530] = t[4529] ^ n[4530];
assign t[4531] = t[4530] ^ n[4531];
assign t[4532] = t[4531] ^ n[4532];
assign t[4533] = t[4532] ^ n[4533];
assign t[4534] = t[4533] ^ n[4534];
assign t[4535] = t[4534] ^ n[4535];
assign t[4536] = t[4535] ^ n[4536];
assign t[4537] = t[4536] ^ n[4537];
assign t[4538] = t[4537] ^ n[4538];
assign t[4539] = t[4538] ^ n[4539];
assign t[4540] = t[4539] ^ n[4540];
assign t[4541] = t[4540] ^ n[4541];
assign t[4542] = t[4541] ^ n[4542];
assign t[4543] = t[4542] ^ n[4543];
assign t[4544] = t[4543] ^ n[4544];
assign t[4545] = t[4544] ^ n[4545];
assign t[4546] = t[4545] ^ n[4546];
assign t[4547] = t[4546] ^ n[4547];
assign t[4548] = t[4547] ^ n[4548];
assign t[4549] = t[4548] ^ n[4549];
assign t[4550] = t[4549] ^ n[4550];
assign t[4551] = t[4550] ^ n[4551];
assign t[4552] = t[4551] ^ n[4552];
assign t[4553] = t[4552] ^ n[4553];
assign t[4554] = t[4553] ^ n[4554];
assign t[4555] = t[4554] ^ n[4555];
assign t[4556] = t[4555] ^ n[4556];
assign t[4557] = t[4556] ^ n[4557];
assign t[4558] = t[4557] ^ n[4558];
assign t[4559] = t[4558] ^ n[4559];
assign t[4560] = t[4559] ^ n[4560];
assign t[4561] = t[4560] ^ n[4561];
assign t[4562] = t[4561] ^ n[4562];
assign t[4563] = t[4562] ^ n[4563];
assign t[4564] = t[4563] ^ n[4564];
assign t[4565] = t[4564] ^ n[4565];
assign t[4566] = t[4565] ^ n[4566];
assign t[4567] = t[4566] ^ n[4567];
assign t[4568] = t[4567] ^ n[4568];
assign t[4569] = t[4568] ^ n[4569];
assign t[4570] = t[4569] ^ n[4570];
assign t[4571] = t[4570] ^ n[4571];
assign t[4572] = t[4571] ^ n[4572];
assign t[4573] = t[4572] ^ n[4573];
assign t[4574] = t[4573] ^ n[4574];
assign t[4575] = t[4574] ^ n[4575];
assign t[4576] = t[4575] ^ n[4576];
assign t[4577] = t[4576] ^ n[4577];
assign t[4578] = t[4577] ^ n[4578];
assign t[4579] = t[4578] ^ n[4579];
assign t[4580] = t[4579] ^ n[4580];
assign t[4581] = t[4580] ^ n[4581];
assign t[4582] = t[4581] ^ n[4582];
assign t[4583] = t[4582] ^ n[4583];
assign t[4584] = t[4583] ^ n[4584];
assign t[4585] = t[4584] ^ n[4585];
assign t[4586] = t[4585] ^ n[4586];
assign t[4587] = t[4586] ^ n[4587];
assign t[4588] = t[4587] ^ n[4588];
assign t[4589] = t[4588] ^ n[4589];
assign t[4590] = t[4589] ^ n[4590];
assign t[4591] = t[4590] ^ n[4591];
assign t[4592] = t[4591] ^ n[4592];
assign t[4593] = t[4592] ^ n[4593];
assign t[4594] = t[4593] ^ n[4594];
assign t[4595] = t[4594] ^ n[4595];
assign t[4596] = t[4595] ^ n[4596];
assign t[4597] = t[4596] ^ n[4597];
assign t[4598] = t[4597] ^ n[4598];
assign t[4599] = t[4598] ^ n[4599];
assign t[4600] = t[4599] ^ n[4600];
assign t[4601] = t[4600] ^ n[4601];
assign t[4602] = t[4601] ^ n[4602];
assign t[4603] = t[4602] ^ n[4603];
assign t[4604] = t[4603] ^ n[4604];
assign t[4605] = t[4604] ^ n[4605];
assign t[4606] = t[4605] ^ n[4606];
assign t[4607] = t[4606] ^ n[4607];
assign t[4608] = t[4607] ^ n[4608];
assign t[4609] = t[4608] ^ n[4609];
assign t[4610] = t[4609] ^ n[4610];
assign t[4611] = t[4610] ^ n[4611];
assign t[4612] = t[4611] ^ n[4612];
assign t[4613] = t[4612] ^ n[4613];
assign t[4614] = t[4613] ^ n[4614];
assign t[4615] = t[4614] ^ n[4615];
assign t[4616] = t[4615] ^ n[4616];
assign t[4617] = t[4616] ^ n[4617];
assign t[4618] = t[4617] ^ n[4618];
assign t[4619] = t[4618] ^ n[4619];
assign t[4620] = t[4619] ^ n[4620];
assign t[4621] = t[4620] ^ n[4621];
assign t[4622] = t[4621] ^ n[4622];
assign t[4623] = t[4622] ^ n[4623];
assign t[4624] = t[4623] ^ n[4624];
assign t[4625] = t[4624] ^ n[4625];
assign t[4626] = t[4625] ^ n[4626];
assign t[4627] = t[4626] ^ n[4627];
assign t[4628] = t[4627] ^ n[4628];
assign t[4629] = t[4628] ^ n[4629];
assign t[4630] = t[4629] ^ n[4630];
assign t[4631] = t[4630] ^ n[4631];
assign t[4632] = t[4631] ^ n[4632];
assign t[4633] = t[4632] ^ n[4633];
assign t[4634] = t[4633] ^ n[4634];
assign t[4635] = t[4634] ^ n[4635];
assign t[4636] = t[4635] ^ n[4636];
assign t[4637] = t[4636] ^ n[4637];
assign t[4638] = t[4637] ^ n[4638];
assign t[4639] = t[4638] ^ n[4639];
assign t[4640] = t[4639] ^ n[4640];
assign t[4641] = t[4640] ^ n[4641];
assign t[4642] = t[4641] ^ n[4642];
assign t[4643] = t[4642] ^ n[4643];
assign t[4644] = t[4643] ^ n[4644];
assign t[4645] = t[4644] ^ n[4645];
assign t[4646] = t[4645] ^ n[4646];
assign t[4647] = t[4646] ^ n[4647];
assign t[4648] = t[4647] ^ n[4648];
assign t[4649] = t[4648] ^ n[4649];
assign t[4650] = t[4649] ^ n[4650];
assign t[4651] = t[4650] ^ n[4651];
assign t[4652] = t[4651] ^ n[4652];
assign t[4653] = t[4652] ^ n[4653];
assign t[4654] = t[4653] ^ n[4654];
assign t[4655] = t[4654] ^ n[4655];
assign t[4656] = t[4655] ^ n[4656];
assign t[4657] = t[4656] ^ n[4657];
assign t[4658] = t[4657] ^ n[4658];
assign t[4659] = t[4658] ^ n[4659];
assign t[4660] = t[4659] ^ n[4660];
assign t[4661] = t[4660] ^ n[4661];
assign t[4662] = t[4661] ^ n[4662];
assign t[4663] = t[4662] ^ n[4663];
assign t[4664] = t[4663] ^ n[4664];
assign t[4665] = t[4664] ^ n[4665];
assign t[4666] = t[4665] ^ n[4666];
assign t[4667] = t[4666] ^ n[4667];
assign t[4668] = t[4667] ^ n[4668];
assign t[4669] = t[4668] ^ n[4669];
assign t[4670] = t[4669] ^ n[4670];
assign t[4671] = t[4670] ^ n[4671];
assign t[4672] = t[4671] ^ n[4672];
assign t[4673] = t[4672] ^ n[4673];
assign t[4674] = t[4673] ^ n[4674];
assign t[4675] = t[4674] ^ n[4675];
assign t[4676] = t[4675] ^ n[4676];
assign t[4677] = t[4676] ^ n[4677];
assign t[4678] = t[4677] ^ n[4678];
assign t[4679] = t[4678] ^ n[4679];
assign t[4680] = t[4679] ^ n[4680];
assign t[4681] = t[4680] ^ n[4681];
assign t[4682] = t[4681] ^ n[4682];
assign t[4683] = t[4682] ^ n[4683];
assign t[4684] = t[4683] ^ n[4684];
assign t[4685] = t[4684] ^ n[4685];
assign t[4686] = t[4685] ^ n[4686];
assign t[4687] = t[4686] ^ n[4687];
assign t[4688] = t[4687] ^ n[4688];
assign t[4689] = t[4688] ^ n[4689];
assign t[4690] = t[4689] ^ n[4690];
assign t[4691] = t[4690] ^ n[4691];
assign t[4692] = t[4691] ^ n[4692];
assign t[4693] = t[4692] ^ n[4693];
assign t[4694] = t[4693] ^ n[4694];
assign t[4695] = t[4694] ^ n[4695];
assign t[4696] = t[4695] ^ n[4696];
assign t[4697] = t[4696] ^ n[4697];
assign t[4698] = t[4697] ^ n[4698];
assign t[4699] = t[4698] ^ n[4699];
assign t[4700] = t[4699] ^ n[4700];
assign t[4701] = t[4700] ^ n[4701];
assign t[4702] = t[4701] ^ n[4702];
assign t[4703] = t[4702] ^ n[4703];
assign t[4704] = t[4703] ^ n[4704];
assign t[4705] = t[4704] ^ n[4705];
assign t[4706] = t[4705] ^ n[4706];
assign t[4707] = t[4706] ^ n[4707];
assign t[4708] = t[4707] ^ n[4708];
assign t[4709] = t[4708] ^ n[4709];
assign t[4710] = t[4709] ^ n[4710];
assign t[4711] = t[4710] ^ n[4711];
assign t[4712] = t[4711] ^ n[4712];
assign t[4713] = t[4712] ^ n[4713];
assign t[4714] = t[4713] ^ n[4714];
assign t[4715] = t[4714] ^ n[4715];
assign t[4716] = t[4715] ^ n[4716];
assign t[4717] = t[4716] ^ n[4717];
assign t[4718] = t[4717] ^ n[4718];
assign t[4719] = t[4718] ^ n[4719];
assign t[4720] = t[4719] ^ n[4720];
assign t[4721] = t[4720] ^ n[4721];
assign t[4722] = t[4721] ^ n[4722];
assign t[4723] = t[4722] ^ n[4723];
assign t[4724] = t[4723] ^ n[4724];
assign t[4725] = t[4724] ^ n[4725];
assign t[4726] = t[4725] ^ n[4726];
assign t[4727] = t[4726] ^ n[4727];
assign t[4728] = t[4727] ^ n[4728];
assign t[4729] = t[4728] ^ n[4729];
assign t[4730] = t[4729] ^ n[4730];
assign t[4731] = t[4730] ^ n[4731];
assign t[4732] = t[4731] ^ n[4732];
assign t[4733] = t[4732] ^ n[4733];
assign t[4734] = t[4733] ^ n[4734];
assign t[4735] = t[4734] ^ n[4735];
assign t[4736] = t[4735] ^ n[4736];
assign t[4737] = t[4736] ^ n[4737];
assign t[4738] = t[4737] ^ n[4738];
assign t[4739] = t[4738] ^ n[4739];
assign t[4740] = t[4739] ^ n[4740];
assign t[4741] = t[4740] ^ n[4741];
assign t[4742] = t[4741] ^ n[4742];
assign t[4743] = t[4742] ^ n[4743];
assign t[4744] = t[4743] ^ n[4744];
assign t[4745] = t[4744] ^ n[4745];
assign t[4746] = t[4745] ^ n[4746];
assign t[4747] = t[4746] ^ n[4747];
assign t[4748] = t[4747] ^ n[4748];
assign t[4749] = t[4748] ^ n[4749];
assign t[4750] = t[4749] ^ n[4750];
assign t[4751] = t[4750] ^ n[4751];
assign t[4752] = t[4751] ^ n[4752];
assign t[4753] = t[4752] ^ n[4753];
assign t[4754] = t[4753] ^ n[4754];
assign t[4755] = t[4754] ^ n[4755];
assign t[4756] = t[4755] ^ n[4756];
assign t[4757] = t[4756] ^ n[4757];
assign t[4758] = t[4757] ^ n[4758];
assign t[4759] = t[4758] ^ n[4759];
assign t[4760] = t[4759] ^ n[4760];
assign t[4761] = t[4760] ^ n[4761];
assign t[4762] = t[4761] ^ n[4762];
assign t[4763] = t[4762] ^ n[4763];
assign t[4764] = t[4763] ^ n[4764];
assign t[4765] = t[4764] ^ n[4765];
assign t[4766] = t[4765] ^ n[4766];
assign t[4767] = t[4766] ^ n[4767];
assign t[4768] = t[4767] ^ n[4768];
assign t[4769] = t[4768] ^ n[4769];
assign t[4770] = t[4769] ^ n[4770];
assign t[4771] = t[4770] ^ n[4771];
assign t[4772] = t[4771] ^ n[4772];
assign t[4773] = t[4772] ^ n[4773];
assign t[4774] = t[4773] ^ n[4774];
assign t[4775] = t[4774] ^ n[4775];
assign t[4776] = t[4775] ^ n[4776];
assign t[4777] = t[4776] ^ n[4777];
assign t[4778] = t[4777] ^ n[4778];
assign t[4779] = t[4778] ^ n[4779];
assign t[4780] = t[4779] ^ n[4780];
assign t[4781] = t[4780] ^ n[4781];
assign t[4782] = t[4781] ^ n[4782];
assign t[4783] = t[4782] ^ n[4783];
assign t[4784] = t[4783] ^ n[4784];
assign t[4785] = t[4784] ^ n[4785];
assign t[4786] = t[4785] ^ n[4786];
assign t[4787] = t[4786] ^ n[4787];
assign t[4788] = t[4787] ^ n[4788];
assign t[4789] = t[4788] ^ n[4789];
assign t[4790] = t[4789] ^ n[4790];
assign t[4791] = t[4790] ^ n[4791];
assign t[4792] = t[4791] ^ n[4792];
assign t[4793] = t[4792] ^ n[4793];
assign t[4794] = t[4793] ^ n[4794];
assign t[4795] = t[4794] ^ n[4795];
assign t[4796] = t[4795] ^ n[4796];
assign t[4797] = t[4796] ^ n[4797];
assign t[4798] = t[4797] ^ n[4798];
assign t[4799] = t[4798] ^ n[4799];
assign t[4800] = t[4799] ^ n[4800];
assign t[4801] = t[4800] ^ n[4801];
assign t[4802] = t[4801] ^ n[4802];
assign t[4803] = t[4802] ^ n[4803];
assign t[4804] = t[4803] ^ n[4804];
assign t[4805] = t[4804] ^ n[4805];
assign t[4806] = t[4805] ^ n[4806];
assign t[4807] = t[4806] ^ n[4807];
assign t[4808] = t[4807] ^ n[4808];
assign t[4809] = t[4808] ^ n[4809];
assign t[4810] = t[4809] ^ n[4810];
assign t[4811] = t[4810] ^ n[4811];
assign t[4812] = t[4811] ^ n[4812];
assign t[4813] = t[4812] ^ n[4813];
assign t[4814] = t[4813] ^ n[4814];
assign t[4815] = t[4814] ^ n[4815];
assign t[4816] = t[4815] ^ n[4816];
assign t[4817] = t[4816] ^ n[4817];
assign t[4818] = t[4817] ^ n[4818];
assign t[4819] = t[4818] ^ n[4819];
assign t[4820] = t[4819] ^ n[4820];
assign t[4821] = t[4820] ^ n[4821];
assign t[4822] = t[4821] ^ n[4822];
assign t[4823] = t[4822] ^ n[4823];
assign t[4824] = t[4823] ^ n[4824];
assign t[4825] = t[4824] ^ n[4825];
assign t[4826] = t[4825] ^ n[4826];
assign t[4827] = t[4826] ^ n[4827];
assign t[4828] = t[4827] ^ n[4828];
assign t[4829] = t[4828] ^ n[4829];
assign t[4830] = t[4829] ^ n[4830];
assign t[4831] = t[4830] ^ n[4831];
assign t[4832] = t[4831] ^ n[4832];
assign t[4833] = t[4832] ^ n[4833];
assign t[4834] = t[4833] ^ n[4834];
assign t[4835] = t[4834] ^ n[4835];
assign t[4836] = t[4835] ^ n[4836];
assign t[4837] = t[4836] ^ n[4837];
assign t[4838] = t[4837] ^ n[4838];
assign t[4839] = t[4838] ^ n[4839];
assign t[4840] = t[4839] ^ n[4840];
assign t[4841] = t[4840] ^ n[4841];
assign t[4842] = t[4841] ^ n[4842];
assign t[4843] = t[4842] ^ n[4843];
assign t[4844] = t[4843] ^ n[4844];
assign t[4845] = t[4844] ^ n[4845];
assign t[4846] = t[4845] ^ n[4846];
assign t[4847] = t[4846] ^ n[4847];
assign t[4848] = t[4847] ^ n[4848];
assign t[4849] = t[4848] ^ n[4849];
assign t[4850] = t[4849] ^ n[4850];
assign t[4851] = t[4850] ^ n[4851];
assign t[4852] = t[4851] ^ n[4852];
assign t[4853] = t[4852] ^ n[4853];
assign t[4854] = t[4853] ^ n[4854];
assign t[4855] = t[4854] ^ n[4855];
assign t[4856] = t[4855] ^ n[4856];
assign t[4857] = t[4856] ^ n[4857];
assign t[4858] = t[4857] ^ n[4858];
assign t[4859] = t[4858] ^ n[4859];
assign t[4860] = t[4859] ^ n[4860];
assign t[4861] = t[4860] ^ n[4861];
assign t[4862] = t[4861] ^ n[4862];
assign t[4863] = t[4862] ^ n[4863];
assign t[4864] = t[4863] ^ n[4864];
assign t[4865] = t[4864] ^ n[4865];
assign t[4866] = t[4865] ^ n[4866];
assign t[4867] = t[4866] ^ n[4867];
assign t[4868] = t[4867] ^ n[4868];
assign t[4869] = t[4868] ^ n[4869];
assign t[4870] = t[4869] ^ n[4870];
assign t[4871] = t[4870] ^ n[4871];
assign t[4872] = t[4871] ^ n[4872];
assign t[4873] = t[4872] ^ n[4873];
assign t[4874] = t[4873] ^ n[4874];
assign t[4875] = t[4874] ^ n[4875];
assign t[4876] = t[4875] ^ n[4876];
assign t[4877] = t[4876] ^ n[4877];
assign t[4878] = t[4877] ^ n[4878];
assign t[4879] = t[4878] ^ n[4879];
assign t[4880] = t[4879] ^ n[4880];
assign t[4881] = t[4880] ^ n[4881];
assign t[4882] = t[4881] ^ n[4882];
assign t[4883] = t[4882] ^ n[4883];
assign t[4884] = t[4883] ^ n[4884];
assign t[4885] = t[4884] ^ n[4885];
assign t[4886] = t[4885] ^ n[4886];
assign t[4887] = t[4886] ^ n[4887];
assign t[4888] = t[4887] ^ n[4888];
assign t[4889] = t[4888] ^ n[4889];
assign t[4890] = t[4889] ^ n[4890];
assign t[4891] = t[4890] ^ n[4891];
assign t[4892] = t[4891] ^ n[4892];
assign t[4893] = t[4892] ^ n[4893];
assign t[4894] = t[4893] ^ n[4894];
assign t[4895] = t[4894] ^ n[4895];
assign t[4896] = t[4895] ^ n[4896];
assign t[4897] = t[4896] ^ n[4897];
assign t[4898] = t[4897] ^ n[4898];
assign t[4899] = t[4898] ^ n[4899];
assign t[4900] = t[4899] ^ n[4900];
assign t[4901] = t[4900] ^ n[4901];
assign t[4902] = t[4901] ^ n[4902];
assign t[4903] = t[4902] ^ n[4903];
assign t[4904] = t[4903] ^ n[4904];
assign t[4905] = t[4904] ^ n[4905];
assign t[4906] = t[4905] ^ n[4906];
assign t[4907] = t[4906] ^ n[4907];
assign t[4908] = t[4907] ^ n[4908];
assign t[4909] = t[4908] ^ n[4909];
assign t[4910] = t[4909] ^ n[4910];
assign t[4911] = t[4910] ^ n[4911];
assign t[4912] = t[4911] ^ n[4912];
assign t[4913] = t[4912] ^ n[4913];
assign t[4914] = t[4913] ^ n[4914];
assign t[4915] = t[4914] ^ n[4915];
assign t[4916] = t[4915] ^ n[4916];
assign t[4917] = t[4916] ^ n[4917];
assign t[4918] = t[4917] ^ n[4918];
assign t[4919] = t[4918] ^ n[4919];
assign t[4920] = t[4919] ^ n[4920];
assign t[4921] = t[4920] ^ n[4921];
assign t[4922] = t[4921] ^ n[4922];
assign t[4923] = t[4922] ^ n[4923];
assign t[4924] = t[4923] ^ n[4924];
assign t[4925] = t[4924] ^ n[4925];
assign t[4926] = t[4925] ^ n[4926];
assign t[4927] = t[4926] ^ n[4927];
assign t[4928] = t[4927] ^ n[4928];
assign t[4929] = t[4928] ^ n[4929];
assign t[4930] = t[4929] ^ n[4930];
assign t[4931] = t[4930] ^ n[4931];
assign t[4932] = t[4931] ^ n[4932];
assign t[4933] = t[4932] ^ n[4933];
assign t[4934] = t[4933] ^ n[4934];
assign t[4935] = t[4934] ^ n[4935];
assign t[4936] = t[4935] ^ n[4936];
assign t[4937] = t[4936] ^ n[4937];
assign t[4938] = t[4937] ^ n[4938];
assign t[4939] = t[4938] ^ n[4939];
assign t[4940] = t[4939] ^ n[4940];
assign t[4941] = t[4940] ^ n[4941];
assign t[4942] = t[4941] ^ n[4942];
assign t[4943] = t[4942] ^ n[4943];
assign t[4944] = t[4943] ^ n[4944];
assign t[4945] = t[4944] ^ n[4945];
assign t[4946] = t[4945] ^ n[4946];
assign t[4947] = t[4946] ^ n[4947];
assign t[4948] = t[4947] ^ n[4948];
assign t[4949] = t[4948] ^ n[4949];
assign t[4950] = t[4949] ^ n[4950];
assign t[4951] = t[4950] ^ n[4951];
assign t[4952] = t[4951] ^ n[4952];
assign t[4953] = t[4952] ^ n[4953];
assign t[4954] = t[4953] ^ n[4954];
assign t[4955] = t[4954] ^ n[4955];
assign t[4956] = t[4955] ^ n[4956];
assign t[4957] = t[4956] ^ n[4957];
assign t[4958] = t[4957] ^ n[4958];
assign t[4959] = t[4958] ^ n[4959];
assign t[4960] = t[4959] ^ n[4960];
assign t[4961] = t[4960] ^ n[4961];
assign t[4962] = t[4961] ^ n[4962];
assign t[4963] = t[4962] ^ n[4963];
assign t[4964] = t[4963] ^ n[4964];
assign t[4965] = t[4964] ^ n[4965];
assign t[4966] = t[4965] ^ n[4966];
assign t[4967] = t[4966] ^ n[4967];
assign t[4968] = t[4967] ^ n[4968];
assign t[4969] = t[4968] ^ n[4969];
assign t[4970] = t[4969] ^ n[4970];
assign t[4971] = t[4970] ^ n[4971];
assign t[4972] = t[4971] ^ n[4972];
assign t[4973] = t[4972] ^ n[4973];
assign t[4974] = t[4973] ^ n[4974];
assign t[4975] = t[4974] ^ n[4975];
assign t[4976] = t[4975] ^ n[4976];
assign t[4977] = t[4976] ^ n[4977];
assign t[4978] = t[4977] ^ n[4978];
assign t[4979] = t[4978] ^ n[4979];
assign t[4980] = t[4979] ^ n[4980];
assign t[4981] = t[4980] ^ n[4981];
assign t[4982] = t[4981] ^ n[4982];
assign t[4983] = t[4982] ^ n[4983];
assign t[4984] = t[4983] ^ n[4984];
assign t[4985] = t[4984] ^ n[4985];
assign t[4986] = t[4985] ^ n[4986];
assign t[4987] = t[4986] ^ n[4987];
assign t[4988] = t[4987] ^ n[4988];
assign t[4989] = t[4988] ^ n[4989];
assign t[4990] = t[4989] ^ n[4990];
assign t[4991] = t[4990] ^ n[4991];
assign t[4992] = t[4991] ^ n[4992];
assign t[4993] = t[4992] ^ n[4993];
assign t[4994] = t[4993] ^ n[4994];
assign t[4995] = t[4994] ^ n[4995];
assign t[4996] = t[4995] ^ n[4996];
assign t[4997] = t[4996] ^ n[4997];
assign t[4998] = t[4997] ^ n[4998];
assign t[4999] = t[4998] ^ n[4999];
assign t[5000] = t[4999] ^ n[5000];
assign t[5001] = t[5000] ^ n[5001];
assign t[5002] = t[5001] ^ n[5002];
assign t[5003] = t[5002] ^ n[5003];
assign t[5004] = t[5003] ^ n[5004];
assign t[5005] = t[5004] ^ n[5005];
assign t[5006] = t[5005] ^ n[5006];
assign t[5007] = t[5006] ^ n[5007];
assign t[5008] = t[5007] ^ n[5008];
assign t[5009] = t[5008] ^ n[5009];
assign t[5010] = t[5009] ^ n[5010];
assign t[5011] = t[5010] ^ n[5011];
assign t[5012] = t[5011] ^ n[5012];
assign t[5013] = t[5012] ^ n[5013];
assign t[5014] = t[5013] ^ n[5014];
assign t[5015] = t[5014] ^ n[5015];
assign t[5016] = t[5015] ^ n[5016];
assign t[5017] = t[5016] ^ n[5017];
assign t[5018] = t[5017] ^ n[5018];
assign t[5019] = t[5018] ^ n[5019];
assign t[5020] = t[5019] ^ n[5020];
assign t[5021] = t[5020] ^ n[5021];
assign t[5022] = t[5021] ^ n[5022];
assign t[5023] = t[5022] ^ n[5023];
assign t[5024] = t[5023] ^ n[5024];
assign t[5025] = t[5024] ^ n[5025];
assign t[5026] = t[5025] ^ n[5026];
assign t[5027] = t[5026] ^ n[5027];
assign t[5028] = t[5027] ^ n[5028];
assign t[5029] = t[5028] ^ n[5029];
assign t[5030] = t[5029] ^ n[5030];
assign t[5031] = t[5030] ^ n[5031];
assign t[5032] = t[5031] ^ n[5032];
assign t[5033] = t[5032] ^ n[5033];
assign t[5034] = t[5033] ^ n[5034];
assign t[5035] = t[5034] ^ n[5035];
assign t[5036] = t[5035] ^ n[5036];
assign t[5037] = t[5036] ^ n[5037];
assign t[5038] = t[5037] ^ n[5038];
assign t[5039] = t[5038] ^ n[5039];
assign t[5040] = t[5039] ^ n[5040];
assign t[5041] = t[5040] ^ n[5041];
assign t[5042] = t[5041] ^ n[5042];
assign t[5043] = t[5042] ^ n[5043];
assign t[5044] = t[5043] ^ n[5044];
assign t[5045] = t[5044] ^ n[5045];
assign t[5046] = t[5045] ^ n[5046];
assign t[5047] = t[5046] ^ n[5047];
assign t[5048] = t[5047] ^ n[5048];
assign t[5049] = t[5048] ^ n[5049];
assign t[5050] = t[5049] ^ n[5050];
assign t[5051] = t[5050] ^ n[5051];
assign t[5052] = t[5051] ^ n[5052];
assign t[5053] = t[5052] ^ n[5053];
assign t[5054] = t[5053] ^ n[5054];
assign t[5055] = t[5054] ^ n[5055];
assign t[5056] = t[5055] ^ n[5056];
assign t[5057] = t[5056] ^ n[5057];
assign t[5058] = t[5057] ^ n[5058];
assign t[5059] = t[5058] ^ n[5059];
assign t[5060] = t[5059] ^ n[5060];
assign t[5061] = t[5060] ^ n[5061];
assign t[5062] = t[5061] ^ n[5062];
assign t[5063] = t[5062] ^ n[5063];
assign t[5064] = t[5063] ^ n[5064];
assign t[5065] = t[5064] ^ n[5065];
assign t[5066] = t[5065] ^ n[5066];
assign t[5067] = t[5066] ^ n[5067];
assign t[5068] = t[5067] ^ n[5068];
assign t[5069] = t[5068] ^ n[5069];
assign t[5070] = t[5069] ^ n[5070];
assign t[5071] = t[5070] ^ n[5071];
assign t[5072] = t[5071] ^ n[5072];
assign t[5073] = t[5072] ^ n[5073];
assign t[5074] = t[5073] ^ n[5074];
assign t[5075] = t[5074] ^ n[5075];
assign t[5076] = t[5075] ^ n[5076];
assign t[5077] = t[5076] ^ n[5077];
assign t[5078] = t[5077] ^ n[5078];
assign t[5079] = t[5078] ^ n[5079];
assign t[5080] = t[5079] ^ n[5080];
assign t[5081] = t[5080] ^ n[5081];
assign t[5082] = t[5081] ^ n[5082];
assign t[5083] = t[5082] ^ n[5083];
assign t[5084] = t[5083] ^ n[5084];
assign t[5085] = t[5084] ^ n[5085];
assign t[5086] = t[5085] ^ n[5086];
assign t[5087] = t[5086] ^ n[5087];
assign t[5088] = t[5087] ^ n[5088];
assign t[5089] = t[5088] ^ n[5089];
assign t[5090] = t[5089] ^ n[5090];
assign t[5091] = t[5090] ^ n[5091];
assign t[5092] = t[5091] ^ n[5092];
assign t[5093] = t[5092] ^ n[5093];
assign t[5094] = t[5093] ^ n[5094];
assign t[5095] = t[5094] ^ n[5095];
assign t[5096] = t[5095] ^ n[5096];
assign t[5097] = t[5096] ^ n[5097];
assign t[5098] = t[5097] ^ n[5098];
assign t[5099] = t[5098] ^ n[5099];
assign t[5100] = t[5099] ^ n[5100];
assign t[5101] = t[5100] ^ n[5101];
assign t[5102] = t[5101] ^ n[5102];
assign t[5103] = t[5102] ^ n[5103];
assign t[5104] = t[5103] ^ n[5104];
assign t[5105] = t[5104] ^ n[5105];
assign t[5106] = t[5105] ^ n[5106];
assign t[5107] = t[5106] ^ n[5107];
assign t[5108] = t[5107] ^ n[5108];
assign t[5109] = t[5108] ^ n[5109];
assign t[5110] = t[5109] ^ n[5110];
assign t[5111] = t[5110] ^ n[5111];
assign t[5112] = t[5111] ^ n[5112];
assign t[5113] = t[5112] ^ n[5113];
assign t[5114] = t[5113] ^ n[5114];
assign t[5115] = t[5114] ^ n[5115];
assign t[5116] = t[5115] ^ n[5116];
assign t[5117] = t[5116] ^ n[5117];
assign t[5118] = t[5117] ^ n[5118];
assign t[5119] = t[5118] ^ n[5119];
assign t[5120] = t[5119] ^ n[5120];
assign t[5121] = t[5120] ^ n[5121];
assign t[5122] = t[5121] ^ n[5122];
assign t[5123] = t[5122] ^ n[5123];
assign t[5124] = t[5123] ^ n[5124];
assign t[5125] = t[5124] ^ n[5125];
assign t[5126] = t[5125] ^ n[5126];
assign t[5127] = t[5126] ^ n[5127];
assign t[5128] = t[5127] ^ n[5128];
assign t[5129] = t[5128] ^ n[5129];
assign t[5130] = t[5129] ^ n[5130];
assign t[5131] = t[5130] ^ n[5131];
assign t[5132] = t[5131] ^ n[5132];
assign t[5133] = t[5132] ^ n[5133];
assign t[5134] = t[5133] ^ n[5134];
assign t[5135] = t[5134] ^ n[5135];
assign t[5136] = t[5135] ^ n[5136];
assign t[5137] = t[5136] ^ n[5137];
assign t[5138] = t[5137] ^ n[5138];
assign t[5139] = t[5138] ^ n[5139];
assign t[5140] = t[5139] ^ n[5140];
assign t[5141] = t[5140] ^ n[5141];
assign t[5142] = t[5141] ^ n[5142];
assign t[5143] = t[5142] ^ n[5143];
assign t[5144] = t[5143] ^ n[5144];
assign t[5145] = t[5144] ^ n[5145];
assign t[5146] = t[5145] ^ n[5146];
assign t[5147] = t[5146] ^ n[5147];
assign t[5148] = t[5147] ^ n[5148];
assign t[5149] = t[5148] ^ n[5149];
assign t[5150] = t[5149] ^ n[5150];
assign t[5151] = t[5150] ^ n[5151];
assign t[5152] = t[5151] ^ n[5152];
assign t[5153] = t[5152] ^ n[5153];
assign t[5154] = t[5153] ^ n[5154];
assign t[5155] = t[5154] ^ n[5155];
assign t[5156] = t[5155] ^ n[5156];
assign t[5157] = t[5156] ^ n[5157];
assign t[5158] = t[5157] ^ n[5158];
assign t[5159] = t[5158] ^ n[5159];
assign t[5160] = t[5159] ^ n[5160];
assign t[5161] = t[5160] ^ n[5161];
assign t[5162] = t[5161] ^ n[5162];
assign t[5163] = t[5162] ^ n[5163];
assign t[5164] = t[5163] ^ n[5164];
assign t[5165] = t[5164] ^ n[5165];
assign t[5166] = t[5165] ^ n[5166];
assign t[5167] = t[5166] ^ n[5167];
assign t[5168] = t[5167] ^ n[5168];
assign t[5169] = t[5168] ^ n[5169];
assign t[5170] = t[5169] ^ n[5170];
assign t[5171] = t[5170] ^ n[5171];
assign t[5172] = t[5171] ^ n[5172];
assign t[5173] = t[5172] ^ n[5173];
assign t[5174] = t[5173] ^ n[5174];
assign t[5175] = t[5174] ^ n[5175];
assign t[5176] = t[5175] ^ n[5176];
assign t[5177] = t[5176] ^ n[5177];
assign t[5178] = t[5177] ^ n[5178];
assign t[5179] = t[5178] ^ n[5179];
assign t[5180] = t[5179] ^ n[5180];
assign t[5181] = t[5180] ^ n[5181];
assign t[5182] = t[5181] ^ n[5182];
assign t[5183] = t[5182] ^ n[5183];
assign t[5184] = t[5183] ^ n[5184];
assign t[5185] = t[5184] ^ n[5185];
assign t[5186] = t[5185] ^ n[5186];
assign t[5187] = t[5186] ^ n[5187];
assign t[5188] = t[5187] ^ n[5188];
assign t[5189] = t[5188] ^ n[5189];
assign t[5190] = t[5189] ^ n[5190];
assign t[5191] = t[5190] ^ n[5191];
assign t[5192] = t[5191] ^ n[5192];
assign t[5193] = t[5192] ^ n[5193];
assign t[5194] = t[5193] ^ n[5194];
assign t[5195] = t[5194] ^ n[5195];
assign t[5196] = t[5195] ^ n[5196];
assign t[5197] = t[5196] ^ n[5197];
assign t[5198] = t[5197] ^ n[5198];
assign t[5199] = t[5198] ^ n[5199];
assign t[5200] = t[5199] ^ n[5200];
assign t[5201] = t[5200] ^ n[5201];
assign t[5202] = t[5201] ^ n[5202];
assign t[5203] = t[5202] ^ n[5203];
assign t[5204] = t[5203] ^ n[5204];
assign t[5205] = t[5204] ^ n[5205];
assign t[5206] = t[5205] ^ n[5206];
assign t[5207] = t[5206] ^ n[5207];
assign t[5208] = t[5207] ^ n[5208];
assign t[5209] = t[5208] ^ n[5209];
assign t[5210] = t[5209] ^ n[5210];
assign t[5211] = t[5210] ^ n[5211];
assign t[5212] = t[5211] ^ n[5212];
assign t[5213] = t[5212] ^ n[5213];
assign t[5214] = t[5213] ^ n[5214];
assign t[5215] = t[5214] ^ n[5215];
assign t[5216] = t[5215] ^ n[5216];
assign t[5217] = t[5216] ^ n[5217];
assign t[5218] = t[5217] ^ n[5218];
assign t[5219] = t[5218] ^ n[5219];
assign t[5220] = t[5219] ^ n[5220];
assign t[5221] = t[5220] ^ n[5221];
assign t[5222] = t[5221] ^ n[5222];
assign t[5223] = t[5222] ^ n[5223];
assign t[5224] = t[5223] ^ n[5224];
assign t[5225] = t[5224] ^ n[5225];
assign t[5226] = t[5225] ^ n[5226];
assign t[5227] = t[5226] ^ n[5227];
assign t[5228] = t[5227] ^ n[5228];
assign t[5229] = t[5228] ^ n[5229];
assign t[5230] = t[5229] ^ n[5230];
assign t[5231] = t[5230] ^ n[5231];
assign t[5232] = t[5231] ^ n[5232];
assign t[5233] = t[5232] ^ n[5233];
assign t[5234] = t[5233] ^ n[5234];
assign t[5235] = t[5234] ^ n[5235];
assign t[5236] = t[5235] ^ n[5236];
assign t[5237] = t[5236] ^ n[5237];
assign t[5238] = t[5237] ^ n[5238];
assign t[5239] = t[5238] ^ n[5239];
assign t[5240] = t[5239] ^ n[5240];
assign t[5241] = t[5240] ^ n[5241];
assign t[5242] = t[5241] ^ n[5242];
assign t[5243] = t[5242] ^ n[5243];
assign t[5244] = t[5243] ^ n[5244];
assign t[5245] = t[5244] ^ n[5245];
assign t[5246] = t[5245] ^ n[5246];
assign t[5247] = t[5246] ^ n[5247];
assign t[5248] = t[5247] ^ n[5248];
assign t[5249] = t[5248] ^ n[5249];
assign t[5250] = t[5249] ^ n[5250];
assign t[5251] = t[5250] ^ n[5251];
assign t[5252] = t[5251] ^ n[5252];
assign t[5253] = t[5252] ^ n[5253];
assign t[5254] = t[5253] ^ n[5254];
assign t[5255] = t[5254] ^ n[5255];
assign t[5256] = t[5255] ^ n[5256];
assign t[5257] = t[5256] ^ n[5257];
assign t[5258] = t[5257] ^ n[5258];
assign t[5259] = t[5258] ^ n[5259];
assign t[5260] = t[5259] ^ n[5260];
assign t[5261] = t[5260] ^ n[5261];
assign t[5262] = t[5261] ^ n[5262];
assign t[5263] = t[5262] ^ n[5263];
assign t[5264] = t[5263] ^ n[5264];
assign t[5265] = t[5264] ^ n[5265];
assign t[5266] = t[5265] ^ n[5266];
assign t[5267] = t[5266] ^ n[5267];
assign t[5268] = t[5267] ^ n[5268];
assign t[5269] = t[5268] ^ n[5269];
assign t[5270] = t[5269] ^ n[5270];
assign t[5271] = t[5270] ^ n[5271];
assign t[5272] = t[5271] ^ n[5272];
assign t[5273] = t[5272] ^ n[5273];
assign t[5274] = t[5273] ^ n[5274];
assign t[5275] = t[5274] ^ n[5275];
assign t[5276] = t[5275] ^ n[5276];
assign t[5277] = t[5276] ^ n[5277];
assign t[5278] = t[5277] ^ n[5278];
assign t[5279] = t[5278] ^ n[5279];
assign t[5280] = t[5279] ^ n[5280];
assign t[5281] = t[5280] ^ n[5281];
assign t[5282] = t[5281] ^ n[5282];
assign t[5283] = t[5282] ^ n[5283];
assign t[5284] = t[5283] ^ n[5284];
assign t[5285] = t[5284] ^ n[5285];
assign t[5286] = t[5285] ^ n[5286];
assign t[5287] = t[5286] ^ n[5287];
assign t[5288] = t[5287] ^ n[5288];
assign t[5289] = t[5288] ^ n[5289];
assign t[5290] = t[5289] ^ n[5290];
assign t[5291] = t[5290] ^ n[5291];
assign t[5292] = t[5291] ^ n[5292];
assign t[5293] = t[5292] ^ n[5293];
assign t[5294] = t[5293] ^ n[5294];
assign t[5295] = t[5294] ^ n[5295];
assign t[5296] = t[5295] ^ n[5296];
assign t[5297] = t[5296] ^ n[5297];
assign t[5298] = t[5297] ^ n[5298];
assign t[5299] = t[5298] ^ n[5299];
assign t[5300] = t[5299] ^ n[5300];
assign t[5301] = t[5300] ^ n[5301];
assign t[5302] = t[5301] ^ n[5302];
assign t[5303] = t[5302] ^ n[5303];
assign t[5304] = t[5303] ^ n[5304];
assign t[5305] = t[5304] ^ n[5305];
assign t[5306] = t[5305] ^ n[5306];
assign t[5307] = t[5306] ^ n[5307];
assign t[5308] = t[5307] ^ n[5308];
assign t[5309] = t[5308] ^ n[5309];
assign t[5310] = t[5309] ^ n[5310];
assign t[5311] = t[5310] ^ n[5311];
assign t[5312] = t[5311] ^ n[5312];
assign t[5313] = t[5312] ^ n[5313];
assign t[5314] = t[5313] ^ n[5314];
assign t[5315] = t[5314] ^ n[5315];
assign t[5316] = t[5315] ^ n[5316];
assign t[5317] = t[5316] ^ n[5317];
assign t[5318] = t[5317] ^ n[5318];
assign t[5319] = t[5318] ^ n[5319];
assign t[5320] = t[5319] ^ n[5320];
assign t[5321] = t[5320] ^ n[5321];
assign t[5322] = t[5321] ^ n[5322];
assign t[5323] = t[5322] ^ n[5323];
assign t[5324] = t[5323] ^ n[5324];
assign t[5325] = t[5324] ^ n[5325];
assign t[5326] = t[5325] ^ n[5326];
assign t[5327] = t[5326] ^ n[5327];
assign t[5328] = t[5327] ^ n[5328];
assign t[5329] = t[5328] ^ n[5329];
assign t[5330] = t[5329] ^ n[5330];
assign t[5331] = t[5330] ^ n[5331];
assign t[5332] = t[5331] ^ n[5332];
assign t[5333] = t[5332] ^ n[5333];
assign t[5334] = t[5333] ^ n[5334];
assign t[5335] = t[5334] ^ n[5335];
assign t[5336] = t[5335] ^ n[5336];
assign t[5337] = t[5336] ^ n[5337];
assign t[5338] = t[5337] ^ n[5338];
assign t[5339] = t[5338] ^ n[5339];
assign t[5340] = t[5339] ^ n[5340];
assign t[5341] = t[5340] ^ n[5341];
assign t[5342] = t[5341] ^ n[5342];
assign t[5343] = t[5342] ^ n[5343];
assign t[5344] = t[5343] ^ n[5344];
assign t[5345] = t[5344] ^ n[5345];
assign t[5346] = t[5345] ^ n[5346];
assign t[5347] = t[5346] ^ n[5347];
assign t[5348] = t[5347] ^ n[5348];
assign t[5349] = t[5348] ^ n[5349];
assign t[5350] = t[5349] ^ n[5350];
assign t[5351] = t[5350] ^ n[5351];
assign t[5352] = t[5351] ^ n[5352];
assign t[5353] = t[5352] ^ n[5353];
assign t[5354] = t[5353] ^ n[5354];
assign t[5355] = t[5354] ^ n[5355];
assign t[5356] = t[5355] ^ n[5356];
assign t[5357] = t[5356] ^ n[5357];
assign t[5358] = t[5357] ^ n[5358];
assign t[5359] = t[5358] ^ n[5359];
assign t[5360] = t[5359] ^ n[5360];
assign t[5361] = t[5360] ^ n[5361];
assign t[5362] = t[5361] ^ n[5362];
assign t[5363] = t[5362] ^ n[5363];
assign t[5364] = t[5363] ^ n[5364];
assign t[5365] = t[5364] ^ n[5365];
assign t[5366] = t[5365] ^ n[5366];
assign t[5367] = t[5366] ^ n[5367];
assign t[5368] = t[5367] ^ n[5368];
assign t[5369] = t[5368] ^ n[5369];
assign t[5370] = t[5369] ^ n[5370];
assign t[5371] = t[5370] ^ n[5371];
assign t[5372] = t[5371] ^ n[5372];
assign t[5373] = t[5372] ^ n[5373];
assign t[5374] = t[5373] ^ n[5374];
assign t[5375] = t[5374] ^ n[5375];
assign t[5376] = t[5375] ^ n[5376];
assign t[5377] = t[5376] ^ n[5377];
assign t[5378] = t[5377] ^ n[5378];
assign t[5379] = t[5378] ^ n[5379];
assign t[5380] = t[5379] ^ n[5380];
assign t[5381] = t[5380] ^ n[5381];
assign t[5382] = t[5381] ^ n[5382];
assign t[5383] = t[5382] ^ n[5383];
assign t[5384] = t[5383] ^ n[5384];
assign t[5385] = t[5384] ^ n[5385];
assign t[5386] = t[5385] ^ n[5386];
assign t[5387] = t[5386] ^ n[5387];
assign t[5388] = t[5387] ^ n[5388];
assign t[5389] = t[5388] ^ n[5389];
assign t[5390] = t[5389] ^ n[5390];
assign t[5391] = t[5390] ^ n[5391];
assign t[5392] = t[5391] ^ n[5392];
assign t[5393] = t[5392] ^ n[5393];
assign t[5394] = t[5393] ^ n[5394];
assign t[5395] = t[5394] ^ n[5395];
assign t[5396] = t[5395] ^ n[5396];
assign t[5397] = t[5396] ^ n[5397];
assign t[5398] = t[5397] ^ n[5398];
assign t[5399] = t[5398] ^ n[5399];
assign t[5400] = t[5399] ^ n[5400];
assign t[5401] = t[5400] ^ n[5401];
assign t[5402] = t[5401] ^ n[5402];
assign t[5403] = t[5402] ^ n[5403];
assign t[5404] = t[5403] ^ n[5404];
assign t[5405] = t[5404] ^ n[5405];
assign t[5406] = t[5405] ^ n[5406];
assign t[5407] = t[5406] ^ n[5407];
assign t[5408] = t[5407] ^ n[5408];
assign t[5409] = t[5408] ^ n[5409];
assign t[5410] = t[5409] ^ n[5410];
assign t[5411] = t[5410] ^ n[5411];
assign t[5412] = t[5411] ^ n[5412];
assign t[5413] = t[5412] ^ n[5413];
assign t[5414] = t[5413] ^ n[5414];
assign t[5415] = t[5414] ^ n[5415];
assign t[5416] = t[5415] ^ n[5416];
assign t[5417] = t[5416] ^ n[5417];
assign t[5418] = t[5417] ^ n[5418];
assign t[5419] = t[5418] ^ n[5419];
assign t[5420] = t[5419] ^ n[5420];
assign t[5421] = t[5420] ^ n[5421];
assign t[5422] = t[5421] ^ n[5422];
assign t[5423] = t[5422] ^ n[5423];
assign t[5424] = t[5423] ^ n[5424];
assign t[5425] = t[5424] ^ n[5425];
assign t[5426] = t[5425] ^ n[5426];
assign t[5427] = t[5426] ^ n[5427];
assign t[5428] = t[5427] ^ n[5428];
assign t[5429] = t[5428] ^ n[5429];
assign t[5430] = t[5429] ^ n[5430];
assign t[5431] = t[5430] ^ n[5431];
assign t[5432] = t[5431] ^ n[5432];
assign t[5433] = t[5432] ^ n[5433];
assign t[5434] = t[5433] ^ n[5434];
assign t[5435] = t[5434] ^ n[5435];
assign t[5436] = t[5435] ^ n[5436];
assign t[5437] = t[5436] ^ n[5437];
assign t[5438] = t[5437] ^ n[5438];
assign t[5439] = t[5438] ^ n[5439];
assign t[5440] = t[5439] ^ n[5440];
assign t[5441] = t[5440] ^ n[5441];
assign t[5442] = t[5441] ^ n[5442];
assign t[5443] = t[5442] ^ n[5443];
assign t[5444] = t[5443] ^ n[5444];
assign t[5445] = t[5444] ^ n[5445];
assign t[5446] = t[5445] ^ n[5446];
assign t[5447] = t[5446] ^ n[5447];
assign t[5448] = t[5447] ^ n[5448];
assign t[5449] = t[5448] ^ n[5449];
assign t[5450] = t[5449] ^ n[5450];
assign t[5451] = t[5450] ^ n[5451];
assign t[5452] = t[5451] ^ n[5452];
assign t[5453] = t[5452] ^ n[5453];
assign t[5454] = t[5453] ^ n[5454];
assign t[5455] = t[5454] ^ n[5455];
assign t[5456] = t[5455] ^ n[5456];
assign t[5457] = t[5456] ^ n[5457];
assign t[5458] = t[5457] ^ n[5458];
assign t[5459] = t[5458] ^ n[5459];
assign t[5460] = t[5459] ^ n[5460];
assign t[5461] = t[5460] ^ n[5461];
assign t[5462] = t[5461] ^ n[5462];
assign t[5463] = t[5462] ^ n[5463];
assign t[5464] = t[5463] ^ n[5464];
assign t[5465] = t[5464] ^ n[5465];
assign t[5466] = t[5465] ^ n[5466];
assign t[5467] = t[5466] ^ n[5467];
assign t[5468] = t[5467] ^ n[5468];
assign t[5469] = t[5468] ^ n[5469];
assign t[5470] = t[5469] ^ n[5470];
assign t[5471] = t[5470] ^ n[5471];
assign t[5472] = t[5471] ^ n[5472];
assign t[5473] = t[5472] ^ n[5473];
assign t[5474] = t[5473] ^ n[5474];
assign t[5475] = t[5474] ^ n[5475];
assign t[5476] = t[5475] ^ n[5476];
assign t[5477] = t[5476] ^ n[5477];
assign t[5478] = t[5477] ^ n[5478];
assign t[5479] = t[5478] ^ n[5479];
assign t[5480] = t[5479] ^ n[5480];
assign t[5481] = t[5480] ^ n[5481];
assign t[5482] = t[5481] ^ n[5482];
assign t[5483] = t[5482] ^ n[5483];
assign t[5484] = t[5483] ^ n[5484];
assign t[5485] = t[5484] ^ n[5485];
assign t[5486] = t[5485] ^ n[5486];
assign t[5487] = t[5486] ^ n[5487];
assign t[5488] = t[5487] ^ n[5488];
assign t[5489] = t[5488] ^ n[5489];
assign t[5490] = t[5489] ^ n[5490];
assign t[5491] = t[5490] ^ n[5491];
assign t[5492] = t[5491] ^ n[5492];
assign t[5493] = t[5492] ^ n[5493];
assign t[5494] = t[5493] ^ n[5494];
assign t[5495] = t[5494] ^ n[5495];
assign t[5496] = t[5495] ^ n[5496];
assign t[5497] = t[5496] ^ n[5497];
assign t[5498] = t[5497] ^ n[5498];
assign t[5499] = t[5498] ^ n[5499];
assign t[5500] = t[5499] ^ n[5500];
assign t[5501] = t[5500] ^ n[5501];
assign t[5502] = t[5501] ^ n[5502];
assign t[5503] = t[5502] ^ n[5503];
assign t[5504] = t[5503] ^ n[5504];
assign t[5505] = t[5504] ^ n[5505];
assign t[5506] = t[5505] ^ n[5506];
assign t[5507] = t[5506] ^ n[5507];
assign t[5508] = t[5507] ^ n[5508];
assign t[5509] = t[5508] ^ n[5509];
assign t[5510] = t[5509] ^ n[5510];
assign t[5511] = t[5510] ^ n[5511];
assign t[5512] = t[5511] ^ n[5512];
assign t[5513] = t[5512] ^ n[5513];
assign t[5514] = t[5513] ^ n[5514];
assign t[5515] = t[5514] ^ n[5515];
assign t[5516] = t[5515] ^ n[5516];
assign t[5517] = t[5516] ^ n[5517];
assign t[5518] = t[5517] ^ n[5518];
assign t[5519] = t[5518] ^ n[5519];
assign t[5520] = t[5519] ^ n[5520];
assign t[5521] = t[5520] ^ n[5521];
assign t[5522] = t[5521] ^ n[5522];
assign t[5523] = t[5522] ^ n[5523];
assign t[5524] = t[5523] ^ n[5524];
assign t[5525] = t[5524] ^ n[5525];
assign t[5526] = t[5525] ^ n[5526];
assign t[5527] = t[5526] ^ n[5527];
assign t[5528] = t[5527] ^ n[5528];
assign t[5529] = t[5528] ^ n[5529];
assign t[5530] = t[5529] ^ n[5530];
assign t[5531] = t[5530] ^ n[5531];
assign t[5532] = t[5531] ^ n[5532];
assign t[5533] = t[5532] ^ n[5533];
assign t[5534] = t[5533] ^ n[5534];
assign t[5535] = t[5534] ^ n[5535];
assign t[5536] = t[5535] ^ n[5536];
assign t[5537] = t[5536] ^ n[5537];
assign t[5538] = t[5537] ^ n[5538];
assign t[5539] = t[5538] ^ n[5539];
assign t[5540] = t[5539] ^ n[5540];
assign t[5541] = t[5540] ^ n[5541];
assign t[5542] = t[5541] ^ n[5542];
assign t[5543] = t[5542] ^ n[5543];
assign t[5544] = t[5543] ^ n[5544];
assign t[5545] = t[5544] ^ n[5545];
assign t[5546] = t[5545] ^ n[5546];
assign t[5547] = t[5546] ^ n[5547];
assign t[5548] = t[5547] ^ n[5548];
assign t[5549] = t[5548] ^ n[5549];
assign t[5550] = t[5549] ^ n[5550];
assign t[5551] = t[5550] ^ n[5551];
assign t[5552] = t[5551] ^ n[5552];
assign t[5553] = t[5552] ^ n[5553];
assign t[5554] = t[5553] ^ n[5554];
assign t[5555] = t[5554] ^ n[5555];
assign t[5556] = t[5555] ^ n[5556];
assign t[5557] = t[5556] ^ n[5557];
assign t[5558] = t[5557] ^ n[5558];
assign t[5559] = t[5558] ^ n[5559];
assign t[5560] = t[5559] ^ n[5560];
assign t[5561] = t[5560] ^ n[5561];
assign t[5562] = t[5561] ^ n[5562];
assign t[5563] = t[5562] ^ n[5563];
assign t[5564] = t[5563] ^ n[5564];
assign t[5565] = t[5564] ^ n[5565];
assign t[5566] = t[5565] ^ n[5566];
assign t[5567] = t[5566] ^ n[5567];
assign t[5568] = t[5567] ^ n[5568];
assign t[5569] = t[5568] ^ n[5569];
assign t[5570] = t[5569] ^ n[5570];
assign t[5571] = t[5570] ^ n[5571];
assign t[5572] = t[5571] ^ n[5572];
assign t[5573] = t[5572] ^ n[5573];
assign t[5574] = t[5573] ^ n[5574];
assign t[5575] = t[5574] ^ n[5575];
assign t[5576] = t[5575] ^ n[5576];
assign t[5577] = t[5576] ^ n[5577];
assign t[5578] = t[5577] ^ n[5578];
assign t[5579] = t[5578] ^ n[5579];
assign t[5580] = t[5579] ^ n[5580];
assign t[5581] = t[5580] ^ n[5581];
assign t[5582] = t[5581] ^ n[5582];
assign t[5583] = t[5582] ^ n[5583];
assign t[5584] = t[5583] ^ n[5584];
assign t[5585] = t[5584] ^ n[5585];
assign t[5586] = t[5585] ^ n[5586];
assign t[5587] = t[5586] ^ n[5587];
assign t[5588] = t[5587] ^ n[5588];
assign t[5589] = t[5588] ^ n[5589];
assign t[5590] = t[5589] ^ n[5590];
assign t[5591] = t[5590] ^ n[5591];
assign t[5592] = t[5591] ^ n[5592];
assign t[5593] = t[5592] ^ n[5593];
assign t[5594] = t[5593] ^ n[5594];
assign t[5595] = t[5594] ^ n[5595];
assign t[5596] = t[5595] ^ n[5596];
assign t[5597] = t[5596] ^ n[5597];
assign t[5598] = t[5597] ^ n[5598];
assign t[5599] = t[5598] ^ n[5599];
assign t[5600] = t[5599] ^ n[5600];
assign t[5601] = t[5600] ^ n[5601];
assign t[5602] = t[5601] ^ n[5602];
assign t[5603] = t[5602] ^ n[5603];
assign t[5604] = t[5603] ^ n[5604];
assign t[5605] = t[5604] ^ n[5605];
assign t[5606] = t[5605] ^ n[5606];
assign t[5607] = t[5606] ^ n[5607];
assign t[5608] = t[5607] ^ n[5608];
assign t[5609] = t[5608] ^ n[5609];
assign t[5610] = t[5609] ^ n[5610];
assign t[5611] = t[5610] ^ n[5611];
assign t[5612] = t[5611] ^ n[5612];
assign t[5613] = t[5612] ^ n[5613];
assign t[5614] = t[5613] ^ n[5614];
assign t[5615] = t[5614] ^ n[5615];
assign t[5616] = t[5615] ^ n[5616];
assign t[5617] = t[5616] ^ n[5617];
assign t[5618] = t[5617] ^ n[5618];
assign t[5619] = t[5618] ^ n[5619];
assign t[5620] = t[5619] ^ n[5620];
assign t[5621] = t[5620] ^ n[5621];
assign t[5622] = t[5621] ^ n[5622];
assign t[5623] = t[5622] ^ n[5623];
assign t[5624] = t[5623] ^ n[5624];
assign t[5625] = t[5624] ^ n[5625];
assign t[5626] = t[5625] ^ n[5626];
assign t[5627] = t[5626] ^ n[5627];
assign t[5628] = t[5627] ^ n[5628];
assign t[5629] = t[5628] ^ n[5629];
assign t[5630] = t[5629] ^ n[5630];
assign t[5631] = t[5630] ^ n[5631];
assign t[5632] = t[5631] ^ n[5632];
assign t[5633] = t[5632] ^ n[5633];
assign t[5634] = t[5633] ^ n[5634];
assign t[5635] = t[5634] ^ n[5635];
assign t[5636] = t[5635] ^ n[5636];
assign t[5637] = t[5636] ^ n[5637];
assign t[5638] = t[5637] ^ n[5638];
assign t[5639] = t[5638] ^ n[5639];
assign t[5640] = t[5639] ^ n[5640];
assign t[5641] = t[5640] ^ n[5641];
assign t[5642] = t[5641] ^ n[5642];
assign t[5643] = t[5642] ^ n[5643];
assign t[5644] = t[5643] ^ n[5644];
assign t[5645] = t[5644] ^ n[5645];
assign t[5646] = t[5645] ^ n[5646];
assign t[5647] = t[5646] ^ n[5647];
assign t[5648] = t[5647] ^ n[5648];
assign t[5649] = t[5648] ^ n[5649];
assign t[5650] = t[5649] ^ n[5650];
assign t[5651] = t[5650] ^ n[5651];
assign t[5652] = t[5651] ^ n[5652];
assign t[5653] = t[5652] ^ n[5653];
assign t[5654] = t[5653] ^ n[5654];
assign t[5655] = t[5654] ^ n[5655];
assign t[5656] = t[5655] ^ n[5656];
assign t[5657] = t[5656] ^ n[5657];
assign t[5658] = t[5657] ^ n[5658];
assign t[5659] = t[5658] ^ n[5659];
assign t[5660] = t[5659] ^ n[5660];
assign t[5661] = t[5660] ^ n[5661];
assign t[5662] = t[5661] ^ n[5662];
assign t[5663] = t[5662] ^ n[5663];
assign t[5664] = t[5663] ^ n[5664];
assign t[5665] = t[5664] ^ n[5665];
assign t[5666] = t[5665] ^ n[5666];
assign t[5667] = t[5666] ^ n[5667];
assign t[5668] = t[5667] ^ n[5668];
assign t[5669] = t[5668] ^ n[5669];
assign t[5670] = t[5669] ^ n[5670];
assign t[5671] = t[5670] ^ n[5671];
assign t[5672] = t[5671] ^ n[5672];
assign t[5673] = t[5672] ^ n[5673];
assign t[5674] = t[5673] ^ n[5674];
assign t[5675] = t[5674] ^ n[5675];
assign t[5676] = t[5675] ^ n[5676];
assign t[5677] = t[5676] ^ n[5677];
assign t[5678] = t[5677] ^ n[5678];
assign t[5679] = t[5678] ^ n[5679];
assign t[5680] = t[5679] ^ n[5680];
assign t[5681] = t[5680] ^ n[5681];
assign t[5682] = t[5681] ^ n[5682];
assign t[5683] = t[5682] ^ n[5683];
assign t[5684] = t[5683] ^ n[5684];
assign t[5685] = t[5684] ^ n[5685];
assign t[5686] = t[5685] ^ n[5686];
assign t[5687] = t[5686] ^ n[5687];
assign t[5688] = t[5687] ^ n[5688];
assign t[5689] = t[5688] ^ n[5689];
assign t[5690] = t[5689] ^ n[5690];
assign t[5691] = t[5690] ^ n[5691];
assign t[5692] = t[5691] ^ n[5692];
assign t[5693] = t[5692] ^ n[5693];
assign t[5694] = t[5693] ^ n[5694];
assign t[5695] = t[5694] ^ n[5695];
assign t[5696] = t[5695] ^ n[5696];
assign t[5697] = t[5696] ^ n[5697];
assign t[5698] = t[5697] ^ n[5698];
assign t[5699] = t[5698] ^ n[5699];
assign t[5700] = t[5699] ^ n[5700];
assign t[5701] = t[5700] ^ n[5701];
assign t[5702] = t[5701] ^ n[5702];
assign t[5703] = t[5702] ^ n[5703];
assign t[5704] = t[5703] ^ n[5704];
assign t[5705] = t[5704] ^ n[5705];
assign t[5706] = t[5705] ^ n[5706];
assign t[5707] = t[5706] ^ n[5707];
assign t[5708] = t[5707] ^ n[5708];
assign t[5709] = t[5708] ^ n[5709];
assign t[5710] = t[5709] ^ n[5710];
assign t[5711] = t[5710] ^ n[5711];
assign t[5712] = t[5711] ^ n[5712];
assign t[5713] = t[5712] ^ n[5713];
assign t[5714] = t[5713] ^ n[5714];
assign t[5715] = t[5714] ^ n[5715];
assign t[5716] = t[5715] ^ n[5716];
assign t[5717] = t[5716] ^ n[5717];
assign t[5718] = t[5717] ^ n[5718];
assign t[5719] = t[5718] ^ n[5719];
assign t[5720] = t[5719] ^ n[5720];
assign t[5721] = t[5720] ^ n[5721];
assign t[5722] = t[5721] ^ n[5722];
assign t[5723] = t[5722] ^ n[5723];
assign t[5724] = t[5723] ^ n[5724];
assign t[5725] = t[5724] ^ n[5725];
assign t[5726] = t[5725] ^ n[5726];
assign t[5727] = t[5726] ^ n[5727];
assign t[5728] = t[5727] ^ n[5728];
assign t[5729] = t[5728] ^ n[5729];
assign t[5730] = t[5729] ^ n[5730];
assign t[5731] = t[5730] ^ n[5731];
assign t[5732] = t[5731] ^ n[5732];
assign t[5733] = t[5732] ^ n[5733];
assign t[5734] = t[5733] ^ n[5734];
assign t[5735] = t[5734] ^ n[5735];
assign t[5736] = t[5735] ^ n[5736];
assign t[5737] = t[5736] ^ n[5737];
assign t[5738] = t[5737] ^ n[5738];
assign t[5739] = t[5738] ^ n[5739];
assign t[5740] = t[5739] ^ n[5740];
assign t[5741] = t[5740] ^ n[5741];
assign t[5742] = t[5741] ^ n[5742];
assign t[5743] = t[5742] ^ n[5743];
assign t[5744] = t[5743] ^ n[5744];
assign t[5745] = t[5744] ^ n[5745];
assign t[5746] = t[5745] ^ n[5746];
assign t[5747] = t[5746] ^ n[5747];
assign t[5748] = t[5747] ^ n[5748];
assign t[5749] = t[5748] ^ n[5749];
assign t[5750] = t[5749] ^ n[5750];
assign t[5751] = t[5750] ^ n[5751];
assign t[5752] = t[5751] ^ n[5752];
assign t[5753] = t[5752] ^ n[5753];
assign t[5754] = t[5753] ^ n[5754];
assign t[5755] = t[5754] ^ n[5755];
assign t[5756] = t[5755] ^ n[5756];
assign t[5757] = t[5756] ^ n[5757];
assign t[5758] = t[5757] ^ n[5758];
assign t[5759] = t[5758] ^ n[5759];
assign t[5760] = t[5759] ^ n[5760];
assign t[5761] = t[5760] ^ n[5761];
assign t[5762] = t[5761] ^ n[5762];
assign t[5763] = t[5762] ^ n[5763];
assign t[5764] = t[5763] ^ n[5764];
assign t[5765] = t[5764] ^ n[5765];
assign t[5766] = t[5765] ^ n[5766];
assign t[5767] = t[5766] ^ n[5767];
assign t[5768] = t[5767] ^ n[5768];
assign t[5769] = t[5768] ^ n[5769];
assign t[5770] = t[5769] ^ n[5770];
assign t[5771] = t[5770] ^ n[5771];
assign t[5772] = t[5771] ^ n[5772];
assign t[5773] = t[5772] ^ n[5773];
assign t[5774] = t[5773] ^ n[5774];
assign t[5775] = t[5774] ^ n[5775];
assign t[5776] = t[5775] ^ n[5776];
assign t[5777] = t[5776] ^ n[5777];
assign t[5778] = t[5777] ^ n[5778];
assign t[5779] = t[5778] ^ n[5779];
assign t[5780] = t[5779] ^ n[5780];
assign t[5781] = t[5780] ^ n[5781];
assign t[5782] = t[5781] ^ n[5782];
assign t[5783] = t[5782] ^ n[5783];
assign t[5784] = t[5783] ^ n[5784];
assign t[5785] = t[5784] ^ n[5785];
assign t[5786] = t[5785] ^ n[5786];
assign t[5787] = t[5786] ^ n[5787];
assign t[5788] = t[5787] ^ n[5788];
assign t[5789] = t[5788] ^ n[5789];
assign t[5790] = t[5789] ^ n[5790];
assign t[5791] = t[5790] ^ n[5791];
assign t[5792] = t[5791] ^ n[5792];
assign t[5793] = t[5792] ^ n[5793];
assign t[5794] = t[5793] ^ n[5794];
assign t[5795] = t[5794] ^ n[5795];
assign t[5796] = t[5795] ^ n[5796];
assign t[5797] = t[5796] ^ n[5797];
assign t[5798] = t[5797] ^ n[5798];
assign t[5799] = t[5798] ^ n[5799];
assign t[5800] = t[5799] ^ n[5800];
assign t[5801] = t[5800] ^ n[5801];
assign t[5802] = t[5801] ^ n[5802];
assign t[5803] = t[5802] ^ n[5803];
assign t[5804] = t[5803] ^ n[5804];
assign t[5805] = t[5804] ^ n[5805];
assign t[5806] = t[5805] ^ n[5806];
assign t[5807] = t[5806] ^ n[5807];
assign t[5808] = t[5807] ^ n[5808];
assign t[5809] = t[5808] ^ n[5809];
assign t[5810] = t[5809] ^ n[5810];
assign t[5811] = t[5810] ^ n[5811];
assign t[5812] = t[5811] ^ n[5812];
assign t[5813] = t[5812] ^ n[5813];
assign t[5814] = t[5813] ^ n[5814];
assign t[5815] = t[5814] ^ n[5815];
assign t[5816] = t[5815] ^ n[5816];
assign t[5817] = t[5816] ^ n[5817];
assign t[5818] = t[5817] ^ n[5818];
assign t[5819] = t[5818] ^ n[5819];
assign t[5820] = t[5819] ^ n[5820];
assign t[5821] = t[5820] ^ n[5821];
assign t[5822] = t[5821] ^ n[5822];
assign t[5823] = t[5822] ^ n[5823];
assign t[5824] = t[5823] ^ n[5824];
assign t[5825] = t[5824] ^ n[5825];
assign t[5826] = t[5825] ^ n[5826];
assign t[5827] = t[5826] ^ n[5827];
assign t[5828] = t[5827] ^ n[5828];
assign t[5829] = t[5828] ^ n[5829];
assign t[5830] = t[5829] ^ n[5830];
assign t[5831] = t[5830] ^ n[5831];
assign t[5832] = t[5831] ^ n[5832];
assign t[5833] = t[5832] ^ n[5833];
assign t[5834] = t[5833] ^ n[5834];
assign t[5835] = t[5834] ^ n[5835];
assign t[5836] = t[5835] ^ n[5836];
assign t[5837] = t[5836] ^ n[5837];
assign t[5838] = t[5837] ^ n[5838];
assign t[5839] = t[5838] ^ n[5839];
assign t[5840] = t[5839] ^ n[5840];
assign t[5841] = t[5840] ^ n[5841];
assign t[5842] = t[5841] ^ n[5842];
assign t[5843] = t[5842] ^ n[5843];
assign t[5844] = t[5843] ^ n[5844];
assign t[5845] = t[5844] ^ n[5845];
assign t[5846] = t[5845] ^ n[5846];
assign t[5847] = t[5846] ^ n[5847];
assign t[5848] = t[5847] ^ n[5848];
assign t[5849] = t[5848] ^ n[5849];
assign t[5850] = t[5849] ^ n[5850];
assign t[5851] = t[5850] ^ n[5851];
assign t[5852] = t[5851] ^ n[5852];
assign t[5853] = t[5852] ^ n[5853];
assign t[5854] = t[5853] ^ n[5854];
assign t[5855] = t[5854] ^ n[5855];
assign t[5856] = t[5855] ^ n[5856];
assign t[5857] = t[5856] ^ n[5857];
assign t[5858] = t[5857] ^ n[5858];
assign t[5859] = t[5858] ^ n[5859];
assign t[5860] = t[5859] ^ n[5860];
assign t[5861] = t[5860] ^ n[5861];
assign t[5862] = t[5861] ^ n[5862];
assign t[5863] = t[5862] ^ n[5863];
assign t[5864] = t[5863] ^ n[5864];
assign t[5865] = t[5864] ^ n[5865];
assign t[5866] = t[5865] ^ n[5866];
assign t[5867] = t[5866] ^ n[5867];
assign t[5868] = t[5867] ^ n[5868];
assign t[5869] = t[5868] ^ n[5869];
assign t[5870] = t[5869] ^ n[5870];
assign t[5871] = t[5870] ^ n[5871];
assign t[5872] = t[5871] ^ n[5872];
assign t[5873] = t[5872] ^ n[5873];
assign t[5874] = t[5873] ^ n[5874];
assign t[5875] = t[5874] ^ n[5875];
assign t[5876] = t[5875] ^ n[5876];
assign t[5877] = t[5876] ^ n[5877];
assign t[5878] = t[5877] ^ n[5878];
assign t[5879] = t[5878] ^ n[5879];
assign t[5880] = t[5879] ^ n[5880];
assign t[5881] = t[5880] ^ n[5881];
assign t[5882] = t[5881] ^ n[5882];
assign t[5883] = t[5882] ^ n[5883];
assign t[5884] = t[5883] ^ n[5884];
assign t[5885] = t[5884] ^ n[5885];
assign t[5886] = t[5885] ^ n[5886];
assign t[5887] = t[5886] ^ n[5887];
assign t[5888] = t[5887] ^ n[5888];
assign t[5889] = t[5888] ^ n[5889];
assign t[5890] = t[5889] ^ n[5890];
assign t[5891] = t[5890] ^ n[5891];
assign t[5892] = t[5891] ^ n[5892];
assign t[5893] = t[5892] ^ n[5893];
assign t[5894] = t[5893] ^ n[5894];
assign t[5895] = t[5894] ^ n[5895];
assign t[5896] = t[5895] ^ n[5896];
assign t[5897] = t[5896] ^ n[5897];
assign t[5898] = t[5897] ^ n[5898];
assign t[5899] = t[5898] ^ n[5899];
assign t[5900] = t[5899] ^ n[5900];
assign t[5901] = t[5900] ^ n[5901];
assign t[5902] = t[5901] ^ n[5902];
assign t[5903] = t[5902] ^ n[5903];
assign t[5904] = t[5903] ^ n[5904];
assign t[5905] = t[5904] ^ n[5905];
assign t[5906] = t[5905] ^ n[5906];
assign t[5907] = t[5906] ^ n[5907];
assign t[5908] = t[5907] ^ n[5908];
assign t[5909] = t[5908] ^ n[5909];
assign t[5910] = t[5909] ^ n[5910];
assign t[5911] = t[5910] ^ n[5911];
assign t[5912] = t[5911] ^ n[5912];
assign t[5913] = t[5912] ^ n[5913];
assign t[5914] = t[5913] ^ n[5914];
assign t[5915] = t[5914] ^ n[5915];
assign t[5916] = t[5915] ^ n[5916];
assign t[5917] = t[5916] ^ n[5917];
assign t[5918] = t[5917] ^ n[5918];
assign t[5919] = t[5918] ^ n[5919];
assign t[5920] = t[5919] ^ n[5920];
assign t[5921] = t[5920] ^ n[5921];
assign t[5922] = t[5921] ^ n[5922];
assign t[5923] = t[5922] ^ n[5923];
assign t[5924] = t[5923] ^ n[5924];
assign t[5925] = t[5924] ^ n[5925];
assign t[5926] = t[5925] ^ n[5926];
assign t[5927] = t[5926] ^ n[5927];
assign t[5928] = t[5927] ^ n[5928];
assign t[5929] = t[5928] ^ n[5929];
assign t[5930] = t[5929] ^ n[5930];
assign t[5931] = t[5930] ^ n[5931];
assign t[5932] = t[5931] ^ n[5932];
assign t[5933] = t[5932] ^ n[5933];
assign t[5934] = t[5933] ^ n[5934];
assign t[5935] = t[5934] ^ n[5935];
assign t[5936] = t[5935] ^ n[5936];
assign t[5937] = t[5936] ^ n[5937];
assign t[5938] = t[5937] ^ n[5938];
assign t[5939] = t[5938] ^ n[5939];
assign t[5940] = t[5939] ^ n[5940];
assign t[5941] = t[5940] ^ n[5941];
assign t[5942] = t[5941] ^ n[5942];
assign t[5943] = t[5942] ^ n[5943];
assign t[5944] = t[5943] ^ n[5944];
assign t[5945] = t[5944] ^ n[5945];
assign t[5946] = t[5945] ^ n[5946];
assign t[5947] = t[5946] ^ n[5947];
assign t[5948] = t[5947] ^ n[5948];
assign t[5949] = t[5948] ^ n[5949];
assign t[5950] = t[5949] ^ n[5950];
assign t[5951] = t[5950] ^ n[5951];
assign t[5952] = t[5951] ^ n[5952];
assign t[5953] = t[5952] ^ n[5953];
assign t[5954] = t[5953] ^ n[5954];
assign t[5955] = t[5954] ^ n[5955];
assign t[5956] = t[5955] ^ n[5956];
assign t[5957] = t[5956] ^ n[5957];
assign t[5958] = t[5957] ^ n[5958];
assign t[5959] = t[5958] ^ n[5959];
assign t[5960] = t[5959] ^ n[5960];
assign t[5961] = t[5960] ^ n[5961];
assign t[5962] = t[5961] ^ n[5962];
assign t[5963] = t[5962] ^ n[5963];
assign t[5964] = t[5963] ^ n[5964];
assign t[5965] = t[5964] ^ n[5965];
assign t[5966] = t[5965] ^ n[5966];
assign t[5967] = t[5966] ^ n[5967];
assign t[5968] = t[5967] ^ n[5968];
assign t[5969] = t[5968] ^ n[5969];
assign t[5970] = t[5969] ^ n[5970];
assign t[5971] = t[5970] ^ n[5971];
assign t[5972] = t[5971] ^ n[5972];
assign t[5973] = t[5972] ^ n[5973];
assign t[5974] = t[5973] ^ n[5974];
assign t[5975] = t[5974] ^ n[5975];
assign t[5976] = t[5975] ^ n[5976];
assign t[5977] = t[5976] ^ n[5977];
assign t[5978] = t[5977] ^ n[5978];
assign t[5979] = t[5978] ^ n[5979];
assign t[5980] = t[5979] ^ n[5980];
assign t[5981] = t[5980] ^ n[5981];
assign t[5982] = t[5981] ^ n[5982];
assign t[5983] = t[5982] ^ n[5983];
assign t[5984] = t[5983] ^ n[5984];
assign t[5985] = t[5984] ^ n[5985];
assign t[5986] = t[5985] ^ n[5986];
assign t[5987] = t[5986] ^ n[5987];
assign t[5988] = t[5987] ^ n[5988];
assign t[5989] = t[5988] ^ n[5989];
assign t[5990] = t[5989] ^ n[5990];
assign t[5991] = t[5990] ^ n[5991];
assign t[5992] = t[5991] ^ n[5992];
assign t[5993] = t[5992] ^ n[5993];
assign t[5994] = t[5993] ^ n[5994];
assign t[5995] = t[5994] ^ n[5995];
assign t[5996] = t[5995] ^ n[5996];
assign t[5997] = t[5996] ^ n[5997];
assign t[5998] = t[5997] ^ n[5998];
assign t[5999] = t[5998] ^ n[5999];
assign t[6000] = t[5999] ^ n[6000];
assign t[6001] = t[6000] ^ n[6001];
assign t[6002] = t[6001] ^ n[6002];
assign t[6003] = t[6002] ^ n[6003];
assign t[6004] = t[6003] ^ n[6004];
assign t[6005] = t[6004] ^ n[6005];
assign t[6006] = t[6005] ^ n[6006];
assign t[6007] = t[6006] ^ n[6007];
assign t[6008] = t[6007] ^ n[6008];
assign t[6009] = t[6008] ^ n[6009];
assign t[6010] = t[6009] ^ n[6010];
assign t[6011] = t[6010] ^ n[6011];
assign t[6012] = t[6011] ^ n[6012];
assign t[6013] = t[6012] ^ n[6013];
assign t[6014] = t[6013] ^ n[6014];
assign t[6015] = t[6014] ^ n[6015];
assign t[6016] = t[6015] ^ n[6016];
assign t[6017] = t[6016] ^ n[6017];
assign t[6018] = t[6017] ^ n[6018];
assign t[6019] = t[6018] ^ n[6019];
assign t[6020] = t[6019] ^ n[6020];
assign t[6021] = t[6020] ^ n[6021];
assign t[6022] = t[6021] ^ n[6022];
assign t[6023] = t[6022] ^ n[6023];
assign t[6024] = t[6023] ^ n[6024];
assign t[6025] = t[6024] ^ n[6025];
assign t[6026] = t[6025] ^ n[6026];
assign t[6027] = t[6026] ^ n[6027];
assign t[6028] = t[6027] ^ n[6028];
assign t[6029] = t[6028] ^ n[6029];
assign t[6030] = t[6029] ^ n[6030];
assign t[6031] = t[6030] ^ n[6031];
assign t[6032] = t[6031] ^ n[6032];
assign t[6033] = t[6032] ^ n[6033];
assign t[6034] = t[6033] ^ n[6034];
assign t[6035] = t[6034] ^ n[6035];
assign t[6036] = t[6035] ^ n[6036];
assign t[6037] = t[6036] ^ n[6037];
assign t[6038] = t[6037] ^ n[6038];
assign t[6039] = t[6038] ^ n[6039];
assign t[6040] = t[6039] ^ n[6040];
assign t[6041] = t[6040] ^ n[6041];
assign t[6042] = t[6041] ^ n[6042];
assign t[6043] = t[6042] ^ n[6043];
assign t[6044] = t[6043] ^ n[6044];
assign t[6045] = t[6044] ^ n[6045];
assign t[6046] = t[6045] ^ n[6046];
assign t[6047] = t[6046] ^ n[6047];
assign t[6048] = t[6047] ^ n[6048];
assign t[6049] = t[6048] ^ n[6049];
assign t[6050] = t[6049] ^ n[6050];
assign t[6051] = t[6050] ^ n[6051];
assign t[6052] = t[6051] ^ n[6052];
assign t[6053] = t[6052] ^ n[6053];
assign t[6054] = t[6053] ^ n[6054];
assign t[6055] = t[6054] ^ n[6055];
assign t[6056] = t[6055] ^ n[6056];
assign t[6057] = t[6056] ^ n[6057];
assign t[6058] = t[6057] ^ n[6058];
assign t[6059] = t[6058] ^ n[6059];
assign t[6060] = t[6059] ^ n[6060];
assign t[6061] = t[6060] ^ n[6061];
assign t[6062] = t[6061] ^ n[6062];
assign t[6063] = t[6062] ^ n[6063];
assign t[6064] = t[6063] ^ n[6064];
assign t[6065] = t[6064] ^ n[6065];
assign t[6066] = t[6065] ^ n[6066];
assign t[6067] = t[6066] ^ n[6067];
assign t[6068] = t[6067] ^ n[6068];
assign t[6069] = t[6068] ^ n[6069];
assign t[6070] = t[6069] ^ n[6070];
assign t[6071] = t[6070] ^ n[6071];
assign t[6072] = t[6071] ^ n[6072];
assign t[6073] = t[6072] ^ n[6073];
assign t[6074] = t[6073] ^ n[6074];
assign t[6075] = t[6074] ^ n[6075];
assign t[6076] = t[6075] ^ n[6076];
assign t[6077] = t[6076] ^ n[6077];
assign t[6078] = t[6077] ^ n[6078];
assign t[6079] = t[6078] ^ n[6079];
assign t[6080] = t[6079] ^ n[6080];
assign t[6081] = t[6080] ^ n[6081];
assign t[6082] = t[6081] ^ n[6082];
assign t[6083] = t[6082] ^ n[6083];
assign t[6084] = t[6083] ^ n[6084];
assign t[6085] = t[6084] ^ n[6085];
assign t[6086] = t[6085] ^ n[6086];
assign t[6087] = t[6086] ^ n[6087];
assign t[6088] = t[6087] ^ n[6088];
assign t[6089] = t[6088] ^ n[6089];
assign t[6090] = t[6089] ^ n[6090];
assign t[6091] = t[6090] ^ n[6091];
assign t[6092] = t[6091] ^ n[6092];
assign t[6093] = t[6092] ^ n[6093];
assign t[6094] = t[6093] ^ n[6094];
assign t[6095] = t[6094] ^ n[6095];
assign t[6096] = t[6095] ^ n[6096];
assign t[6097] = t[6096] ^ n[6097];
assign t[6098] = t[6097] ^ n[6098];
assign t[6099] = t[6098] ^ n[6099];
assign t[6100] = t[6099] ^ n[6100];
assign t[6101] = t[6100] ^ n[6101];
assign t[6102] = t[6101] ^ n[6102];
assign t[6103] = t[6102] ^ n[6103];
assign t[6104] = t[6103] ^ n[6104];
assign t[6105] = t[6104] ^ n[6105];
assign t[6106] = t[6105] ^ n[6106];
assign t[6107] = t[6106] ^ n[6107];
assign t[6108] = t[6107] ^ n[6108];
assign t[6109] = t[6108] ^ n[6109];
assign t[6110] = t[6109] ^ n[6110];
assign t[6111] = t[6110] ^ n[6111];
assign t[6112] = t[6111] ^ n[6112];
assign t[6113] = t[6112] ^ n[6113];
assign t[6114] = t[6113] ^ n[6114];
assign t[6115] = t[6114] ^ n[6115];
assign t[6116] = t[6115] ^ n[6116];
assign t[6117] = t[6116] ^ n[6117];
assign t[6118] = t[6117] ^ n[6118];
assign t[6119] = t[6118] ^ n[6119];
assign t[6120] = t[6119] ^ n[6120];
assign t[6121] = t[6120] ^ n[6121];
assign t[6122] = t[6121] ^ n[6122];
assign t[6123] = t[6122] ^ n[6123];
assign t[6124] = t[6123] ^ n[6124];
assign t[6125] = t[6124] ^ n[6125];
assign t[6126] = t[6125] ^ n[6126];
assign t[6127] = t[6126] ^ n[6127];
assign t[6128] = t[6127] ^ n[6128];
assign t[6129] = t[6128] ^ n[6129];
assign t[6130] = t[6129] ^ n[6130];
assign t[6131] = t[6130] ^ n[6131];
assign t[6132] = t[6131] ^ n[6132];
assign t[6133] = t[6132] ^ n[6133];
assign t[6134] = t[6133] ^ n[6134];
assign t[6135] = t[6134] ^ n[6135];
assign t[6136] = t[6135] ^ n[6136];
assign t[6137] = t[6136] ^ n[6137];
assign t[6138] = t[6137] ^ n[6138];
assign t[6139] = t[6138] ^ n[6139];
assign t[6140] = t[6139] ^ n[6140];
assign t[6141] = t[6140] ^ n[6141];
assign t[6142] = t[6141] ^ n[6142];
assign t[6143] = t[6142] ^ n[6143];
assign t[6144] = t[6143] ^ n[6144];
assign t[6145] = t[6144] ^ n[6145];
assign t[6146] = t[6145] ^ n[6146];
assign t[6147] = t[6146] ^ n[6147];
assign t[6148] = t[6147] ^ n[6148];
assign t[6149] = t[6148] ^ n[6149];
assign t[6150] = t[6149] ^ n[6150];
assign t[6151] = t[6150] ^ n[6151];
assign t[6152] = t[6151] ^ n[6152];
assign t[6153] = t[6152] ^ n[6153];
assign t[6154] = t[6153] ^ n[6154];
assign t[6155] = t[6154] ^ n[6155];
assign t[6156] = t[6155] ^ n[6156];
assign t[6157] = t[6156] ^ n[6157];
assign t[6158] = t[6157] ^ n[6158];
assign t[6159] = t[6158] ^ n[6159];
assign t[6160] = t[6159] ^ n[6160];
assign t[6161] = t[6160] ^ n[6161];
assign t[6162] = t[6161] ^ n[6162];
assign t[6163] = t[6162] ^ n[6163];
assign t[6164] = t[6163] ^ n[6164];
assign t[6165] = t[6164] ^ n[6165];
assign t[6166] = t[6165] ^ n[6166];
assign t[6167] = t[6166] ^ n[6167];
assign t[6168] = t[6167] ^ n[6168];
assign t[6169] = t[6168] ^ n[6169];
assign t[6170] = t[6169] ^ n[6170];
assign t[6171] = t[6170] ^ n[6171];
assign t[6172] = t[6171] ^ n[6172];
assign t[6173] = t[6172] ^ n[6173];
assign t[6174] = t[6173] ^ n[6174];
assign t[6175] = t[6174] ^ n[6175];
assign t[6176] = t[6175] ^ n[6176];
assign t[6177] = t[6176] ^ n[6177];
assign t[6178] = t[6177] ^ n[6178];
assign t[6179] = t[6178] ^ n[6179];
assign t[6180] = t[6179] ^ n[6180];
assign t[6181] = t[6180] ^ n[6181];
assign t[6182] = t[6181] ^ n[6182];
assign t[6183] = t[6182] ^ n[6183];
assign t[6184] = t[6183] ^ n[6184];
assign t[6185] = t[6184] ^ n[6185];
assign t[6186] = t[6185] ^ n[6186];
assign t[6187] = t[6186] ^ n[6187];
assign t[6188] = t[6187] ^ n[6188];
assign t[6189] = t[6188] ^ n[6189];
assign t[6190] = t[6189] ^ n[6190];
assign t[6191] = t[6190] ^ n[6191];
assign t[6192] = t[6191] ^ n[6192];
assign t[6193] = t[6192] ^ n[6193];
assign t[6194] = t[6193] ^ n[6194];
assign t[6195] = t[6194] ^ n[6195];
assign t[6196] = t[6195] ^ n[6196];
assign t[6197] = t[6196] ^ n[6197];
assign t[6198] = t[6197] ^ n[6198];
assign t[6199] = t[6198] ^ n[6199];
assign t[6200] = t[6199] ^ n[6200];
assign t[6201] = t[6200] ^ n[6201];
assign t[6202] = t[6201] ^ n[6202];
assign t[6203] = t[6202] ^ n[6203];
assign t[6204] = t[6203] ^ n[6204];
assign t[6205] = t[6204] ^ n[6205];
assign t[6206] = t[6205] ^ n[6206];
assign t[6207] = t[6206] ^ n[6207];
assign t[6208] = t[6207] ^ n[6208];
assign t[6209] = t[6208] ^ n[6209];
assign t[6210] = t[6209] ^ n[6210];
assign t[6211] = t[6210] ^ n[6211];
assign t[6212] = t[6211] ^ n[6212];
assign t[6213] = t[6212] ^ n[6213];
assign t[6214] = t[6213] ^ n[6214];
assign t[6215] = t[6214] ^ n[6215];
assign t[6216] = t[6215] ^ n[6216];
assign t[6217] = t[6216] ^ n[6217];
assign t[6218] = t[6217] ^ n[6218];
assign t[6219] = t[6218] ^ n[6219];
assign t[6220] = t[6219] ^ n[6220];
assign t[6221] = t[6220] ^ n[6221];
assign t[6222] = t[6221] ^ n[6222];
assign t[6223] = t[6222] ^ n[6223];
assign t[6224] = t[6223] ^ n[6224];
assign t[6225] = t[6224] ^ n[6225];
assign t[6226] = t[6225] ^ n[6226];
assign t[6227] = t[6226] ^ n[6227];
assign t[6228] = t[6227] ^ n[6228];
assign t[6229] = t[6228] ^ n[6229];
assign t[6230] = t[6229] ^ n[6230];
assign t[6231] = t[6230] ^ n[6231];
assign t[6232] = t[6231] ^ n[6232];
assign t[6233] = t[6232] ^ n[6233];
assign t[6234] = t[6233] ^ n[6234];
assign t[6235] = t[6234] ^ n[6235];
assign t[6236] = t[6235] ^ n[6236];
assign t[6237] = t[6236] ^ n[6237];
assign t[6238] = t[6237] ^ n[6238];
assign t[6239] = t[6238] ^ n[6239];
assign t[6240] = t[6239] ^ n[6240];
assign t[6241] = t[6240] ^ n[6241];
assign t[6242] = t[6241] ^ n[6242];
assign t[6243] = t[6242] ^ n[6243];
assign t[6244] = t[6243] ^ n[6244];
assign t[6245] = t[6244] ^ n[6245];
assign t[6246] = t[6245] ^ n[6246];
assign t[6247] = t[6246] ^ n[6247];
assign t[6248] = t[6247] ^ n[6248];
assign t[6249] = t[6248] ^ n[6249];
assign t[6250] = t[6249] ^ n[6250];
assign t[6251] = t[6250] ^ n[6251];
assign t[6252] = t[6251] ^ n[6252];
assign t[6253] = t[6252] ^ n[6253];
assign t[6254] = t[6253] ^ n[6254];
assign t[6255] = t[6254] ^ n[6255];
assign t[6256] = t[6255] ^ n[6256];
assign t[6257] = t[6256] ^ n[6257];
assign t[6258] = t[6257] ^ n[6258];
assign t[6259] = t[6258] ^ n[6259];
assign t[6260] = t[6259] ^ n[6260];
assign t[6261] = t[6260] ^ n[6261];
assign t[6262] = t[6261] ^ n[6262];
assign t[6263] = t[6262] ^ n[6263];
assign t[6264] = t[6263] ^ n[6264];
assign t[6265] = t[6264] ^ n[6265];
assign t[6266] = t[6265] ^ n[6266];
assign t[6267] = t[6266] ^ n[6267];
assign t[6268] = t[6267] ^ n[6268];
assign t[6269] = t[6268] ^ n[6269];
assign t[6270] = t[6269] ^ n[6270];
assign t[6271] = t[6270] ^ n[6271];
assign t[6272] = t[6271] ^ n[6272];
assign t[6273] = t[6272] ^ n[6273];
assign t[6274] = t[6273] ^ n[6274];
assign t[6275] = t[6274] ^ n[6275];
assign t[6276] = t[6275] ^ n[6276];
assign t[6277] = t[6276] ^ n[6277];
assign t[6278] = t[6277] ^ n[6278];
assign t[6279] = t[6278] ^ n[6279];
assign t[6280] = t[6279] ^ n[6280];
assign t[6281] = t[6280] ^ n[6281];
assign t[6282] = t[6281] ^ n[6282];
assign t[6283] = t[6282] ^ n[6283];
assign t[6284] = t[6283] ^ n[6284];
assign t[6285] = t[6284] ^ n[6285];
assign t[6286] = t[6285] ^ n[6286];
assign t[6287] = t[6286] ^ n[6287];
assign t[6288] = t[6287] ^ n[6288];
assign t[6289] = t[6288] ^ n[6289];
assign t[6290] = t[6289] ^ n[6290];
assign t[6291] = t[6290] ^ n[6291];
assign t[6292] = t[6291] ^ n[6292];
assign t[6293] = t[6292] ^ n[6293];
assign t[6294] = t[6293] ^ n[6294];
assign t[6295] = t[6294] ^ n[6295];
assign t[6296] = t[6295] ^ n[6296];
assign t[6297] = t[6296] ^ n[6297];
assign t[6298] = t[6297] ^ n[6298];
assign t[6299] = t[6298] ^ n[6299];
assign t[6300] = t[6299] ^ n[6300];
assign t[6301] = t[6300] ^ n[6301];
assign t[6302] = t[6301] ^ n[6302];
assign t[6303] = t[6302] ^ n[6303];
assign t[6304] = t[6303] ^ n[6304];
assign t[6305] = t[6304] ^ n[6305];
assign t[6306] = t[6305] ^ n[6306];
assign t[6307] = t[6306] ^ n[6307];
assign t[6308] = t[6307] ^ n[6308];
assign t[6309] = t[6308] ^ n[6309];
assign t[6310] = t[6309] ^ n[6310];
assign t[6311] = t[6310] ^ n[6311];
assign t[6312] = t[6311] ^ n[6312];
assign t[6313] = t[6312] ^ n[6313];
assign t[6314] = t[6313] ^ n[6314];
assign t[6315] = t[6314] ^ n[6315];
assign t[6316] = t[6315] ^ n[6316];
assign t[6317] = t[6316] ^ n[6317];
assign t[6318] = t[6317] ^ n[6318];
assign t[6319] = t[6318] ^ n[6319];
assign t[6320] = t[6319] ^ n[6320];
assign t[6321] = t[6320] ^ n[6321];
assign t[6322] = t[6321] ^ n[6322];
assign t[6323] = t[6322] ^ n[6323];
assign t[6324] = t[6323] ^ n[6324];
assign t[6325] = t[6324] ^ n[6325];
assign t[6326] = t[6325] ^ n[6326];
assign t[6327] = t[6326] ^ n[6327];
assign t[6328] = t[6327] ^ n[6328];
assign t[6329] = t[6328] ^ n[6329];
assign t[6330] = t[6329] ^ n[6330];
assign t[6331] = t[6330] ^ n[6331];
assign t[6332] = t[6331] ^ n[6332];
assign t[6333] = t[6332] ^ n[6333];
assign t[6334] = t[6333] ^ n[6334];
assign t[6335] = t[6334] ^ n[6335];
assign t[6336] = t[6335] ^ n[6336];
assign t[6337] = t[6336] ^ n[6337];
assign t[6338] = t[6337] ^ n[6338];
assign t[6339] = t[6338] ^ n[6339];
assign t[6340] = t[6339] ^ n[6340];
assign t[6341] = t[6340] ^ n[6341];
assign t[6342] = t[6341] ^ n[6342];
assign t[6343] = t[6342] ^ n[6343];
assign t[6344] = t[6343] ^ n[6344];
assign t[6345] = t[6344] ^ n[6345];
assign t[6346] = t[6345] ^ n[6346];
assign t[6347] = t[6346] ^ n[6347];
assign t[6348] = t[6347] ^ n[6348];
assign t[6349] = t[6348] ^ n[6349];
assign t[6350] = t[6349] ^ n[6350];
assign t[6351] = t[6350] ^ n[6351];
assign t[6352] = t[6351] ^ n[6352];
assign t[6353] = t[6352] ^ n[6353];
assign t[6354] = t[6353] ^ n[6354];
assign t[6355] = t[6354] ^ n[6355];
assign t[6356] = t[6355] ^ n[6356];
assign t[6357] = t[6356] ^ n[6357];
assign t[6358] = t[6357] ^ n[6358];
assign t[6359] = t[6358] ^ n[6359];
assign t[6360] = t[6359] ^ n[6360];
assign t[6361] = t[6360] ^ n[6361];
assign t[6362] = t[6361] ^ n[6362];
assign t[6363] = t[6362] ^ n[6363];
assign t[6364] = t[6363] ^ n[6364];
assign t[6365] = t[6364] ^ n[6365];
assign t[6366] = t[6365] ^ n[6366];
assign t[6367] = t[6366] ^ n[6367];
assign t[6368] = t[6367] ^ n[6368];
assign t[6369] = t[6368] ^ n[6369];
assign t[6370] = t[6369] ^ n[6370];
assign t[6371] = t[6370] ^ n[6371];
assign t[6372] = t[6371] ^ n[6372];
assign t[6373] = t[6372] ^ n[6373];
assign t[6374] = t[6373] ^ n[6374];
assign t[6375] = t[6374] ^ n[6375];
assign t[6376] = t[6375] ^ n[6376];
assign t[6377] = t[6376] ^ n[6377];
assign t[6378] = t[6377] ^ n[6378];
assign t[6379] = t[6378] ^ n[6379];
assign t[6380] = t[6379] ^ n[6380];
assign t[6381] = t[6380] ^ n[6381];
assign t[6382] = t[6381] ^ n[6382];
assign t[6383] = t[6382] ^ n[6383];
assign t[6384] = t[6383] ^ n[6384];
assign t[6385] = t[6384] ^ n[6385];
assign t[6386] = t[6385] ^ n[6386];
assign t[6387] = t[6386] ^ n[6387];
assign t[6388] = t[6387] ^ n[6388];
assign t[6389] = t[6388] ^ n[6389];
assign t[6390] = t[6389] ^ n[6390];
assign t[6391] = t[6390] ^ n[6391];
assign t[6392] = t[6391] ^ n[6392];
assign t[6393] = t[6392] ^ n[6393];
assign t[6394] = t[6393] ^ n[6394];
assign t[6395] = t[6394] ^ n[6395];
assign t[6396] = t[6395] ^ n[6396];
assign t[6397] = t[6396] ^ n[6397];
assign t[6398] = t[6397] ^ n[6398];
assign t[6399] = t[6398] ^ n[6399];
assign t[6400] = t[6399] ^ n[6400];
assign t[6401] = t[6400] ^ n[6401];
assign t[6402] = t[6401] ^ n[6402];
assign t[6403] = t[6402] ^ n[6403];
assign t[6404] = t[6403] ^ n[6404];
assign t[6405] = t[6404] ^ n[6405];
assign t[6406] = t[6405] ^ n[6406];
assign t[6407] = t[6406] ^ n[6407];
assign t[6408] = t[6407] ^ n[6408];
assign t[6409] = t[6408] ^ n[6409];
assign t[6410] = t[6409] ^ n[6410];
assign t[6411] = t[6410] ^ n[6411];
assign t[6412] = t[6411] ^ n[6412];
assign t[6413] = t[6412] ^ n[6413];
assign t[6414] = t[6413] ^ n[6414];
assign t[6415] = t[6414] ^ n[6415];
assign t[6416] = t[6415] ^ n[6416];
assign t[6417] = t[6416] ^ n[6417];
assign t[6418] = t[6417] ^ n[6418];
assign t[6419] = t[6418] ^ n[6419];
assign t[6420] = t[6419] ^ n[6420];
assign t[6421] = t[6420] ^ n[6421];
assign t[6422] = t[6421] ^ n[6422];
assign t[6423] = t[6422] ^ n[6423];
assign t[6424] = t[6423] ^ n[6424];
assign t[6425] = t[6424] ^ n[6425];
assign t[6426] = t[6425] ^ n[6426];
assign t[6427] = t[6426] ^ n[6427];
assign t[6428] = t[6427] ^ n[6428];
assign t[6429] = t[6428] ^ n[6429];
assign t[6430] = t[6429] ^ n[6430];
assign t[6431] = t[6430] ^ n[6431];
assign t[6432] = t[6431] ^ n[6432];
assign t[6433] = t[6432] ^ n[6433];
assign t[6434] = t[6433] ^ n[6434];
assign t[6435] = t[6434] ^ n[6435];
assign t[6436] = t[6435] ^ n[6436];
assign t[6437] = t[6436] ^ n[6437];
assign t[6438] = t[6437] ^ n[6438];
assign t[6439] = t[6438] ^ n[6439];
assign t[6440] = t[6439] ^ n[6440];
assign t[6441] = t[6440] ^ n[6441];
assign t[6442] = t[6441] ^ n[6442];
assign t[6443] = t[6442] ^ n[6443];
assign t[6444] = t[6443] ^ n[6444];
assign t[6445] = t[6444] ^ n[6445];
assign t[6446] = t[6445] ^ n[6446];
assign t[6447] = t[6446] ^ n[6447];
assign t[6448] = t[6447] ^ n[6448];
assign t[6449] = t[6448] ^ n[6449];
assign t[6450] = t[6449] ^ n[6450];
assign t[6451] = t[6450] ^ n[6451];
assign t[6452] = t[6451] ^ n[6452];
assign t[6453] = t[6452] ^ n[6453];
assign t[6454] = t[6453] ^ n[6454];
assign t[6455] = t[6454] ^ n[6455];
assign t[6456] = t[6455] ^ n[6456];
assign t[6457] = t[6456] ^ n[6457];
assign t[6458] = t[6457] ^ n[6458];
assign t[6459] = t[6458] ^ n[6459];
assign t[6460] = t[6459] ^ n[6460];
assign t[6461] = t[6460] ^ n[6461];
assign t[6462] = t[6461] ^ n[6462];
assign t[6463] = t[6462] ^ n[6463];
assign t[6464] = t[6463] ^ n[6464];
assign t[6465] = t[6464] ^ n[6465];
assign t[6466] = t[6465] ^ n[6466];
assign t[6467] = t[6466] ^ n[6467];
assign t[6468] = t[6467] ^ n[6468];
assign t[6469] = t[6468] ^ n[6469];
assign t[6470] = t[6469] ^ n[6470];
assign t[6471] = t[6470] ^ n[6471];
assign t[6472] = t[6471] ^ n[6472];
assign t[6473] = t[6472] ^ n[6473];
assign t[6474] = t[6473] ^ n[6474];
assign t[6475] = t[6474] ^ n[6475];
assign t[6476] = t[6475] ^ n[6476];
assign t[6477] = t[6476] ^ n[6477];
assign t[6478] = t[6477] ^ n[6478];
assign t[6479] = t[6478] ^ n[6479];
assign t[6480] = t[6479] ^ n[6480];
assign t[6481] = t[6480] ^ n[6481];
assign t[6482] = t[6481] ^ n[6482];
assign t[6483] = t[6482] ^ n[6483];
assign t[6484] = t[6483] ^ n[6484];
assign t[6485] = t[6484] ^ n[6485];
assign t[6486] = t[6485] ^ n[6486];
assign t[6487] = t[6486] ^ n[6487];
assign t[6488] = t[6487] ^ n[6488];
assign t[6489] = t[6488] ^ n[6489];
assign t[6490] = t[6489] ^ n[6490];
assign t[6491] = t[6490] ^ n[6491];
assign t[6492] = t[6491] ^ n[6492];
assign t[6493] = t[6492] ^ n[6493];
assign t[6494] = t[6493] ^ n[6494];
assign t[6495] = t[6494] ^ n[6495];
assign t[6496] = t[6495] ^ n[6496];
assign t[6497] = t[6496] ^ n[6497];
assign t[6498] = t[6497] ^ n[6498];
assign t[6499] = t[6498] ^ n[6499];
assign t[6500] = t[6499] ^ n[6500];
assign t[6501] = t[6500] ^ n[6501];
assign t[6502] = t[6501] ^ n[6502];
assign t[6503] = t[6502] ^ n[6503];
assign t[6504] = t[6503] ^ n[6504];
assign t[6505] = t[6504] ^ n[6505];
assign t[6506] = t[6505] ^ n[6506];
assign t[6507] = t[6506] ^ n[6507];
assign t[6508] = t[6507] ^ n[6508];
assign t[6509] = t[6508] ^ n[6509];
assign t[6510] = t[6509] ^ n[6510];
assign t[6511] = t[6510] ^ n[6511];
assign t[6512] = t[6511] ^ n[6512];
assign t[6513] = t[6512] ^ n[6513];
assign t[6514] = t[6513] ^ n[6514];
assign t[6515] = t[6514] ^ n[6515];
assign t[6516] = t[6515] ^ n[6516];
assign t[6517] = t[6516] ^ n[6517];
assign t[6518] = t[6517] ^ n[6518];
assign t[6519] = t[6518] ^ n[6519];
assign t[6520] = t[6519] ^ n[6520];
assign t[6521] = t[6520] ^ n[6521];
assign t[6522] = t[6521] ^ n[6522];
assign t[6523] = t[6522] ^ n[6523];
assign t[6524] = t[6523] ^ n[6524];
assign t[6525] = t[6524] ^ n[6525];
assign t[6526] = t[6525] ^ n[6526];
assign t[6527] = t[6526] ^ n[6527];
assign t[6528] = t[6527] ^ n[6528];
assign t[6529] = t[6528] ^ n[6529];
assign t[6530] = t[6529] ^ n[6530];
assign t[6531] = t[6530] ^ n[6531];
assign t[6532] = t[6531] ^ n[6532];
assign t[6533] = t[6532] ^ n[6533];
assign t[6534] = t[6533] ^ n[6534];
assign t[6535] = t[6534] ^ n[6535];
assign t[6536] = t[6535] ^ n[6536];
assign t[6537] = t[6536] ^ n[6537];
assign t[6538] = t[6537] ^ n[6538];
assign t[6539] = t[6538] ^ n[6539];
assign t[6540] = t[6539] ^ n[6540];
assign t[6541] = t[6540] ^ n[6541];
assign t[6542] = t[6541] ^ n[6542];
assign t[6543] = t[6542] ^ n[6543];
assign t[6544] = t[6543] ^ n[6544];
assign t[6545] = t[6544] ^ n[6545];
assign t[6546] = t[6545] ^ n[6546];
assign t[6547] = t[6546] ^ n[6547];
assign t[6548] = t[6547] ^ n[6548];
assign t[6549] = t[6548] ^ n[6549];
assign t[6550] = t[6549] ^ n[6550];
assign t[6551] = t[6550] ^ n[6551];
assign t[6552] = t[6551] ^ n[6552];
assign t[6553] = t[6552] ^ n[6553];
assign t[6554] = t[6553] ^ n[6554];
assign t[6555] = t[6554] ^ n[6555];
assign t[6556] = t[6555] ^ n[6556];
assign t[6557] = t[6556] ^ n[6557];
assign t[6558] = t[6557] ^ n[6558];
assign t[6559] = t[6558] ^ n[6559];
assign t[6560] = t[6559] ^ n[6560];
assign t[6561] = t[6560] ^ n[6561];
assign t[6562] = t[6561] ^ n[6562];
assign t[6563] = t[6562] ^ n[6563];
assign t[6564] = t[6563] ^ n[6564];
assign t[6565] = t[6564] ^ n[6565];
assign t[6566] = t[6565] ^ n[6566];
assign t[6567] = t[6566] ^ n[6567];
assign t[6568] = t[6567] ^ n[6568];
assign t[6569] = t[6568] ^ n[6569];
assign t[6570] = t[6569] ^ n[6570];
assign t[6571] = t[6570] ^ n[6571];
assign t[6572] = t[6571] ^ n[6572];
assign t[6573] = t[6572] ^ n[6573];
assign t[6574] = t[6573] ^ n[6574];
assign t[6575] = t[6574] ^ n[6575];
assign t[6576] = t[6575] ^ n[6576];
assign t[6577] = t[6576] ^ n[6577];
assign t[6578] = t[6577] ^ n[6578];
assign t[6579] = t[6578] ^ n[6579];
assign t[6580] = t[6579] ^ n[6580];
assign t[6581] = t[6580] ^ n[6581];
assign t[6582] = t[6581] ^ n[6582];
assign t[6583] = t[6582] ^ n[6583];
assign t[6584] = t[6583] ^ n[6584];
assign t[6585] = t[6584] ^ n[6585];
assign t[6586] = t[6585] ^ n[6586];
assign t[6587] = t[6586] ^ n[6587];
assign t[6588] = t[6587] ^ n[6588];
assign t[6589] = t[6588] ^ n[6589];
assign t[6590] = t[6589] ^ n[6590];
assign t[6591] = t[6590] ^ n[6591];
assign t[6592] = t[6591] ^ n[6592];
assign t[6593] = t[6592] ^ n[6593];
assign t[6594] = t[6593] ^ n[6594];
assign t[6595] = t[6594] ^ n[6595];
assign t[6596] = t[6595] ^ n[6596];
assign t[6597] = t[6596] ^ n[6597];
assign t[6598] = t[6597] ^ n[6598];
assign t[6599] = t[6598] ^ n[6599];
assign t[6600] = t[6599] ^ n[6600];
assign t[6601] = t[6600] ^ n[6601];
assign t[6602] = t[6601] ^ n[6602];
assign t[6603] = t[6602] ^ n[6603];
assign t[6604] = t[6603] ^ n[6604];
assign t[6605] = t[6604] ^ n[6605];
assign t[6606] = t[6605] ^ n[6606];
assign t[6607] = t[6606] ^ n[6607];
assign t[6608] = t[6607] ^ n[6608];
assign t[6609] = t[6608] ^ n[6609];
assign t[6610] = t[6609] ^ n[6610];
assign t[6611] = t[6610] ^ n[6611];
assign t[6612] = t[6611] ^ n[6612];
assign t[6613] = t[6612] ^ n[6613];
assign t[6614] = t[6613] ^ n[6614];
assign t[6615] = t[6614] ^ n[6615];
assign t[6616] = t[6615] ^ n[6616];
assign t[6617] = t[6616] ^ n[6617];
assign t[6618] = t[6617] ^ n[6618];
assign t[6619] = t[6618] ^ n[6619];
assign t[6620] = t[6619] ^ n[6620];
assign t[6621] = t[6620] ^ n[6621];
assign t[6622] = t[6621] ^ n[6622];
assign t[6623] = t[6622] ^ n[6623];
assign t[6624] = t[6623] ^ n[6624];
assign t[6625] = t[6624] ^ n[6625];
assign t[6626] = t[6625] ^ n[6626];
assign t[6627] = t[6626] ^ n[6627];
assign t[6628] = t[6627] ^ n[6628];
assign t[6629] = t[6628] ^ n[6629];
assign t[6630] = t[6629] ^ n[6630];
assign t[6631] = t[6630] ^ n[6631];
assign t[6632] = t[6631] ^ n[6632];
assign t[6633] = t[6632] ^ n[6633];
assign t[6634] = t[6633] ^ n[6634];
assign t[6635] = t[6634] ^ n[6635];
assign t[6636] = t[6635] ^ n[6636];
assign t[6637] = t[6636] ^ n[6637];
assign t[6638] = t[6637] ^ n[6638];
assign t[6639] = t[6638] ^ n[6639];
assign t[6640] = t[6639] ^ n[6640];
assign t[6641] = t[6640] ^ n[6641];
assign t[6642] = t[6641] ^ n[6642];
assign t[6643] = t[6642] ^ n[6643];
assign t[6644] = t[6643] ^ n[6644];
assign t[6645] = t[6644] ^ n[6645];
assign t[6646] = t[6645] ^ n[6646];
assign t[6647] = t[6646] ^ n[6647];
assign t[6648] = t[6647] ^ n[6648];
assign t[6649] = t[6648] ^ n[6649];
assign t[6650] = t[6649] ^ n[6650];
assign t[6651] = t[6650] ^ n[6651];
assign t[6652] = t[6651] ^ n[6652];
assign t[6653] = t[6652] ^ n[6653];
assign t[6654] = t[6653] ^ n[6654];
assign t[6655] = t[6654] ^ n[6655];
assign t[6656] = t[6655] ^ n[6656];
assign t[6657] = t[6656] ^ n[6657];
assign t[6658] = t[6657] ^ n[6658];
assign t[6659] = t[6658] ^ n[6659];
assign t[6660] = t[6659] ^ n[6660];
assign t[6661] = t[6660] ^ n[6661];
assign t[6662] = t[6661] ^ n[6662];
assign t[6663] = t[6662] ^ n[6663];
assign t[6664] = t[6663] ^ n[6664];
assign t[6665] = t[6664] ^ n[6665];
assign t[6666] = t[6665] ^ n[6666];
assign t[6667] = t[6666] ^ n[6667];
assign t[6668] = t[6667] ^ n[6668];
assign t[6669] = t[6668] ^ n[6669];
assign t[6670] = t[6669] ^ n[6670];
assign t[6671] = t[6670] ^ n[6671];
assign t[6672] = t[6671] ^ n[6672];
assign t[6673] = t[6672] ^ n[6673];
assign t[6674] = t[6673] ^ n[6674];
assign t[6675] = t[6674] ^ n[6675];
assign t[6676] = t[6675] ^ n[6676];
assign t[6677] = t[6676] ^ n[6677];
assign t[6678] = t[6677] ^ n[6678];
assign t[6679] = t[6678] ^ n[6679];
assign t[6680] = t[6679] ^ n[6680];
assign t[6681] = t[6680] ^ n[6681];
assign t[6682] = t[6681] ^ n[6682];
assign t[6683] = t[6682] ^ n[6683];
assign t[6684] = t[6683] ^ n[6684];
assign t[6685] = t[6684] ^ n[6685];
assign t[6686] = t[6685] ^ n[6686];
assign t[6687] = t[6686] ^ n[6687];
assign t[6688] = t[6687] ^ n[6688];
assign t[6689] = t[6688] ^ n[6689];
assign t[6690] = t[6689] ^ n[6690];
assign t[6691] = t[6690] ^ n[6691];
assign t[6692] = t[6691] ^ n[6692];
assign t[6693] = t[6692] ^ n[6693];
assign t[6694] = t[6693] ^ n[6694];
assign t[6695] = t[6694] ^ n[6695];
assign t[6696] = t[6695] ^ n[6696];
assign t[6697] = t[6696] ^ n[6697];
assign t[6698] = t[6697] ^ n[6698];
assign t[6699] = t[6698] ^ n[6699];
assign t[6700] = t[6699] ^ n[6700];
assign t[6701] = t[6700] ^ n[6701];
assign t[6702] = t[6701] ^ n[6702];
assign t[6703] = t[6702] ^ n[6703];
assign t[6704] = t[6703] ^ n[6704];
assign t[6705] = t[6704] ^ n[6705];
assign t[6706] = t[6705] ^ n[6706];
assign t[6707] = t[6706] ^ n[6707];
assign t[6708] = t[6707] ^ n[6708];
assign t[6709] = t[6708] ^ n[6709];
assign t[6710] = t[6709] ^ n[6710];
assign t[6711] = t[6710] ^ n[6711];
assign t[6712] = t[6711] ^ n[6712];
assign t[6713] = t[6712] ^ n[6713];
assign t[6714] = t[6713] ^ n[6714];
assign t[6715] = t[6714] ^ n[6715];
assign t[6716] = t[6715] ^ n[6716];
assign t[6717] = t[6716] ^ n[6717];
assign t[6718] = t[6717] ^ n[6718];
assign t[6719] = t[6718] ^ n[6719];
assign t[6720] = t[6719] ^ n[6720];
assign t[6721] = t[6720] ^ n[6721];
assign t[6722] = t[6721] ^ n[6722];
assign t[6723] = t[6722] ^ n[6723];
assign t[6724] = t[6723] ^ n[6724];
assign t[6725] = t[6724] ^ n[6725];
assign t[6726] = t[6725] ^ n[6726];
assign t[6727] = t[6726] ^ n[6727];
assign t[6728] = t[6727] ^ n[6728];
assign t[6729] = t[6728] ^ n[6729];
assign t[6730] = t[6729] ^ n[6730];
assign t[6731] = t[6730] ^ n[6731];
assign t[6732] = t[6731] ^ n[6732];
assign t[6733] = t[6732] ^ n[6733];
assign t[6734] = t[6733] ^ n[6734];
assign t[6735] = t[6734] ^ n[6735];
assign t[6736] = t[6735] ^ n[6736];
assign t[6737] = t[6736] ^ n[6737];
assign t[6738] = t[6737] ^ n[6738];
assign t[6739] = t[6738] ^ n[6739];
assign t[6740] = t[6739] ^ n[6740];
assign t[6741] = t[6740] ^ n[6741];
assign t[6742] = t[6741] ^ n[6742];
assign t[6743] = t[6742] ^ n[6743];
assign t[6744] = t[6743] ^ n[6744];
assign t[6745] = t[6744] ^ n[6745];
assign t[6746] = t[6745] ^ n[6746];
assign t[6747] = t[6746] ^ n[6747];
assign t[6748] = t[6747] ^ n[6748];
assign t[6749] = t[6748] ^ n[6749];
assign t[6750] = t[6749] ^ n[6750];
assign t[6751] = t[6750] ^ n[6751];
assign t[6752] = t[6751] ^ n[6752];
assign t[6753] = t[6752] ^ n[6753];
assign t[6754] = t[6753] ^ n[6754];
assign t[6755] = t[6754] ^ n[6755];
assign t[6756] = t[6755] ^ n[6756];
assign t[6757] = t[6756] ^ n[6757];
assign t[6758] = t[6757] ^ n[6758];
assign t[6759] = t[6758] ^ n[6759];
assign t[6760] = t[6759] ^ n[6760];
assign t[6761] = t[6760] ^ n[6761];
assign t[6762] = t[6761] ^ n[6762];
assign t[6763] = t[6762] ^ n[6763];
assign t[6764] = t[6763] ^ n[6764];
assign t[6765] = t[6764] ^ n[6765];
assign t[6766] = t[6765] ^ n[6766];
assign t[6767] = t[6766] ^ n[6767];
assign t[6768] = t[6767] ^ n[6768];
assign t[6769] = t[6768] ^ n[6769];
assign t[6770] = t[6769] ^ n[6770];
assign t[6771] = t[6770] ^ n[6771];
assign t[6772] = t[6771] ^ n[6772];
assign t[6773] = t[6772] ^ n[6773];
assign t[6774] = t[6773] ^ n[6774];
assign t[6775] = t[6774] ^ n[6775];
assign t[6776] = t[6775] ^ n[6776];
assign t[6777] = t[6776] ^ n[6777];
assign t[6778] = t[6777] ^ n[6778];
assign t[6779] = t[6778] ^ n[6779];
assign t[6780] = t[6779] ^ n[6780];
assign t[6781] = t[6780] ^ n[6781];
assign t[6782] = t[6781] ^ n[6782];
assign t[6783] = t[6782] ^ n[6783];
assign t[6784] = t[6783] ^ n[6784];
assign t[6785] = t[6784] ^ n[6785];
assign t[6786] = t[6785] ^ n[6786];
assign t[6787] = t[6786] ^ n[6787];
assign t[6788] = t[6787] ^ n[6788];
assign t[6789] = t[6788] ^ n[6789];
assign t[6790] = t[6789] ^ n[6790];
assign t[6791] = t[6790] ^ n[6791];
assign t[6792] = t[6791] ^ n[6792];
assign t[6793] = t[6792] ^ n[6793];
assign t[6794] = t[6793] ^ n[6794];
assign t[6795] = t[6794] ^ n[6795];
assign t[6796] = t[6795] ^ n[6796];
assign t[6797] = t[6796] ^ n[6797];
assign t[6798] = t[6797] ^ n[6798];
assign t[6799] = t[6798] ^ n[6799];
assign t[6800] = t[6799] ^ n[6800];
assign t[6801] = t[6800] ^ n[6801];
assign t[6802] = t[6801] ^ n[6802];
assign t[6803] = t[6802] ^ n[6803];
assign t[6804] = t[6803] ^ n[6804];
assign t[6805] = t[6804] ^ n[6805];
assign t[6806] = t[6805] ^ n[6806];
assign t[6807] = t[6806] ^ n[6807];
assign t[6808] = t[6807] ^ n[6808];
assign t[6809] = t[6808] ^ n[6809];
assign t[6810] = t[6809] ^ n[6810];
assign t[6811] = t[6810] ^ n[6811];
assign t[6812] = t[6811] ^ n[6812];
assign t[6813] = t[6812] ^ n[6813];
assign t[6814] = t[6813] ^ n[6814];
assign t[6815] = t[6814] ^ n[6815];
assign t[6816] = t[6815] ^ n[6816];
assign t[6817] = t[6816] ^ n[6817];
assign t[6818] = t[6817] ^ n[6818];
assign t[6819] = t[6818] ^ n[6819];
assign t[6820] = t[6819] ^ n[6820];
assign t[6821] = t[6820] ^ n[6821];
assign t[6822] = t[6821] ^ n[6822];
assign t[6823] = t[6822] ^ n[6823];
assign t[6824] = t[6823] ^ n[6824];
assign t[6825] = t[6824] ^ n[6825];
assign t[6826] = t[6825] ^ n[6826];
assign t[6827] = t[6826] ^ n[6827];
assign t[6828] = t[6827] ^ n[6828];
assign t[6829] = t[6828] ^ n[6829];
assign t[6830] = t[6829] ^ n[6830];
assign t[6831] = t[6830] ^ n[6831];
assign t[6832] = t[6831] ^ n[6832];
assign t[6833] = t[6832] ^ n[6833];
assign t[6834] = t[6833] ^ n[6834];
assign t[6835] = t[6834] ^ n[6835];
assign t[6836] = t[6835] ^ n[6836];
assign t[6837] = t[6836] ^ n[6837];
assign t[6838] = t[6837] ^ n[6838];
assign t[6839] = t[6838] ^ n[6839];
assign t[6840] = t[6839] ^ n[6840];
assign t[6841] = t[6840] ^ n[6841];
assign t[6842] = t[6841] ^ n[6842];
assign t[6843] = t[6842] ^ n[6843];
assign t[6844] = t[6843] ^ n[6844];
assign t[6845] = t[6844] ^ n[6845];
assign t[6846] = t[6845] ^ n[6846];
assign t[6847] = t[6846] ^ n[6847];
assign t[6848] = t[6847] ^ n[6848];
assign t[6849] = t[6848] ^ n[6849];
assign t[6850] = t[6849] ^ n[6850];
assign t[6851] = t[6850] ^ n[6851];
assign t[6852] = t[6851] ^ n[6852];
assign t[6853] = t[6852] ^ n[6853];
assign t[6854] = t[6853] ^ n[6854];
assign t[6855] = t[6854] ^ n[6855];
assign t[6856] = t[6855] ^ n[6856];
assign t[6857] = t[6856] ^ n[6857];
assign t[6858] = t[6857] ^ n[6858];
assign t[6859] = t[6858] ^ n[6859];
assign t[6860] = t[6859] ^ n[6860];
assign t[6861] = t[6860] ^ n[6861];
assign t[6862] = t[6861] ^ n[6862];
assign t[6863] = t[6862] ^ n[6863];
assign t[6864] = t[6863] ^ n[6864];
assign t[6865] = t[6864] ^ n[6865];
assign t[6866] = t[6865] ^ n[6866];
assign t[6867] = t[6866] ^ n[6867];
assign t[6868] = t[6867] ^ n[6868];
assign t[6869] = t[6868] ^ n[6869];
assign t[6870] = t[6869] ^ n[6870];
assign t[6871] = t[6870] ^ n[6871];
assign t[6872] = t[6871] ^ n[6872];
assign t[6873] = t[6872] ^ n[6873];
assign t[6874] = t[6873] ^ n[6874];
assign t[6875] = t[6874] ^ n[6875];
assign t[6876] = t[6875] ^ n[6876];
assign t[6877] = t[6876] ^ n[6877];
assign t[6878] = t[6877] ^ n[6878];
assign t[6879] = t[6878] ^ n[6879];
assign t[6880] = t[6879] ^ n[6880];
assign t[6881] = t[6880] ^ n[6881];
assign t[6882] = t[6881] ^ n[6882];
assign t[6883] = t[6882] ^ n[6883];
assign t[6884] = t[6883] ^ n[6884];
assign t[6885] = t[6884] ^ n[6885];
assign t[6886] = t[6885] ^ n[6886];
assign t[6887] = t[6886] ^ n[6887];
assign t[6888] = t[6887] ^ n[6888];
assign t[6889] = t[6888] ^ n[6889];
assign t[6890] = t[6889] ^ n[6890];
assign t[6891] = t[6890] ^ n[6891];
assign t[6892] = t[6891] ^ n[6892];
assign t[6893] = t[6892] ^ n[6893];
assign t[6894] = t[6893] ^ n[6894];
assign t[6895] = t[6894] ^ n[6895];
assign t[6896] = t[6895] ^ n[6896];
assign t[6897] = t[6896] ^ n[6897];
assign t[6898] = t[6897] ^ n[6898];
assign t[6899] = t[6898] ^ n[6899];
assign t[6900] = t[6899] ^ n[6900];
assign t[6901] = t[6900] ^ n[6901];
assign t[6902] = t[6901] ^ n[6902];
assign t[6903] = t[6902] ^ n[6903];
assign t[6904] = t[6903] ^ n[6904];
assign t[6905] = t[6904] ^ n[6905];
assign t[6906] = t[6905] ^ n[6906];
assign t[6907] = t[6906] ^ n[6907];
assign t[6908] = t[6907] ^ n[6908];
assign t[6909] = t[6908] ^ n[6909];
assign t[6910] = t[6909] ^ n[6910];
assign t[6911] = t[6910] ^ n[6911];
assign t[6912] = t[6911] ^ n[6912];
assign t[6913] = t[6912] ^ n[6913];
assign t[6914] = t[6913] ^ n[6914];
assign t[6915] = t[6914] ^ n[6915];
assign t[6916] = t[6915] ^ n[6916];
assign t[6917] = t[6916] ^ n[6917];
assign t[6918] = t[6917] ^ n[6918];
assign t[6919] = t[6918] ^ n[6919];
assign t[6920] = t[6919] ^ n[6920];
assign t[6921] = t[6920] ^ n[6921];
assign t[6922] = t[6921] ^ n[6922];
assign t[6923] = t[6922] ^ n[6923];
assign t[6924] = t[6923] ^ n[6924];
assign t[6925] = t[6924] ^ n[6925];
assign t[6926] = t[6925] ^ n[6926];
assign t[6927] = t[6926] ^ n[6927];
assign t[6928] = t[6927] ^ n[6928];
assign t[6929] = t[6928] ^ n[6929];
assign t[6930] = t[6929] ^ n[6930];
assign t[6931] = t[6930] ^ n[6931];
assign t[6932] = t[6931] ^ n[6932];
assign t[6933] = t[6932] ^ n[6933];
assign t[6934] = t[6933] ^ n[6934];
assign t[6935] = t[6934] ^ n[6935];
assign t[6936] = t[6935] ^ n[6936];
assign t[6937] = t[6936] ^ n[6937];
assign t[6938] = t[6937] ^ n[6938];
assign t[6939] = t[6938] ^ n[6939];
assign t[6940] = t[6939] ^ n[6940];
assign t[6941] = t[6940] ^ n[6941];
assign t[6942] = t[6941] ^ n[6942];
assign t[6943] = t[6942] ^ n[6943];
assign t[6944] = t[6943] ^ n[6944];
assign t[6945] = t[6944] ^ n[6945];
assign t[6946] = t[6945] ^ n[6946];
assign t[6947] = t[6946] ^ n[6947];
assign t[6948] = t[6947] ^ n[6948];
assign t[6949] = t[6948] ^ n[6949];
assign t[6950] = t[6949] ^ n[6950];
assign t[6951] = t[6950] ^ n[6951];
assign t[6952] = t[6951] ^ n[6952];
assign t[6953] = t[6952] ^ n[6953];
assign t[6954] = t[6953] ^ n[6954];
assign t[6955] = t[6954] ^ n[6955];
assign t[6956] = t[6955] ^ n[6956];
assign t[6957] = t[6956] ^ n[6957];
assign t[6958] = t[6957] ^ n[6958];
assign t[6959] = t[6958] ^ n[6959];
assign t[6960] = t[6959] ^ n[6960];
assign t[6961] = t[6960] ^ n[6961];
assign t[6962] = t[6961] ^ n[6962];
assign t[6963] = t[6962] ^ n[6963];
assign t[6964] = t[6963] ^ n[6964];
assign t[6965] = t[6964] ^ n[6965];
assign t[6966] = t[6965] ^ n[6966];
assign t[6967] = t[6966] ^ n[6967];
assign t[6968] = t[6967] ^ n[6968];
assign t[6969] = t[6968] ^ n[6969];
assign t[6970] = t[6969] ^ n[6970];
assign t[6971] = t[6970] ^ n[6971];
assign t[6972] = t[6971] ^ n[6972];
assign t[6973] = t[6972] ^ n[6973];
assign t[6974] = t[6973] ^ n[6974];
assign t[6975] = t[6974] ^ n[6975];
assign t[6976] = t[6975] ^ n[6976];
assign t[6977] = t[6976] ^ n[6977];
assign t[6978] = t[6977] ^ n[6978];
assign t[6979] = t[6978] ^ n[6979];
assign t[6980] = t[6979] ^ n[6980];
assign t[6981] = t[6980] ^ n[6981];
assign t[6982] = t[6981] ^ n[6982];
assign t[6983] = t[6982] ^ n[6983];
assign t[6984] = t[6983] ^ n[6984];
assign t[6985] = t[6984] ^ n[6985];
assign t[6986] = t[6985] ^ n[6986];
assign t[6987] = t[6986] ^ n[6987];
assign t[6988] = t[6987] ^ n[6988];
assign t[6989] = t[6988] ^ n[6989];
assign t[6990] = t[6989] ^ n[6990];
assign t[6991] = t[6990] ^ n[6991];
assign t[6992] = t[6991] ^ n[6992];
assign t[6993] = t[6992] ^ n[6993];
assign t[6994] = t[6993] ^ n[6994];
assign t[6995] = t[6994] ^ n[6995];
assign t[6996] = t[6995] ^ n[6996];
assign t[6997] = t[6996] ^ n[6997];
assign t[6998] = t[6997] ^ n[6998];
assign t[6999] = t[6998] ^ n[6999];
assign t[7000] = t[6999] ^ n[7000];
assign t[7001] = t[7000] ^ n[7001];
assign t[7002] = t[7001] ^ n[7002];
assign t[7003] = t[7002] ^ n[7003];
assign t[7004] = t[7003] ^ n[7004];
assign t[7005] = t[7004] ^ n[7005];
assign t[7006] = t[7005] ^ n[7006];
assign t[7007] = t[7006] ^ n[7007];
assign t[7008] = t[7007] ^ n[7008];
assign t[7009] = t[7008] ^ n[7009];
assign t[7010] = t[7009] ^ n[7010];
assign t[7011] = t[7010] ^ n[7011];
assign t[7012] = t[7011] ^ n[7012];
assign t[7013] = t[7012] ^ n[7013];
assign t[7014] = t[7013] ^ n[7014];
assign t[7015] = t[7014] ^ n[7015];
assign t[7016] = t[7015] ^ n[7016];
assign t[7017] = t[7016] ^ n[7017];
assign t[7018] = t[7017] ^ n[7018];
assign t[7019] = t[7018] ^ n[7019];
assign t[7020] = t[7019] ^ n[7020];
assign t[7021] = t[7020] ^ n[7021];
assign t[7022] = t[7021] ^ n[7022];
assign t[7023] = t[7022] ^ n[7023];
assign t[7024] = t[7023] ^ n[7024];
assign t[7025] = t[7024] ^ n[7025];
assign t[7026] = t[7025] ^ n[7026];
assign t[7027] = t[7026] ^ n[7027];
assign t[7028] = t[7027] ^ n[7028];
assign t[7029] = t[7028] ^ n[7029];
assign t[7030] = t[7029] ^ n[7030];
assign t[7031] = t[7030] ^ n[7031];
assign t[7032] = t[7031] ^ n[7032];
assign t[7033] = t[7032] ^ n[7033];
assign t[7034] = t[7033] ^ n[7034];
assign t[7035] = t[7034] ^ n[7035];
assign t[7036] = t[7035] ^ n[7036];
assign t[7037] = t[7036] ^ n[7037];
assign t[7038] = t[7037] ^ n[7038];
assign t[7039] = t[7038] ^ n[7039];
assign t[7040] = t[7039] ^ n[7040];
assign t[7041] = t[7040] ^ n[7041];
assign t[7042] = t[7041] ^ n[7042];
assign t[7043] = t[7042] ^ n[7043];
assign t[7044] = t[7043] ^ n[7044];
assign t[7045] = t[7044] ^ n[7045];
assign t[7046] = t[7045] ^ n[7046];
assign t[7047] = t[7046] ^ n[7047];
assign t[7048] = t[7047] ^ n[7048];
assign t[7049] = t[7048] ^ n[7049];
assign t[7050] = t[7049] ^ n[7050];
assign t[7051] = t[7050] ^ n[7051];
assign t[7052] = t[7051] ^ n[7052];
assign t[7053] = t[7052] ^ n[7053];
assign t[7054] = t[7053] ^ n[7054];
assign t[7055] = t[7054] ^ n[7055];
assign t[7056] = t[7055] ^ n[7056];
assign t[7057] = t[7056] ^ n[7057];
assign t[7058] = t[7057] ^ n[7058];
assign t[7059] = t[7058] ^ n[7059];
assign t[7060] = t[7059] ^ n[7060];
assign t[7061] = t[7060] ^ n[7061];
assign t[7062] = t[7061] ^ n[7062];
assign t[7063] = t[7062] ^ n[7063];
assign t[7064] = t[7063] ^ n[7064];
assign t[7065] = t[7064] ^ n[7065];
assign t[7066] = t[7065] ^ n[7066];
assign t[7067] = t[7066] ^ n[7067];
assign t[7068] = t[7067] ^ n[7068];
assign t[7069] = t[7068] ^ n[7069];
assign t[7070] = t[7069] ^ n[7070];
assign t[7071] = t[7070] ^ n[7071];
assign t[7072] = t[7071] ^ n[7072];
assign t[7073] = t[7072] ^ n[7073];
assign t[7074] = t[7073] ^ n[7074];
assign t[7075] = t[7074] ^ n[7075];
assign t[7076] = t[7075] ^ n[7076];
assign t[7077] = t[7076] ^ n[7077];
assign t[7078] = t[7077] ^ n[7078];
assign t[7079] = t[7078] ^ n[7079];
assign t[7080] = t[7079] ^ n[7080];
assign t[7081] = t[7080] ^ n[7081];
assign t[7082] = t[7081] ^ n[7082];
assign t[7083] = t[7082] ^ n[7083];
assign t[7084] = t[7083] ^ n[7084];
assign t[7085] = t[7084] ^ n[7085];
assign t[7086] = t[7085] ^ n[7086];
assign t[7087] = t[7086] ^ n[7087];
assign t[7088] = t[7087] ^ n[7088];
assign t[7089] = t[7088] ^ n[7089];
assign t[7090] = t[7089] ^ n[7090];
assign t[7091] = t[7090] ^ n[7091];
assign t[7092] = t[7091] ^ n[7092];
assign t[7093] = t[7092] ^ n[7093];
assign t[7094] = t[7093] ^ n[7094];
assign t[7095] = t[7094] ^ n[7095];
assign t[7096] = t[7095] ^ n[7096];
assign t[7097] = t[7096] ^ n[7097];
assign t[7098] = t[7097] ^ n[7098];
assign t[7099] = t[7098] ^ n[7099];
assign t[7100] = t[7099] ^ n[7100];
assign t[7101] = t[7100] ^ n[7101];
assign t[7102] = t[7101] ^ n[7102];
assign t[7103] = t[7102] ^ n[7103];
assign t[7104] = t[7103] ^ n[7104];
assign t[7105] = t[7104] ^ n[7105];
assign t[7106] = t[7105] ^ n[7106];
assign t[7107] = t[7106] ^ n[7107];
assign t[7108] = t[7107] ^ n[7108];
assign t[7109] = t[7108] ^ n[7109];
assign t[7110] = t[7109] ^ n[7110];
assign t[7111] = t[7110] ^ n[7111];
assign t[7112] = t[7111] ^ n[7112];
assign t[7113] = t[7112] ^ n[7113];
assign t[7114] = t[7113] ^ n[7114];
assign t[7115] = t[7114] ^ n[7115];
assign t[7116] = t[7115] ^ n[7116];
assign t[7117] = t[7116] ^ n[7117];
assign t[7118] = t[7117] ^ n[7118];
assign t[7119] = t[7118] ^ n[7119];
assign t[7120] = t[7119] ^ n[7120];
assign t[7121] = t[7120] ^ n[7121];
assign t[7122] = t[7121] ^ n[7122];
assign t[7123] = t[7122] ^ n[7123];
assign t[7124] = t[7123] ^ n[7124];
assign t[7125] = t[7124] ^ n[7125];
assign t[7126] = t[7125] ^ n[7126];
assign t[7127] = t[7126] ^ n[7127];
assign t[7128] = t[7127] ^ n[7128];
assign t[7129] = t[7128] ^ n[7129];
assign t[7130] = t[7129] ^ n[7130];
assign t[7131] = t[7130] ^ n[7131];
assign t[7132] = t[7131] ^ n[7132];
assign t[7133] = t[7132] ^ n[7133];
assign t[7134] = t[7133] ^ n[7134];
assign t[7135] = t[7134] ^ n[7135];
assign t[7136] = t[7135] ^ n[7136];
assign t[7137] = t[7136] ^ n[7137];
assign t[7138] = t[7137] ^ n[7138];
assign t[7139] = t[7138] ^ n[7139];
assign t[7140] = t[7139] ^ n[7140];
assign t[7141] = t[7140] ^ n[7141];
assign t[7142] = t[7141] ^ n[7142];
assign t[7143] = t[7142] ^ n[7143];
assign t[7144] = t[7143] ^ n[7144];
assign t[7145] = t[7144] ^ n[7145];
assign t[7146] = t[7145] ^ n[7146];
assign t[7147] = t[7146] ^ n[7147];
assign t[7148] = t[7147] ^ n[7148];
assign t[7149] = t[7148] ^ n[7149];
assign t[7150] = t[7149] ^ n[7150];
assign t[7151] = t[7150] ^ n[7151];
assign t[7152] = t[7151] ^ n[7152];
assign t[7153] = t[7152] ^ n[7153];
assign t[7154] = t[7153] ^ n[7154];
assign t[7155] = t[7154] ^ n[7155];
assign t[7156] = t[7155] ^ n[7156];
assign t[7157] = t[7156] ^ n[7157];
assign t[7158] = t[7157] ^ n[7158];
assign t[7159] = t[7158] ^ n[7159];
assign t[7160] = t[7159] ^ n[7160];
assign t[7161] = t[7160] ^ n[7161];
assign t[7162] = t[7161] ^ n[7162];
assign t[7163] = t[7162] ^ n[7163];
assign t[7164] = t[7163] ^ n[7164];
assign t[7165] = t[7164] ^ n[7165];
assign t[7166] = t[7165] ^ n[7166];
assign t[7167] = t[7166] ^ n[7167];
assign t[7168] = t[7167] ^ n[7168];
assign t[7169] = t[7168] ^ n[7169];
assign t[7170] = t[7169] ^ n[7170];
assign t[7171] = t[7170] ^ n[7171];
assign t[7172] = t[7171] ^ n[7172];
assign t[7173] = t[7172] ^ n[7173];
assign t[7174] = t[7173] ^ n[7174];
assign t[7175] = t[7174] ^ n[7175];
assign t[7176] = t[7175] ^ n[7176];
assign t[7177] = t[7176] ^ n[7177];
assign t[7178] = t[7177] ^ n[7178];
assign t[7179] = t[7178] ^ n[7179];
assign t[7180] = t[7179] ^ n[7180];
assign t[7181] = t[7180] ^ n[7181];
assign t[7182] = t[7181] ^ n[7182];
assign t[7183] = t[7182] ^ n[7183];
assign t[7184] = t[7183] ^ n[7184];
assign t[7185] = t[7184] ^ n[7185];
assign t[7186] = t[7185] ^ n[7186];
assign t[7187] = t[7186] ^ n[7187];
assign t[7188] = t[7187] ^ n[7188];
assign t[7189] = t[7188] ^ n[7189];
assign t[7190] = t[7189] ^ n[7190];
assign t[7191] = t[7190] ^ n[7191];
assign t[7192] = t[7191] ^ n[7192];
assign t[7193] = t[7192] ^ n[7193];
assign t[7194] = t[7193] ^ n[7194];
assign t[7195] = t[7194] ^ n[7195];
assign t[7196] = t[7195] ^ n[7196];
assign t[7197] = t[7196] ^ n[7197];
assign t[7198] = t[7197] ^ n[7198];
assign t[7199] = t[7198] ^ n[7199];
assign t[7200] = t[7199] ^ n[7200];
assign t[7201] = t[7200] ^ n[7201];
assign t[7202] = t[7201] ^ n[7202];
assign t[7203] = t[7202] ^ n[7203];
assign t[7204] = t[7203] ^ n[7204];
assign t[7205] = t[7204] ^ n[7205];
assign t[7206] = t[7205] ^ n[7206];
assign t[7207] = t[7206] ^ n[7207];
assign t[7208] = t[7207] ^ n[7208];
assign t[7209] = t[7208] ^ n[7209];
assign t[7210] = t[7209] ^ n[7210];
assign t[7211] = t[7210] ^ n[7211];
assign t[7212] = t[7211] ^ n[7212];
assign t[7213] = t[7212] ^ n[7213];
assign t[7214] = t[7213] ^ n[7214];
assign t[7215] = t[7214] ^ n[7215];
assign t[7216] = t[7215] ^ n[7216];
assign t[7217] = t[7216] ^ n[7217];
assign t[7218] = t[7217] ^ n[7218];
assign t[7219] = t[7218] ^ n[7219];
assign t[7220] = t[7219] ^ n[7220];
assign t[7221] = t[7220] ^ n[7221];
assign t[7222] = t[7221] ^ n[7222];
assign t[7223] = t[7222] ^ n[7223];
assign t[7224] = t[7223] ^ n[7224];
assign t[7225] = t[7224] ^ n[7225];
assign t[7226] = t[7225] ^ n[7226];
assign t[7227] = t[7226] ^ n[7227];
assign t[7228] = t[7227] ^ n[7228];
assign t[7229] = t[7228] ^ n[7229];
assign t[7230] = t[7229] ^ n[7230];
assign t[7231] = t[7230] ^ n[7231];
assign t[7232] = t[7231] ^ n[7232];
assign t[7233] = t[7232] ^ n[7233];
assign t[7234] = t[7233] ^ n[7234];
assign t[7235] = t[7234] ^ n[7235];
assign t[7236] = t[7235] ^ n[7236];
assign t[7237] = t[7236] ^ n[7237];
assign t[7238] = t[7237] ^ n[7238];
assign t[7239] = t[7238] ^ n[7239];
assign t[7240] = t[7239] ^ n[7240];
assign t[7241] = t[7240] ^ n[7241];
assign t[7242] = t[7241] ^ n[7242];
assign t[7243] = t[7242] ^ n[7243];
assign t[7244] = t[7243] ^ n[7244];
assign t[7245] = t[7244] ^ n[7245];
assign t[7246] = t[7245] ^ n[7246];
assign t[7247] = t[7246] ^ n[7247];
assign t[7248] = t[7247] ^ n[7248];
assign t[7249] = t[7248] ^ n[7249];
assign t[7250] = t[7249] ^ n[7250];
assign t[7251] = t[7250] ^ n[7251];
assign t[7252] = t[7251] ^ n[7252];
assign t[7253] = t[7252] ^ n[7253];
assign t[7254] = t[7253] ^ n[7254];
assign t[7255] = t[7254] ^ n[7255];
assign t[7256] = t[7255] ^ n[7256];
assign t[7257] = t[7256] ^ n[7257];
assign t[7258] = t[7257] ^ n[7258];
assign t[7259] = t[7258] ^ n[7259];
assign t[7260] = t[7259] ^ n[7260];
assign t[7261] = t[7260] ^ n[7261];
assign t[7262] = t[7261] ^ n[7262];
assign t[7263] = t[7262] ^ n[7263];
assign t[7264] = t[7263] ^ n[7264];
assign t[7265] = t[7264] ^ n[7265];
assign t[7266] = t[7265] ^ n[7266];
assign t[7267] = t[7266] ^ n[7267];
assign t[7268] = t[7267] ^ n[7268];
assign t[7269] = t[7268] ^ n[7269];
assign t[7270] = t[7269] ^ n[7270];
assign t[7271] = t[7270] ^ n[7271];
assign t[7272] = t[7271] ^ n[7272];
assign t[7273] = t[7272] ^ n[7273];
assign t[7274] = t[7273] ^ n[7274];
assign t[7275] = t[7274] ^ n[7275];
assign t[7276] = t[7275] ^ n[7276];
assign t[7277] = t[7276] ^ n[7277];
assign t[7278] = t[7277] ^ n[7278];
assign t[7279] = t[7278] ^ n[7279];
assign t[7280] = t[7279] ^ n[7280];
assign t[7281] = t[7280] ^ n[7281];
assign t[7282] = t[7281] ^ n[7282];
assign t[7283] = t[7282] ^ n[7283];
assign t[7284] = t[7283] ^ n[7284];
assign t[7285] = t[7284] ^ n[7285];
assign t[7286] = t[7285] ^ n[7286];
assign t[7287] = t[7286] ^ n[7287];
assign t[7288] = t[7287] ^ n[7288];
assign t[7289] = t[7288] ^ n[7289];
assign t[7290] = t[7289] ^ n[7290];
assign t[7291] = t[7290] ^ n[7291];
assign t[7292] = t[7291] ^ n[7292];
assign t[7293] = t[7292] ^ n[7293];
assign t[7294] = t[7293] ^ n[7294];
assign t[7295] = t[7294] ^ n[7295];
assign t[7296] = t[7295] ^ n[7296];
assign t[7297] = t[7296] ^ n[7297];
assign t[7298] = t[7297] ^ n[7298];
assign t[7299] = t[7298] ^ n[7299];
assign t[7300] = t[7299] ^ n[7300];
assign t[7301] = t[7300] ^ n[7301];
assign t[7302] = t[7301] ^ n[7302];
assign t[7303] = t[7302] ^ n[7303];
assign t[7304] = t[7303] ^ n[7304];
assign t[7305] = t[7304] ^ n[7305];
assign t[7306] = t[7305] ^ n[7306];
assign t[7307] = t[7306] ^ n[7307];
assign t[7308] = t[7307] ^ n[7308];
assign t[7309] = t[7308] ^ n[7309];
assign t[7310] = t[7309] ^ n[7310];
assign t[7311] = t[7310] ^ n[7311];
assign t[7312] = t[7311] ^ n[7312];
assign t[7313] = t[7312] ^ n[7313];
assign t[7314] = t[7313] ^ n[7314];
assign t[7315] = t[7314] ^ n[7315];
assign t[7316] = t[7315] ^ n[7316];
assign t[7317] = t[7316] ^ n[7317];
assign t[7318] = t[7317] ^ n[7318];
assign t[7319] = t[7318] ^ n[7319];
assign t[7320] = t[7319] ^ n[7320];
assign t[7321] = t[7320] ^ n[7321];
assign t[7322] = t[7321] ^ n[7322];
assign t[7323] = t[7322] ^ n[7323];
assign t[7324] = t[7323] ^ n[7324];
assign t[7325] = t[7324] ^ n[7325];
assign t[7326] = t[7325] ^ n[7326];
assign t[7327] = t[7326] ^ n[7327];
assign t[7328] = t[7327] ^ n[7328];
assign t[7329] = t[7328] ^ n[7329];
assign t[7330] = t[7329] ^ n[7330];
assign t[7331] = t[7330] ^ n[7331];
assign t[7332] = t[7331] ^ n[7332];
assign t[7333] = t[7332] ^ n[7333];
assign t[7334] = t[7333] ^ n[7334];
assign t[7335] = t[7334] ^ n[7335];
assign t[7336] = t[7335] ^ n[7336];
assign t[7337] = t[7336] ^ n[7337];
assign t[7338] = t[7337] ^ n[7338];
assign t[7339] = t[7338] ^ n[7339];
assign t[7340] = t[7339] ^ n[7340];
assign t[7341] = t[7340] ^ n[7341];
assign t[7342] = t[7341] ^ n[7342];
assign t[7343] = t[7342] ^ n[7343];
assign t[7344] = t[7343] ^ n[7344];
assign t[7345] = t[7344] ^ n[7345];
assign t[7346] = t[7345] ^ n[7346];
assign t[7347] = t[7346] ^ n[7347];
assign t[7348] = t[7347] ^ n[7348];
assign t[7349] = t[7348] ^ n[7349];
assign t[7350] = t[7349] ^ n[7350];
assign t[7351] = t[7350] ^ n[7351];
assign t[7352] = t[7351] ^ n[7352];
assign t[7353] = t[7352] ^ n[7353];
assign t[7354] = t[7353] ^ n[7354];
assign t[7355] = t[7354] ^ n[7355];
assign t[7356] = t[7355] ^ n[7356];
assign t[7357] = t[7356] ^ n[7357];
assign t[7358] = t[7357] ^ n[7358];
assign t[7359] = t[7358] ^ n[7359];
assign t[7360] = t[7359] ^ n[7360];
assign t[7361] = t[7360] ^ n[7361];
assign t[7362] = t[7361] ^ n[7362];
assign t[7363] = t[7362] ^ n[7363];
assign t[7364] = t[7363] ^ n[7364];
assign t[7365] = t[7364] ^ n[7365];
assign t[7366] = t[7365] ^ n[7366];
assign t[7367] = t[7366] ^ n[7367];
assign t[7368] = t[7367] ^ n[7368];
assign t[7369] = t[7368] ^ n[7369];
assign t[7370] = t[7369] ^ n[7370];
assign t[7371] = t[7370] ^ n[7371];
assign t[7372] = t[7371] ^ n[7372];
assign t[7373] = t[7372] ^ n[7373];
assign t[7374] = t[7373] ^ n[7374];
assign t[7375] = t[7374] ^ n[7375];
assign t[7376] = t[7375] ^ n[7376];
assign t[7377] = t[7376] ^ n[7377];
assign t[7378] = t[7377] ^ n[7378];
assign t[7379] = t[7378] ^ n[7379];
assign t[7380] = t[7379] ^ n[7380];
assign t[7381] = t[7380] ^ n[7381];
assign t[7382] = t[7381] ^ n[7382];
assign t[7383] = t[7382] ^ n[7383];
assign t[7384] = t[7383] ^ n[7384];
assign t[7385] = t[7384] ^ n[7385];
assign t[7386] = t[7385] ^ n[7386];
assign t[7387] = t[7386] ^ n[7387];
assign t[7388] = t[7387] ^ n[7388];
assign t[7389] = t[7388] ^ n[7389];
assign t[7390] = t[7389] ^ n[7390];
assign t[7391] = t[7390] ^ n[7391];
assign t[7392] = t[7391] ^ n[7392];
assign t[7393] = t[7392] ^ n[7393];
assign t[7394] = t[7393] ^ n[7394];
assign t[7395] = t[7394] ^ n[7395];
assign t[7396] = t[7395] ^ n[7396];
assign t[7397] = t[7396] ^ n[7397];
assign t[7398] = t[7397] ^ n[7398];
assign t[7399] = t[7398] ^ n[7399];
assign t[7400] = t[7399] ^ n[7400];
assign t[7401] = t[7400] ^ n[7401];
assign t[7402] = t[7401] ^ n[7402];
assign t[7403] = t[7402] ^ n[7403];
assign t[7404] = t[7403] ^ n[7404];
assign t[7405] = t[7404] ^ n[7405];
assign t[7406] = t[7405] ^ n[7406];
assign t[7407] = t[7406] ^ n[7407];
assign t[7408] = t[7407] ^ n[7408];
assign t[7409] = t[7408] ^ n[7409];
assign t[7410] = t[7409] ^ n[7410];
assign t[7411] = t[7410] ^ n[7411];
assign t[7412] = t[7411] ^ n[7412];
assign t[7413] = t[7412] ^ n[7413];
assign t[7414] = t[7413] ^ n[7414];
assign t[7415] = t[7414] ^ n[7415];
assign t[7416] = t[7415] ^ n[7416];
assign t[7417] = t[7416] ^ n[7417];
assign t[7418] = t[7417] ^ n[7418];
assign t[7419] = t[7418] ^ n[7419];
assign t[7420] = t[7419] ^ n[7420];
assign t[7421] = t[7420] ^ n[7421];
assign t[7422] = t[7421] ^ n[7422];
assign t[7423] = t[7422] ^ n[7423];
assign t[7424] = t[7423] ^ n[7424];
assign t[7425] = t[7424] ^ n[7425];
assign t[7426] = t[7425] ^ n[7426];
assign t[7427] = t[7426] ^ n[7427];
assign t[7428] = t[7427] ^ n[7428];
assign t[7429] = t[7428] ^ n[7429];
assign t[7430] = t[7429] ^ n[7430];
assign t[7431] = t[7430] ^ n[7431];
assign t[7432] = t[7431] ^ n[7432];
assign t[7433] = t[7432] ^ n[7433];
assign t[7434] = t[7433] ^ n[7434];
assign t[7435] = t[7434] ^ n[7435];
assign t[7436] = t[7435] ^ n[7436];
assign t[7437] = t[7436] ^ n[7437];
assign t[7438] = t[7437] ^ n[7438];
assign t[7439] = t[7438] ^ n[7439];
assign t[7440] = t[7439] ^ n[7440];
assign t[7441] = t[7440] ^ n[7441];
assign t[7442] = t[7441] ^ n[7442];
assign t[7443] = t[7442] ^ n[7443];
assign t[7444] = t[7443] ^ n[7444];
assign t[7445] = t[7444] ^ n[7445];
assign t[7446] = t[7445] ^ n[7446];
assign t[7447] = t[7446] ^ n[7447];
assign t[7448] = t[7447] ^ n[7448];
assign t[7449] = t[7448] ^ n[7449];
assign t[7450] = t[7449] ^ n[7450];
assign t[7451] = t[7450] ^ n[7451];
assign t[7452] = t[7451] ^ n[7452];
assign t[7453] = t[7452] ^ n[7453];
assign t[7454] = t[7453] ^ n[7454];
assign t[7455] = t[7454] ^ n[7455];
assign t[7456] = t[7455] ^ n[7456];
assign t[7457] = t[7456] ^ n[7457];
assign t[7458] = t[7457] ^ n[7458];
assign t[7459] = t[7458] ^ n[7459];
assign t[7460] = t[7459] ^ n[7460];
assign t[7461] = t[7460] ^ n[7461];
assign t[7462] = t[7461] ^ n[7462];
assign t[7463] = t[7462] ^ n[7463];
assign t[7464] = t[7463] ^ n[7464];
assign t[7465] = t[7464] ^ n[7465];
assign t[7466] = t[7465] ^ n[7466];
assign t[7467] = t[7466] ^ n[7467];
assign t[7468] = t[7467] ^ n[7468];
assign t[7469] = t[7468] ^ n[7469];
assign t[7470] = t[7469] ^ n[7470];
assign t[7471] = t[7470] ^ n[7471];
assign t[7472] = t[7471] ^ n[7472];
assign t[7473] = t[7472] ^ n[7473];
assign t[7474] = t[7473] ^ n[7474];
assign t[7475] = t[7474] ^ n[7475];
assign t[7476] = t[7475] ^ n[7476];
assign t[7477] = t[7476] ^ n[7477];
assign t[7478] = t[7477] ^ n[7478];
assign t[7479] = t[7478] ^ n[7479];
assign t[7480] = t[7479] ^ n[7480];
assign t[7481] = t[7480] ^ n[7481];
assign t[7482] = t[7481] ^ n[7482];
assign t[7483] = t[7482] ^ n[7483];
assign t[7484] = t[7483] ^ n[7484];
assign t[7485] = t[7484] ^ n[7485];
assign t[7486] = t[7485] ^ n[7486];
assign t[7487] = t[7486] ^ n[7487];
assign t[7488] = t[7487] ^ n[7488];
assign t[7489] = t[7488] ^ n[7489];
assign t[7490] = t[7489] ^ n[7490];
assign t[7491] = t[7490] ^ n[7491];
assign t[7492] = t[7491] ^ n[7492];
assign t[7493] = t[7492] ^ n[7493];
assign t[7494] = t[7493] ^ n[7494];
assign t[7495] = t[7494] ^ n[7495];
assign t[7496] = t[7495] ^ n[7496];
assign t[7497] = t[7496] ^ n[7497];
assign t[7498] = t[7497] ^ n[7498];
assign t[7499] = t[7498] ^ n[7499];
assign t[7500] = t[7499] ^ n[7500];
assign t[7501] = t[7500] ^ n[7501];
assign t[7502] = t[7501] ^ n[7502];
assign t[7503] = t[7502] ^ n[7503];
assign t[7504] = t[7503] ^ n[7504];
assign t[7505] = t[7504] ^ n[7505];
assign t[7506] = t[7505] ^ n[7506];
assign t[7507] = t[7506] ^ n[7507];
assign t[7508] = t[7507] ^ n[7508];
assign t[7509] = t[7508] ^ n[7509];
assign t[7510] = t[7509] ^ n[7510];
assign t[7511] = t[7510] ^ n[7511];
assign t[7512] = t[7511] ^ n[7512];
assign t[7513] = t[7512] ^ n[7513];
assign t[7514] = t[7513] ^ n[7514];
assign t[7515] = t[7514] ^ n[7515];
assign t[7516] = t[7515] ^ n[7516];
assign t[7517] = t[7516] ^ n[7517];
assign t[7518] = t[7517] ^ n[7518];
assign t[7519] = t[7518] ^ n[7519];
assign t[7520] = t[7519] ^ n[7520];
assign t[7521] = t[7520] ^ n[7521];
assign t[7522] = t[7521] ^ n[7522];
assign t[7523] = t[7522] ^ n[7523];
assign t[7524] = t[7523] ^ n[7524];
assign t[7525] = t[7524] ^ n[7525];
assign t[7526] = t[7525] ^ n[7526];
assign t[7527] = t[7526] ^ n[7527];
assign t[7528] = t[7527] ^ n[7528];
assign t[7529] = t[7528] ^ n[7529];
assign t[7530] = t[7529] ^ n[7530];
assign t[7531] = t[7530] ^ n[7531];
assign t[7532] = t[7531] ^ n[7532];
assign t[7533] = t[7532] ^ n[7533];
assign t[7534] = t[7533] ^ n[7534];
assign t[7535] = t[7534] ^ n[7535];
assign t[7536] = t[7535] ^ n[7536];
assign t[7537] = t[7536] ^ n[7537];
assign t[7538] = t[7537] ^ n[7538];
assign t[7539] = t[7538] ^ n[7539];
assign t[7540] = t[7539] ^ n[7540];
assign t[7541] = t[7540] ^ n[7541];
assign t[7542] = t[7541] ^ n[7542];
assign t[7543] = t[7542] ^ n[7543];
assign t[7544] = t[7543] ^ n[7544];
assign t[7545] = t[7544] ^ n[7545];
assign t[7546] = t[7545] ^ n[7546];
assign t[7547] = t[7546] ^ n[7547];
assign t[7548] = t[7547] ^ n[7548];
assign t[7549] = t[7548] ^ n[7549];
assign t[7550] = t[7549] ^ n[7550];
assign t[7551] = t[7550] ^ n[7551];
assign t[7552] = t[7551] ^ n[7552];
assign t[7553] = t[7552] ^ n[7553];
assign t[7554] = t[7553] ^ n[7554];
assign t[7555] = t[7554] ^ n[7555];
assign t[7556] = t[7555] ^ n[7556];
assign t[7557] = t[7556] ^ n[7557];
assign t[7558] = t[7557] ^ n[7558];
assign t[7559] = t[7558] ^ n[7559];
assign t[7560] = t[7559] ^ n[7560];
assign t[7561] = t[7560] ^ n[7561];
assign t[7562] = t[7561] ^ n[7562];
assign t[7563] = t[7562] ^ n[7563];
assign t[7564] = t[7563] ^ n[7564];
assign t[7565] = t[7564] ^ n[7565];
assign t[7566] = t[7565] ^ n[7566];
assign t[7567] = t[7566] ^ n[7567];
assign t[7568] = t[7567] ^ n[7568];
assign t[7569] = t[7568] ^ n[7569];
assign t[7570] = t[7569] ^ n[7570];
assign t[7571] = t[7570] ^ n[7571];
assign t[7572] = t[7571] ^ n[7572];
assign t[7573] = t[7572] ^ n[7573];
assign t[7574] = t[7573] ^ n[7574];
assign t[7575] = t[7574] ^ n[7575];
assign t[7576] = t[7575] ^ n[7576];
assign t[7577] = t[7576] ^ n[7577];
assign t[7578] = t[7577] ^ n[7578];
assign t[7579] = t[7578] ^ n[7579];
assign t[7580] = t[7579] ^ n[7580];
assign t[7581] = t[7580] ^ n[7581];
assign t[7582] = t[7581] ^ n[7582];
assign t[7583] = t[7582] ^ n[7583];
assign t[7584] = t[7583] ^ n[7584];
assign t[7585] = t[7584] ^ n[7585];
assign t[7586] = t[7585] ^ n[7586];
assign t[7587] = t[7586] ^ n[7587];
assign t[7588] = t[7587] ^ n[7588];
assign t[7589] = t[7588] ^ n[7589];
assign t[7590] = t[7589] ^ n[7590];
assign t[7591] = t[7590] ^ n[7591];
assign t[7592] = t[7591] ^ n[7592];
assign t[7593] = t[7592] ^ n[7593];
assign t[7594] = t[7593] ^ n[7594];
assign t[7595] = t[7594] ^ n[7595];
assign t[7596] = t[7595] ^ n[7596];
assign t[7597] = t[7596] ^ n[7597];
assign t[7598] = t[7597] ^ n[7598];
assign t[7599] = t[7598] ^ n[7599];
assign t[7600] = t[7599] ^ n[7600];
assign t[7601] = t[7600] ^ n[7601];
assign t[7602] = t[7601] ^ n[7602];
assign t[7603] = t[7602] ^ n[7603];
assign t[7604] = t[7603] ^ n[7604];
assign t[7605] = t[7604] ^ n[7605];
assign t[7606] = t[7605] ^ n[7606];
assign t[7607] = t[7606] ^ n[7607];
assign t[7608] = t[7607] ^ n[7608];
assign t[7609] = t[7608] ^ n[7609];
assign t[7610] = t[7609] ^ n[7610];
assign t[7611] = t[7610] ^ n[7611];
assign t[7612] = t[7611] ^ n[7612];
assign t[7613] = t[7612] ^ n[7613];
assign t[7614] = t[7613] ^ n[7614];
assign t[7615] = t[7614] ^ n[7615];
assign t[7616] = t[7615] ^ n[7616];
assign t[7617] = t[7616] ^ n[7617];
assign t[7618] = t[7617] ^ n[7618];
assign t[7619] = t[7618] ^ n[7619];
assign t[7620] = t[7619] ^ n[7620];
assign t[7621] = t[7620] ^ n[7621];
assign t[7622] = t[7621] ^ n[7622];
assign t[7623] = t[7622] ^ n[7623];
assign t[7624] = t[7623] ^ n[7624];
assign t[7625] = t[7624] ^ n[7625];
assign t[7626] = t[7625] ^ n[7626];
assign t[7627] = t[7626] ^ n[7627];
assign t[7628] = t[7627] ^ n[7628];
assign t[7629] = t[7628] ^ n[7629];
assign t[7630] = t[7629] ^ n[7630];
assign t[7631] = t[7630] ^ n[7631];
assign t[7632] = t[7631] ^ n[7632];
assign t[7633] = t[7632] ^ n[7633];
assign t[7634] = t[7633] ^ n[7634];
assign t[7635] = t[7634] ^ n[7635];
assign t[7636] = t[7635] ^ n[7636];
assign t[7637] = t[7636] ^ n[7637];
assign t[7638] = t[7637] ^ n[7638];
assign t[7639] = t[7638] ^ n[7639];
assign t[7640] = t[7639] ^ n[7640];
assign t[7641] = t[7640] ^ n[7641];
assign t[7642] = t[7641] ^ n[7642];
assign t[7643] = t[7642] ^ n[7643];
assign t[7644] = t[7643] ^ n[7644];
assign t[7645] = t[7644] ^ n[7645];
assign t[7646] = t[7645] ^ n[7646];
assign t[7647] = t[7646] ^ n[7647];
assign t[7648] = t[7647] ^ n[7648];
assign t[7649] = t[7648] ^ n[7649];
assign t[7650] = t[7649] ^ n[7650];
assign t[7651] = t[7650] ^ n[7651];
assign t[7652] = t[7651] ^ n[7652];
assign t[7653] = t[7652] ^ n[7653];
assign t[7654] = t[7653] ^ n[7654];
assign t[7655] = t[7654] ^ n[7655];
assign t[7656] = t[7655] ^ n[7656];
assign t[7657] = t[7656] ^ n[7657];
assign t[7658] = t[7657] ^ n[7658];
assign t[7659] = t[7658] ^ n[7659];
assign t[7660] = t[7659] ^ n[7660];
assign t[7661] = t[7660] ^ n[7661];
assign t[7662] = t[7661] ^ n[7662];
assign t[7663] = t[7662] ^ n[7663];
assign t[7664] = t[7663] ^ n[7664];
assign t[7665] = t[7664] ^ n[7665];
assign t[7666] = t[7665] ^ n[7666];
assign t[7667] = t[7666] ^ n[7667];
assign t[7668] = t[7667] ^ n[7668];
assign t[7669] = t[7668] ^ n[7669];
assign t[7670] = t[7669] ^ n[7670];
assign t[7671] = t[7670] ^ n[7671];
assign t[7672] = t[7671] ^ n[7672];
assign t[7673] = t[7672] ^ n[7673];
assign t[7674] = t[7673] ^ n[7674];
assign t[7675] = t[7674] ^ n[7675];
assign t[7676] = t[7675] ^ n[7676];
assign t[7677] = t[7676] ^ n[7677];
assign t[7678] = t[7677] ^ n[7678];
assign t[7679] = t[7678] ^ n[7679];
assign t[7680] = t[7679] ^ n[7680];
assign t[7681] = t[7680] ^ n[7681];
assign t[7682] = t[7681] ^ n[7682];
assign t[7683] = t[7682] ^ n[7683];
assign t[7684] = t[7683] ^ n[7684];
assign t[7685] = t[7684] ^ n[7685];
assign t[7686] = t[7685] ^ n[7686];
assign t[7687] = t[7686] ^ n[7687];
assign t[7688] = t[7687] ^ n[7688];
assign t[7689] = t[7688] ^ n[7689];
assign t[7690] = t[7689] ^ n[7690];
assign t[7691] = t[7690] ^ n[7691];
assign t[7692] = t[7691] ^ n[7692];
assign t[7693] = t[7692] ^ n[7693];
assign t[7694] = t[7693] ^ n[7694];
assign t[7695] = t[7694] ^ n[7695];
assign t[7696] = t[7695] ^ n[7696];
assign t[7697] = t[7696] ^ n[7697];
assign t[7698] = t[7697] ^ n[7698];
assign t[7699] = t[7698] ^ n[7699];
assign t[7700] = t[7699] ^ n[7700];
assign t[7701] = t[7700] ^ n[7701];
assign t[7702] = t[7701] ^ n[7702];
assign t[7703] = t[7702] ^ n[7703];
assign t[7704] = t[7703] ^ n[7704];
assign t[7705] = t[7704] ^ n[7705];
assign t[7706] = t[7705] ^ n[7706];
assign t[7707] = t[7706] ^ n[7707];
assign t[7708] = t[7707] ^ n[7708];
assign t[7709] = t[7708] ^ n[7709];
assign t[7710] = t[7709] ^ n[7710];
assign t[7711] = t[7710] ^ n[7711];
assign t[7712] = t[7711] ^ n[7712];
assign t[7713] = t[7712] ^ n[7713];
assign t[7714] = t[7713] ^ n[7714];
assign t[7715] = t[7714] ^ n[7715];
assign t[7716] = t[7715] ^ n[7716];
assign t[7717] = t[7716] ^ n[7717];
assign t[7718] = t[7717] ^ n[7718];
assign t[7719] = t[7718] ^ n[7719];
assign t[7720] = t[7719] ^ n[7720];
assign t[7721] = t[7720] ^ n[7721];
assign t[7722] = t[7721] ^ n[7722];
assign t[7723] = t[7722] ^ n[7723];
assign t[7724] = t[7723] ^ n[7724];
assign t[7725] = t[7724] ^ n[7725];
assign t[7726] = t[7725] ^ n[7726];
assign t[7727] = t[7726] ^ n[7727];
assign t[7728] = t[7727] ^ n[7728];
assign t[7729] = t[7728] ^ n[7729];
assign t[7730] = t[7729] ^ n[7730];
assign t[7731] = t[7730] ^ n[7731];
assign t[7732] = t[7731] ^ n[7732];
assign t[7733] = t[7732] ^ n[7733];
assign t[7734] = t[7733] ^ n[7734];
assign t[7735] = t[7734] ^ n[7735];
assign t[7736] = t[7735] ^ n[7736];
assign t[7737] = t[7736] ^ n[7737];
assign t[7738] = t[7737] ^ n[7738];
assign t[7739] = t[7738] ^ n[7739];
assign t[7740] = t[7739] ^ n[7740];
assign t[7741] = t[7740] ^ n[7741];
assign t[7742] = t[7741] ^ n[7742];
assign t[7743] = t[7742] ^ n[7743];
assign t[7744] = t[7743] ^ n[7744];
assign t[7745] = t[7744] ^ n[7745];
assign t[7746] = t[7745] ^ n[7746];
assign t[7747] = t[7746] ^ n[7747];
assign t[7748] = t[7747] ^ n[7748];
assign t[7749] = t[7748] ^ n[7749];
assign t[7750] = t[7749] ^ n[7750];
assign t[7751] = t[7750] ^ n[7751];
assign t[7752] = t[7751] ^ n[7752];
assign t[7753] = t[7752] ^ n[7753];
assign t[7754] = t[7753] ^ n[7754];
assign t[7755] = t[7754] ^ n[7755];
assign t[7756] = t[7755] ^ n[7756];
assign t[7757] = t[7756] ^ n[7757];
assign t[7758] = t[7757] ^ n[7758];
assign t[7759] = t[7758] ^ n[7759];
assign t[7760] = t[7759] ^ n[7760];
assign t[7761] = t[7760] ^ n[7761];
assign t[7762] = t[7761] ^ n[7762];
assign t[7763] = t[7762] ^ n[7763];
assign t[7764] = t[7763] ^ n[7764];
assign t[7765] = t[7764] ^ n[7765];
assign t[7766] = t[7765] ^ n[7766];
assign t[7767] = t[7766] ^ n[7767];
assign t[7768] = t[7767] ^ n[7768];
assign t[7769] = t[7768] ^ n[7769];
assign t[7770] = t[7769] ^ n[7770];
assign t[7771] = t[7770] ^ n[7771];
assign t[7772] = t[7771] ^ n[7772];
assign t[7773] = t[7772] ^ n[7773];
assign t[7774] = t[7773] ^ n[7774];
assign t[7775] = t[7774] ^ n[7775];
assign t[7776] = t[7775] ^ n[7776];
assign t[7777] = t[7776] ^ n[7777];
assign t[7778] = t[7777] ^ n[7778];
assign t[7779] = t[7778] ^ n[7779];
assign t[7780] = t[7779] ^ n[7780];
assign t[7781] = t[7780] ^ n[7781];
assign t[7782] = t[7781] ^ n[7782];
assign t[7783] = t[7782] ^ n[7783];
assign t[7784] = t[7783] ^ n[7784];
assign t[7785] = t[7784] ^ n[7785];
assign t[7786] = t[7785] ^ n[7786];
assign t[7787] = t[7786] ^ n[7787];
assign t[7788] = t[7787] ^ n[7788];
assign t[7789] = t[7788] ^ n[7789];
assign t[7790] = t[7789] ^ n[7790];
assign t[7791] = t[7790] ^ n[7791];
assign t[7792] = t[7791] ^ n[7792];
assign t[7793] = t[7792] ^ n[7793];
assign t[7794] = t[7793] ^ n[7794];
assign t[7795] = t[7794] ^ n[7795];
assign t[7796] = t[7795] ^ n[7796];
assign t[7797] = t[7796] ^ n[7797];
assign t[7798] = t[7797] ^ n[7798];
assign t[7799] = t[7798] ^ n[7799];
assign t[7800] = t[7799] ^ n[7800];
assign t[7801] = t[7800] ^ n[7801];
assign t[7802] = t[7801] ^ n[7802];
assign t[7803] = t[7802] ^ n[7803];
assign t[7804] = t[7803] ^ n[7804];
assign t[7805] = t[7804] ^ n[7805];
assign t[7806] = t[7805] ^ n[7806];
assign t[7807] = t[7806] ^ n[7807];
assign t[7808] = t[7807] ^ n[7808];
assign t[7809] = t[7808] ^ n[7809];
assign t[7810] = t[7809] ^ n[7810];
assign t[7811] = t[7810] ^ n[7811];
assign t[7812] = t[7811] ^ n[7812];
assign t[7813] = t[7812] ^ n[7813];
assign t[7814] = t[7813] ^ n[7814];
assign t[7815] = t[7814] ^ n[7815];
assign t[7816] = t[7815] ^ n[7816];
assign t[7817] = t[7816] ^ n[7817];
assign t[7818] = t[7817] ^ n[7818];
assign t[7819] = t[7818] ^ n[7819];
assign t[7820] = t[7819] ^ n[7820];
assign t[7821] = t[7820] ^ n[7821];
assign t[7822] = t[7821] ^ n[7822];
assign t[7823] = t[7822] ^ n[7823];
assign t[7824] = t[7823] ^ n[7824];
assign t[7825] = t[7824] ^ n[7825];
assign t[7826] = t[7825] ^ n[7826];
assign t[7827] = t[7826] ^ n[7827];
assign t[7828] = t[7827] ^ n[7828];
assign t[7829] = t[7828] ^ n[7829];
assign t[7830] = t[7829] ^ n[7830];
assign t[7831] = t[7830] ^ n[7831];
assign t[7832] = t[7831] ^ n[7832];
assign t[7833] = t[7832] ^ n[7833];
assign t[7834] = t[7833] ^ n[7834];
assign t[7835] = t[7834] ^ n[7835];
assign t[7836] = t[7835] ^ n[7836];
assign t[7837] = t[7836] ^ n[7837];
assign t[7838] = t[7837] ^ n[7838];
assign t[7839] = t[7838] ^ n[7839];
assign t[7840] = t[7839] ^ n[7840];
assign t[7841] = t[7840] ^ n[7841];
assign t[7842] = t[7841] ^ n[7842];
assign t[7843] = t[7842] ^ n[7843];
assign t[7844] = t[7843] ^ n[7844];
assign t[7845] = t[7844] ^ n[7845];
assign t[7846] = t[7845] ^ n[7846];
assign t[7847] = t[7846] ^ n[7847];
assign t[7848] = t[7847] ^ n[7848];
assign t[7849] = t[7848] ^ n[7849];
assign t[7850] = t[7849] ^ n[7850];
assign t[7851] = t[7850] ^ n[7851];
assign t[7852] = t[7851] ^ n[7852];
assign t[7853] = t[7852] ^ n[7853];
assign t[7854] = t[7853] ^ n[7854];
assign t[7855] = t[7854] ^ n[7855];
assign t[7856] = t[7855] ^ n[7856];
assign t[7857] = t[7856] ^ n[7857];
assign t[7858] = t[7857] ^ n[7858];
assign t[7859] = t[7858] ^ n[7859];
assign t[7860] = t[7859] ^ n[7860];
assign t[7861] = t[7860] ^ n[7861];
assign t[7862] = t[7861] ^ n[7862];
assign t[7863] = t[7862] ^ n[7863];
assign t[7864] = t[7863] ^ n[7864];
assign t[7865] = t[7864] ^ n[7865];
assign t[7866] = t[7865] ^ n[7866];
assign t[7867] = t[7866] ^ n[7867];
assign t[7868] = t[7867] ^ n[7868];
assign t[7869] = t[7868] ^ n[7869];
assign t[7870] = t[7869] ^ n[7870];
assign t[7871] = t[7870] ^ n[7871];
assign t[7872] = t[7871] ^ n[7872];
assign t[7873] = t[7872] ^ n[7873];
assign t[7874] = t[7873] ^ n[7874];
assign t[7875] = t[7874] ^ n[7875];
assign t[7876] = t[7875] ^ n[7876];
assign t[7877] = t[7876] ^ n[7877];
assign t[7878] = t[7877] ^ n[7878];
assign t[7879] = t[7878] ^ n[7879];
assign t[7880] = t[7879] ^ n[7880];
assign t[7881] = t[7880] ^ n[7881];
assign t[7882] = t[7881] ^ n[7882];
assign t[7883] = t[7882] ^ n[7883];
assign t[7884] = t[7883] ^ n[7884];
assign t[7885] = t[7884] ^ n[7885];
assign t[7886] = t[7885] ^ n[7886];
assign t[7887] = t[7886] ^ n[7887];
assign t[7888] = t[7887] ^ n[7888];
assign t[7889] = t[7888] ^ n[7889];
assign t[7890] = t[7889] ^ n[7890];
assign t[7891] = t[7890] ^ n[7891];
assign t[7892] = t[7891] ^ n[7892];
assign t[7893] = t[7892] ^ n[7893];
assign t[7894] = t[7893] ^ n[7894];
assign t[7895] = t[7894] ^ n[7895];
assign t[7896] = t[7895] ^ n[7896];
assign t[7897] = t[7896] ^ n[7897];
assign t[7898] = t[7897] ^ n[7898];
assign t[7899] = t[7898] ^ n[7899];
assign t[7900] = t[7899] ^ n[7900];
assign t[7901] = t[7900] ^ n[7901];
assign t[7902] = t[7901] ^ n[7902];
assign t[7903] = t[7902] ^ n[7903];
assign t[7904] = t[7903] ^ n[7904];
assign t[7905] = t[7904] ^ n[7905];
assign t[7906] = t[7905] ^ n[7906];
assign t[7907] = t[7906] ^ n[7907];
assign t[7908] = t[7907] ^ n[7908];
assign t[7909] = t[7908] ^ n[7909];
assign t[7910] = t[7909] ^ n[7910];
assign t[7911] = t[7910] ^ n[7911];
assign t[7912] = t[7911] ^ n[7912];
assign t[7913] = t[7912] ^ n[7913];
assign t[7914] = t[7913] ^ n[7914];
assign t[7915] = t[7914] ^ n[7915];
assign t[7916] = t[7915] ^ n[7916];
assign t[7917] = t[7916] ^ n[7917];
assign t[7918] = t[7917] ^ n[7918];
assign t[7919] = t[7918] ^ n[7919];
assign t[7920] = t[7919] ^ n[7920];
assign t[7921] = t[7920] ^ n[7921];
assign t[7922] = t[7921] ^ n[7922];
assign t[7923] = t[7922] ^ n[7923];
assign t[7924] = t[7923] ^ n[7924];
assign t[7925] = t[7924] ^ n[7925];
assign t[7926] = t[7925] ^ n[7926];
assign t[7927] = t[7926] ^ n[7927];
assign t[7928] = t[7927] ^ n[7928];
assign t[7929] = t[7928] ^ n[7929];
assign t[7930] = t[7929] ^ n[7930];
assign t[7931] = t[7930] ^ n[7931];
assign t[7932] = t[7931] ^ n[7932];
assign t[7933] = t[7932] ^ n[7933];
assign t[7934] = t[7933] ^ n[7934];
assign t[7935] = t[7934] ^ n[7935];
assign t[7936] = t[7935] ^ n[7936];
assign t[7937] = t[7936] ^ n[7937];
assign t[7938] = t[7937] ^ n[7938];
assign t[7939] = t[7938] ^ n[7939];
assign t[7940] = t[7939] ^ n[7940];
assign t[7941] = t[7940] ^ n[7941];
assign t[7942] = t[7941] ^ n[7942];
assign t[7943] = t[7942] ^ n[7943];
assign t[7944] = t[7943] ^ n[7944];
assign t[7945] = t[7944] ^ n[7945];
assign t[7946] = t[7945] ^ n[7946];
assign t[7947] = t[7946] ^ n[7947];
assign t[7948] = t[7947] ^ n[7948];
assign t[7949] = t[7948] ^ n[7949];
assign t[7950] = t[7949] ^ n[7950];
assign t[7951] = t[7950] ^ n[7951];
assign t[7952] = t[7951] ^ n[7952];
assign t[7953] = t[7952] ^ n[7953];
assign t[7954] = t[7953] ^ n[7954];
assign t[7955] = t[7954] ^ n[7955];
assign t[7956] = t[7955] ^ n[7956];
assign t[7957] = t[7956] ^ n[7957];
assign t[7958] = t[7957] ^ n[7958];
assign t[7959] = t[7958] ^ n[7959];
assign t[7960] = t[7959] ^ n[7960];
assign t[7961] = t[7960] ^ n[7961];
assign t[7962] = t[7961] ^ n[7962];
assign t[7963] = t[7962] ^ n[7963];
assign t[7964] = t[7963] ^ n[7964];
assign t[7965] = t[7964] ^ n[7965];
assign t[7966] = t[7965] ^ n[7966];
assign t[7967] = t[7966] ^ n[7967];
assign t[7968] = t[7967] ^ n[7968];
assign t[7969] = t[7968] ^ n[7969];
assign t[7970] = t[7969] ^ n[7970];
assign t[7971] = t[7970] ^ n[7971];
assign t[7972] = t[7971] ^ n[7972];
assign t[7973] = t[7972] ^ n[7973];
assign t[7974] = t[7973] ^ n[7974];
assign t[7975] = t[7974] ^ n[7975];
assign t[7976] = t[7975] ^ n[7976];
assign t[7977] = t[7976] ^ n[7977];
assign t[7978] = t[7977] ^ n[7978];
assign t[7979] = t[7978] ^ n[7979];
assign t[7980] = t[7979] ^ n[7980];
assign t[7981] = t[7980] ^ n[7981];
assign t[7982] = t[7981] ^ n[7982];
assign t[7983] = t[7982] ^ n[7983];
assign t[7984] = t[7983] ^ n[7984];
assign t[7985] = t[7984] ^ n[7985];
assign t[7986] = t[7985] ^ n[7986];
assign t[7987] = t[7986] ^ n[7987];
assign t[7988] = t[7987] ^ n[7988];
assign t[7989] = t[7988] ^ n[7989];
assign t[7990] = t[7989] ^ n[7990];
assign t[7991] = t[7990] ^ n[7991];
assign t[7992] = t[7991] ^ n[7992];
assign t[7993] = t[7992] ^ n[7993];
assign t[7994] = t[7993] ^ n[7994];
assign t[7995] = t[7994] ^ n[7995];
assign t[7996] = t[7995] ^ n[7996];
assign t[7997] = t[7996] ^ n[7997];
assign t[7998] = t[7997] ^ n[7998];
assign t[7999] = t[7998] ^ n[7999];
assign t[8000] = t[7999] ^ n[8000];
assign t[8001] = t[8000] ^ n[8001];
assign t[8002] = t[8001] ^ n[8002];
assign t[8003] = t[8002] ^ n[8003];
assign t[8004] = t[8003] ^ n[8004];
assign t[8005] = t[8004] ^ n[8005];
assign t[8006] = t[8005] ^ n[8006];
assign t[8007] = t[8006] ^ n[8007];
assign t[8008] = t[8007] ^ n[8008];
assign t[8009] = t[8008] ^ n[8009];
assign t[8010] = t[8009] ^ n[8010];
assign t[8011] = t[8010] ^ n[8011];
assign t[8012] = t[8011] ^ n[8012];
assign t[8013] = t[8012] ^ n[8013];
assign t[8014] = t[8013] ^ n[8014];
assign t[8015] = t[8014] ^ n[8015];
assign t[8016] = t[8015] ^ n[8016];
assign t[8017] = t[8016] ^ n[8017];
assign t[8018] = t[8017] ^ n[8018];
assign t[8019] = t[8018] ^ n[8019];
assign t[8020] = t[8019] ^ n[8020];
assign t[8021] = t[8020] ^ n[8021];
assign t[8022] = t[8021] ^ n[8022];
assign t[8023] = t[8022] ^ n[8023];
assign t[8024] = t[8023] ^ n[8024];
assign t[8025] = t[8024] ^ n[8025];
assign t[8026] = t[8025] ^ n[8026];
assign t[8027] = t[8026] ^ n[8027];
assign t[8028] = t[8027] ^ n[8028];
assign t[8029] = t[8028] ^ n[8029];
assign t[8030] = t[8029] ^ n[8030];
assign t[8031] = t[8030] ^ n[8031];
assign t[8032] = t[8031] ^ n[8032];
assign t[8033] = t[8032] ^ n[8033];
assign t[8034] = t[8033] ^ n[8034];
assign t[8035] = t[8034] ^ n[8035];
assign t[8036] = t[8035] ^ n[8036];
assign t[8037] = t[8036] ^ n[8037];
assign t[8038] = t[8037] ^ n[8038];
assign t[8039] = t[8038] ^ n[8039];
assign t[8040] = t[8039] ^ n[8040];
assign t[8041] = t[8040] ^ n[8041];
assign t[8042] = t[8041] ^ n[8042];
assign t[8043] = t[8042] ^ n[8043];
assign t[8044] = t[8043] ^ n[8044];
assign t[8045] = t[8044] ^ n[8045];
assign t[8046] = t[8045] ^ n[8046];
assign t[8047] = t[8046] ^ n[8047];
assign t[8048] = t[8047] ^ n[8048];
assign t[8049] = t[8048] ^ n[8049];
assign t[8050] = t[8049] ^ n[8050];
assign t[8051] = t[8050] ^ n[8051];
assign t[8052] = t[8051] ^ n[8052];
assign t[8053] = t[8052] ^ n[8053];
assign t[8054] = t[8053] ^ n[8054];
assign t[8055] = t[8054] ^ n[8055];
assign t[8056] = t[8055] ^ n[8056];
assign t[8057] = t[8056] ^ n[8057];
assign t[8058] = t[8057] ^ n[8058];
assign t[8059] = t[8058] ^ n[8059];
assign t[8060] = t[8059] ^ n[8060];
assign t[8061] = t[8060] ^ n[8061];
assign t[8062] = t[8061] ^ n[8062];
assign t[8063] = t[8062] ^ n[8063];
assign t[8064] = t[8063] ^ n[8064];
assign t[8065] = t[8064] ^ n[8065];
assign t[8066] = t[8065] ^ n[8066];
assign t[8067] = t[8066] ^ n[8067];
assign t[8068] = t[8067] ^ n[8068];
assign t[8069] = t[8068] ^ n[8069];
assign t[8070] = t[8069] ^ n[8070];
assign t[8071] = t[8070] ^ n[8071];
assign t[8072] = t[8071] ^ n[8072];
assign t[8073] = t[8072] ^ n[8073];
assign t[8074] = t[8073] ^ n[8074];
assign t[8075] = t[8074] ^ n[8075];
assign t[8076] = t[8075] ^ n[8076];
assign t[8077] = t[8076] ^ n[8077];
assign t[8078] = t[8077] ^ n[8078];
assign t[8079] = t[8078] ^ n[8079];
assign t[8080] = t[8079] ^ n[8080];
assign t[8081] = t[8080] ^ n[8081];
assign t[8082] = t[8081] ^ n[8082];
assign t[8083] = t[8082] ^ n[8083];
assign t[8084] = t[8083] ^ n[8084];
assign t[8085] = t[8084] ^ n[8085];
assign t[8086] = t[8085] ^ n[8086];
assign t[8087] = t[8086] ^ n[8087];
assign t[8088] = t[8087] ^ n[8088];
assign t[8089] = t[8088] ^ n[8089];
assign t[8090] = t[8089] ^ n[8090];
assign t[8091] = t[8090] ^ n[8091];
assign t[8092] = t[8091] ^ n[8092];
assign t[8093] = t[8092] ^ n[8093];
assign t[8094] = t[8093] ^ n[8094];
assign t[8095] = t[8094] ^ n[8095];
assign t[8096] = t[8095] ^ n[8096];
assign t[8097] = t[8096] ^ n[8097];
assign t[8098] = t[8097] ^ n[8098];
assign t[8099] = t[8098] ^ n[8099];
assign t[8100] = t[8099] ^ n[8100];
assign t[8101] = t[8100] ^ n[8101];
assign t[8102] = t[8101] ^ n[8102];
assign t[8103] = t[8102] ^ n[8103];
assign t[8104] = t[8103] ^ n[8104];
assign t[8105] = t[8104] ^ n[8105];
assign t[8106] = t[8105] ^ n[8106];
assign t[8107] = t[8106] ^ n[8107];
assign t[8108] = t[8107] ^ n[8108];
assign t[8109] = t[8108] ^ n[8109];
assign t[8110] = t[8109] ^ n[8110];
assign t[8111] = t[8110] ^ n[8111];
assign t[8112] = t[8111] ^ n[8112];
assign t[8113] = t[8112] ^ n[8113];
assign t[8114] = t[8113] ^ n[8114];
assign t[8115] = t[8114] ^ n[8115];
assign t[8116] = t[8115] ^ n[8116];
assign t[8117] = t[8116] ^ n[8117];
assign t[8118] = t[8117] ^ n[8118];
assign t[8119] = t[8118] ^ n[8119];
assign t[8120] = t[8119] ^ n[8120];
assign t[8121] = t[8120] ^ n[8121];
assign t[8122] = t[8121] ^ n[8122];
assign t[8123] = t[8122] ^ n[8123];
assign t[8124] = t[8123] ^ n[8124];
assign t[8125] = t[8124] ^ n[8125];
assign t[8126] = t[8125] ^ n[8126];
assign t[8127] = t[8126] ^ n[8127];
assign t[8128] = t[8127] ^ n[8128];
assign t[8129] = t[8128] ^ n[8129];
assign t[8130] = t[8129] ^ n[8130];
assign t[8131] = t[8130] ^ n[8131];
assign t[8132] = t[8131] ^ n[8132];
assign t[8133] = t[8132] ^ n[8133];
assign t[8134] = t[8133] ^ n[8134];
assign t[8135] = t[8134] ^ n[8135];
assign t[8136] = t[8135] ^ n[8136];
assign t[8137] = t[8136] ^ n[8137];
assign t[8138] = t[8137] ^ n[8138];
assign t[8139] = t[8138] ^ n[8139];
assign t[8140] = t[8139] ^ n[8140];
assign t[8141] = t[8140] ^ n[8141];
assign t[8142] = t[8141] ^ n[8142];
assign t[8143] = t[8142] ^ n[8143];
assign t[8144] = t[8143] ^ n[8144];
assign t[8145] = t[8144] ^ n[8145];
assign t[8146] = t[8145] ^ n[8146];
assign t[8147] = t[8146] ^ n[8147];
assign t[8148] = t[8147] ^ n[8148];
assign t[8149] = t[8148] ^ n[8149];
assign t[8150] = t[8149] ^ n[8150];
assign t[8151] = t[8150] ^ n[8151];
assign t[8152] = t[8151] ^ n[8152];
assign t[8153] = t[8152] ^ n[8153];
assign t[8154] = t[8153] ^ n[8154];
assign t[8155] = t[8154] ^ n[8155];
assign t[8156] = t[8155] ^ n[8156];
assign t[8157] = t[8156] ^ n[8157];
assign t[8158] = t[8157] ^ n[8158];
assign t[8159] = t[8158] ^ n[8159];
assign t[8160] = t[8159] ^ n[8160];
assign t[8161] = t[8160] ^ n[8161];
assign t[8162] = t[8161] ^ n[8162];
assign t[8163] = t[8162] ^ n[8163];
assign t[8164] = t[8163] ^ n[8164];
assign t[8165] = t[8164] ^ n[8165];
assign t[8166] = t[8165] ^ n[8166];
assign t[8167] = t[8166] ^ n[8167];
assign t[8168] = t[8167] ^ n[8168];
assign t[8169] = t[8168] ^ n[8169];
assign t[8170] = t[8169] ^ n[8170];
assign t[8171] = t[8170] ^ n[8171];
assign t[8172] = t[8171] ^ n[8172];
assign t[8173] = t[8172] ^ n[8173];
assign t[8174] = t[8173] ^ n[8174];
assign t[8175] = t[8174] ^ n[8175];
assign t[8176] = t[8175] ^ n[8176];

assign s[11] = ( a[11] ^ b [11] ) ^ t[8176];

endmodule