
module gen_linear_part ( a, b, c_in, n, s );
  input [6:0] a;
  input [6:0] b;
  input [500:0] n;
  output [7:0] s;
  input c_in;
  wire   t_245, t_244, t_243, t_242, t_241, t_240, t_239, t_238, t_237, t_236,
         t_235, t_234, t_233, t_232, t_231, t_230, t_229, t_228, t_227, t_226,
         t_225, t_224, t_223, t_222, t_221, t_220, t_219, t_218, t_217, t_216,
         t_215, t_214, t_213, t_212, t_211, t_210, t_209, t_208, t_207, t_206,
         t_205, t_204, t_203, t_202, t_201, t_200, t_199, t_198, t_197, t_196,
         t_195, t_194, t_193, t_192, t_191, t_190, t_189, t_188, t_187, t_186,
         t_185, t_184, t_183, t_182, t_181, t_180, t_179, t_178, t_177, t_176,
         t_175, t_174, t_173, t_172, t_171, t_170, t_169, t_168, t_167, t_166,
         t_165, t_164, t_163, t_162, t_161, t_160, t_159, t_158, t_157, t_156,
         t_155, t_154, t_153, t_152, t_151, t_150, t_149, t_148, t_147, t_146,
         t_145, t_144, t_143, t_142, t_141, t_140, t_139, t_138, t_137, t_136,
         t_135, t_134, t_133, t_132, t_131, t_130, t_129, t_128, t_127, t_126,
         t_125, t_124, t_123, t_122, t_121, t_120, t_118, t_117, t_116, t_115,
         t_114, t_113, t_112, t_111, t_110, t_109, t_108, t_107, t_106, t_105,
         t_104, t_103, t_102, t_101, t_100, t_99, t_98, t_97, t_96, t_95, t_94,
         t_93, t_92, t_91, t_90, t_89, t_88, t_87, t_86, t_85, t_84, t_83,
         t_82, t_81, t_80, t_79, t_78, t_77, t_76, t_75, t_74, t_73, t_72,
         t_71, t_70, t_69, t_68, t_67, t_66, t_65, t_64, t_63, t_62, t_61,
         t_60, t_59, t_58, t_57, t_55, t_54, t_53, t_52, t_51, t_50, t_49,
         t_48, t_47, t_46, t_45, t_44, t_43, t_42, t_41, t_40, t_39, t_38,
         t_37, t_36, t_35, t_34, t_33, t_32, t_31, t_30, t_29, t_28, t_27,
         t_26, t_24, t_23, t_22, t_21, t_20, t_19, t_18, t_17, t_16, t_15,
         t_14, t_13, t_12, t_11, t_9, t_8, t_7, t_6, t_5, t_4, t_2, t_1, N0,
         N1, N2, N3, N4, N5, N6;
  wire   [499:247] t;

  CKXOR2D1 C1014 ( .A1(t[499]), .A2(n[500]), .Z(s[7]) );
  CKXOR2D1 C1013 ( .A1(t[498]), .A2(n[499]), .Z(t[499]) );
  CKXOR2D1 C1012 ( .A1(t[497]), .A2(n[498]), .Z(t[498]) );
  CKXOR2D1 C1011 ( .A1(t[496]), .A2(n[497]), .Z(t[497]) );
  CKXOR2D1 C1010 ( .A1(t[495]), .A2(n[496]), .Z(t[496]) );
  CKXOR2D1 C1009 ( .A1(t[494]), .A2(n[495]), .Z(t[495]) );
  CKXOR2D1 C1008 ( .A1(t[493]), .A2(n[494]), .Z(t[494]) );
  CKXOR2D1 C1007 ( .A1(t[492]), .A2(n[493]), .Z(t[493]) );
  CKXOR2D1 C1006 ( .A1(t[491]), .A2(n[492]), .Z(t[492]) );
  CKXOR2D1 C1005 ( .A1(t[490]), .A2(n[491]), .Z(t[491]) );
  CKXOR2D1 C1004 ( .A1(t[489]), .A2(n[490]), .Z(t[490]) );
  CKXOR2D1 C1003 ( .A1(t[488]), .A2(n[489]), .Z(t[489]) );
  CKXOR2D1 C1002 ( .A1(t[487]), .A2(n[488]), .Z(t[488]) );
  CKXOR2D1 C1001 ( .A1(t[486]), .A2(n[487]), .Z(t[487]) );
  CKXOR2D1 C1000 ( .A1(t[485]), .A2(n[486]), .Z(t[486]) );
  CKXOR2D1 C999 ( .A1(t[484]), .A2(n[485]), .Z(t[485]) );
  CKXOR2D1 C998 ( .A1(t[483]), .A2(n[484]), .Z(t[484]) );
  CKXOR2D1 C997 ( .A1(t[482]), .A2(n[483]), .Z(t[483]) );
  CKXOR2D1 C996 ( .A1(t[481]), .A2(n[482]), .Z(t[482]) );
  CKXOR2D1 C995 ( .A1(t[480]), .A2(n[481]), .Z(t[481]) );
  CKXOR2D1 C994 ( .A1(t[479]), .A2(n[480]), .Z(t[480]) );
  CKXOR2D1 C993 ( .A1(t[478]), .A2(n[479]), .Z(t[479]) );
  CKXOR2D1 C992 ( .A1(t[477]), .A2(n[478]), .Z(t[478]) );
  CKXOR2D1 C991 ( .A1(t[476]), .A2(n[477]), .Z(t[477]) );
  CKXOR2D1 C990 ( .A1(t[475]), .A2(n[476]), .Z(t[476]) );
  CKXOR2D1 C989 ( .A1(t[474]), .A2(n[475]), .Z(t[475]) );
  CKXOR2D1 C988 ( .A1(t[473]), .A2(n[474]), .Z(t[474]) );
  CKXOR2D1 C987 ( .A1(t[472]), .A2(n[473]), .Z(t[473]) );
  CKXOR2D1 C986 ( .A1(t[471]), .A2(n[472]), .Z(t[472]) );
  CKXOR2D1 C985 ( .A1(t[470]), .A2(n[471]), .Z(t[471]) );
  CKXOR2D1 C984 ( .A1(t[469]), .A2(n[470]), .Z(t[470]) );
  CKXOR2D1 C983 ( .A1(t[468]), .A2(n[469]), .Z(t[469]) );
  CKXOR2D1 C982 ( .A1(t[467]), .A2(n[468]), .Z(t[468]) );
  CKXOR2D1 C981 ( .A1(t[466]), .A2(n[467]), .Z(t[467]) );
  CKXOR2D1 C980 ( .A1(t[465]), .A2(n[466]), .Z(t[466]) );
  CKXOR2D1 C979 ( .A1(t[464]), .A2(n[465]), .Z(t[465]) );
  CKXOR2D1 C978 ( .A1(t[463]), .A2(n[464]), .Z(t[464]) );
  CKXOR2D1 C977 ( .A1(t[462]), .A2(n[463]), .Z(t[463]) );
  CKXOR2D1 C976 ( .A1(t[461]), .A2(n[462]), .Z(t[462]) );
  CKXOR2D1 C975 ( .A1(t[460]), .A2(n[461]), .Z(t[461]) );
  CKXOR2D1 C974 ( .A1(t[459]), .A2(n[460]), .Z(t[460]) );
  CKXOR2D1 C973 ( .A1(t[458]), .A2(n[459]), .Z(t[459]) );
  CKXOR2D1 C972 ( .A1(t[457]), .A2(n[458]), .Z(t[458]) );
  CKXOR2D1 C971 ( .A1(t[456]), .A2(n[457]), .Z(t[457]) );
  CKXOR2D1 C970 ( .A1(t[455]), .A2(n[456]), .Z(t[456]) );
  CKXOR2D1 C969 ( .A1(t[454]), .A2(n[455]), .Z(t[455]) );
  CKXOR2D1 C968 ( .A1(t[453]), .A2(n[454]), .Z(t[454]) );
  CKXOR2D1 C967 ( .A1(t[452]), .A2(n[453]), .Z(t[453]) );
  CKXOR2D1 C966 ( .A1(t[451]), .A2(n[452]), .Z(t[452]) );
  CKXOR2D1 C965 ( .A1(t[450]), .A2(n[451]), .Z(t[451]) );
  CKXOR2D1 C964 ( .A1(t[449]), .A2(n[450]), .Z(t[450]) );
  CKXOR2D1 C963 ( .A1(t[448]), .A2(n[449]), .Z(t[449]) );
  CKXOR2D1 C962 ( .A1(t[447]), .A2(n[448]), .Z(t[448]) );
  CKXOR2D1 C961 ( .A1(t[446]), .A2(n[447]), .Z(t[447]) );
  CKXOR2D1 C960 ( .A1(t[445]), .A2(n[446]), .Z(t[446]) );
  CKXOR2D1 C959 ( .A1(t[444]), .A2(n[445]), .Z(t[445]) );
  CKXOR2D1 C958 ( .A1(t[443]), .A2(n[444]), .Z(t[444]) );
  CKXOR2D1 C957 ( .A1(t[442]), .A2(n[443]), .Z(t[443]) );
  CKXOR2D1 C956 ( .A1(t[441]), .A2(n[442]), .Z(t[442]) );
  CKXOR2D1 C955 ( .A1(t[440]), .A2(n[441]), .Z(t[441]) );
  CKXOR2D1 C954 ( .A1(t[439]), .A2(n[440]), .Z(t[440]) );
  CKXOR2D1 C953 ( .A1(t[438]), .A2(n[439]), .Z(t[439]) );
  CKXOR2D1 C952 ( .A1(t[437]), .A2(n[438]), .Z(t[438]) );
  CKXOR2D1 C951 ( .A1(t[436]), .A2(n[437]), .Z(t[437]) );
  CKXOR2D1 C950 ( .A1(t[435]), .A2(n[436]), .Z(t[436]) );
  CKXOR2D1 C949 ( .A1(t[434]), .A2(n[435]), .Z(t[435]) );
  CKXOR2D1 C948 ( .A1(t[433]), .A2(n[434]), .Z(t[434]) );
  CKXOR2D1 C947 ( .A1(t[432]), .A2(n[433]), .Z(t[433]) );
  CKXOR2D1 C946 ( .A1(t[431]), .A2(n[432]), .Z(t[432]) );
  CKXOR2D1 C945 ( .A1(t[430]), .A2(n[431]), .Z(t[431]) );
  CKXOR2D1 C944 ( .A1(t[429]), .A2(n[430]), .Z(t[430]) );
  CKXOR2D1 C943 ( .A1(t[428]), .A2(n[429]), .Z(t[429]) );
  CKXOR2D1 C942 ( .A1(t[427]), .A2(n[428]), .Z(t[428]) );
  CKXOR2D1 C941 ( .A1(t[426]), .A2(n[427]), .Z(t[427]) );
  CKXOR2D1 C940 ( .A1(t[425]), .A2(n[426]), .Z(t[426]) );
  CKXOR2D1 C939 ( .A1(t[424]), .A2(n[425]), .Z(t[425]) );
  CKXOR2D1 C938 ( .A1(t[423]), .A2(n[424]), .Z(t[424]) );
  CKXOR2D1 C937 ( .A1(t[422]), .A2(n[423]), .Z(t[423]) );
  CKXOR2D1 C936 ( .A1(t[421]), .A2(n[422]), .Z(t[422]) );
  CKXOR2D1 C935 ( .A1(t[420]), .A2(n[421]), .Z(t[421]) );
  CKXOR2D1 C934 ( .A1(t[419]), .A2(n[420]), .Z(t[420]) );
  CKXOR2D1 C933 ( .A1(t[418]), .A2(n[419]), .Z(t[419]) );
  CKXOR2D1 C932 ( .A1(t[417]), .A2(n[418]), .Z(t[418]) );
  CKXOR2D1 C931 ( .A1(t[416]), .A2(n[417]), .Z(t[417]) );
  CKXOR2D1 C930 ( .A1(t[415]), .A2(n[416]), .Z(t[416]) );
  CKXOR2D1 C929 ( .A1(t[414]), .A2(n[415]), .Z(t[415]) );
  CKXOR2D1 C928 ( .A1(t[413]), .A2(n[414]), .Z(t[414]) );
  CKXOR2D1 C927 ( .A1(t[412]), .A2(n[413]), .Z(t[413]) );
  CKXOR2D1 C926 ( .A1(t[411]), .A2(n[412]), .Z(t[412]) );
  CKXOR2D1 C925 ( .A1(t[410]), .A2(n[411]), .Z(t[411]) );
  CKXOR2D1 C924 ( .A1(t[409]), .A2(n[410]), .Z(t[410]) );
  CKXOR2D1 C923 ( .A1(t[408]), .A2(n[409]), .Z(t[409]) );
  CKXOR2D1 C922 ( .A1(t[407]), .A2(n[408]), .Z(t[408]) );
  CKXOR2D1 C921 ( .A1(t[406]), .A2(n[407]), .Z(t[407]) );
  CKXOR2D1 C920 ( .A1(t[405]), .A2(n[406]), .Z(t[406]) );
  CKXOR2D1 C919 ( .A1(t[404]), .A2(n[405]), .Z(t[405]) );
  CKXOR2D1 C918 ( .A1(t[403]), .A2(n[404]), .Z(t[404]) );
  CKXOR2D1 C917 ( .A1(t[402]), .A2(n[403]), .Z(t[403]) );
  CKXOR2D1 C916 ( .A1(t[401]), .A2(n[402]), .Z(t[402]) );
  CKXOR2D1 C915 ( .A1(t[400]), .A2(n[401]), .Z(t[401]) );
  CKXOR2D1 C914 ( .A1(t[399]), .A2(n[400]), .Z(t[400]) );
  CKXOR2D1 C913 ( .A1(t[398]), .A2(n[399]), .Z(t[399]) );
  CKXOR2D1 C912 ( .A1(t[397]), .A2(n[398]), .Z(t[398]) );
  CKXOR2D1 C911 ( .A1(t[396]), .A2(n[397]), .Z(t[397]) );
  CKXOR2D1 C910 ( .A1(t[395]), .A2(n[396]), .Z(t[396]) );
  CKXOR2D1 C909 ( .A1(t[394]), .A2(n[395]), .Z(t[395]) );
  CKXOR2D1 C908 ( .A1(t[393]), .A2(n[394]), .Z(t[394]) );
  CKXOR2D1 C907 ( .A1(t[392]), .A2(n[393]), .Z(t[393]) );
  CKXOR2D1 C906 ( .A1(t[391]), .A2(n[392]), .Z(t[392]) );
  CKXOR2D1 C905 ( .A1(t[390]), .A2(n[391]), .Z(t[391]) );
  CKXOR2D1 C904 ( .A1(t[389]), .A2(n[390]), .Z(t[390]) );
  CKXOR2D1 C903 ( .A1(t[388]), .A2(n[389]), .Z(t[389]) );
  CKXOR2D1 C902 ( .A1(t[387]), .A2(n[388]), .Z(t[388]) );
  CKXOR2D1 C901 ( .A1(t[386]), .A2(n[387]), .Z(t[387]) );
  CKXOR2D1 C900 ( .A1(t[385]), .A2(n[386]), .Z(t[386]) );
  CKXOR2D1 C899 ( .A1(t[384]), .A2(n[385]), .Z(t[385]) );
  CKXOR2D1 C898 ( .A1(t[383]), .A2(n[384]), .Z(t[384]) );
  CKXOR2D1 C897 ( .A1(t[382]), .A2(n[383]), .Z(t[383]) );
  CKXOR2D1 C896 ( .A1(t[381]), .A2(n[382]), .Z(t[382]) );
  CKXOR2D1 C895 ( .A1(t[380]), .A2(n[381]), .Z(t[381]) );
  CKXOR2D1 C894 ( .A1(t[379]), .A2(n[380]), .Z(t[380]) );
  CKXOR2D1 C893 ( .A1(t[378]), .A2(n[379]), .Z(t[379]) );
  CKXOR2D1 C892 ( .A1(t[377]), .A2(n[378]), .Z(t[378]) );
  CKXOR2D1 C891 ( .A1(t[376]), .A2(n[377]), .Z(t[377]) );
  CKXOR2D1 C890 ( .A1(t[375]), .A2(n[376]), .Z(t[376]) );
  CKXOR2D1 C889 ( .A1(t[374]), .A2(n[375]), .Z(t[375]) );
  CKXOR2D1 C888 ( .A1(t[373]), .A2(n[374]), .Z(t[374]) );
  CKXOR2D1 C887 ( .A1(t[372]), .A2(n[373]), .Z(t[373]) );
  CKXOR2D1 C886 ( .A1(t[371]), .A2(n[372]), .Z(t[372]) );
  CKXOR2D1 C885 ( .A1(t[370]), .A2(n[371]), .Z(t[371]) );
  CKXOR2D1 C884 ( .A1(t[369]), .A2(n[370]), .Z(t[370]) );
  CKXOR2D1 C883 ( .A1(t[368]), .A2(n[369]), .Z(t[369]) );
  CKXOR2D1 C882 ( .A1(t[367]), .A2(n[368]), .Z(t[368]) );
  CKXOR2D1 C881 ( .A1(t[366]), .A2(n[367]), .Z(t[367]) );
  CKXOR2D1 C880 ( .A1(t[365]), .A2(n[366]), .Z(t[366]) );
  CKXOR2D1 C879 ( .A1(t[364]), .A2(n[365]), .Z(t[365]) );
  CKXOR2D1 C878 ( .A1(t[363]), .A2(n[364]), .Z(t[364]) );
  CKXOR2D1 C877 ( .A1(t[362]), .A2(n[363]), .Z(t[363]) );
  CKXOR2D1 C876 ( .A1(t[361]), .A2(n[362]), .Z(t[362]) );
  CKXOR2D1 C875 ( .A1(t[360]), .A2(n[361]), .Z(t[361]) );
  CKXOR2D1 C874 ( .A1(t[359]), .A2(n[360]), .Z(t[360]) );
  CKXOR2D1 C873 ( .A1(t[358]), .A2(n[359]), .Z(t[359]) );
  CKXOR2D1 C872 ( .A1(t[357]), .A2(n[358]), .Z(t[358]) );
  CKXOR2D1 C871 ( .A1(t[356]), .A2(n[357]), .Z(t[357]) );
  CKXOR2D1 C870 ( .A1(t[355]), .A2(n[356]), .Z(t[356]) );
  CKXOR2D1 C869 ( .A1(t[354]), .A2(n[355]), .Z(t[355]) );
  CKXOR2D1 C868 ( .A1(t[353]), .A2(n[354]), .Z(t[354]) );
  CKXOR2D1 C867 ( .A1(t[352]), .A2(n[353]), .Z(t[353]) );
  CKXOR2D1 C866 ( .A1(t[351]), .A2(n[352]), .Z(t[352]) );
  CKXOR2D1 C865 ( .A1(t[350]), .A2(n[351]), .Z(t[351]) );
  CKXOR2D1 C864 ( .A1(t[349]), .A2(n[350]), .Z(t[350]) );
  CKXOR2D1 C863 ( .A1(t[348]), .A2(n[349]), .Z(t[349]) );
  CKXOR2D1 C862 ( .A1(t[347]), .A2(n[348]), .Z(t[348]) );
  CKXOR2D1 C861 ( .A1(t[346]), .A2(n[347]), .Z(t[347]) );
  CKXOR2D1 C860 ( .A1(t[345]), .A2(n[346]), .Z(t[346]) );
  CKXOR2D1 C859 ( .A1(t[344]), .A2(n[345]), .Z(t[345]) );
  CKXOR2D1 C858 ( .A1(t[343]), .A2(n[344]), .Z(t[344]) );
  CKXOR2D1 C857 ( .A1(t[342]), .A2(n[343]), .Z(t[343]) );
  CKXOR2D1 C856 ( .A1(t[341]), .A2(n[342]), .Z(t[342]) );
  CKXOR2D1 C855 ( .A1(t[340]), .A2(n[341]), .Z(t[341]) );
  CKXOR2D1 C854 ( .A1(t[339]), .A2(n[340]), .Z(t[340]) );
  CKXOR2D1 C853 ( .A1(t[338]), .A2(n[339]), .Z(t[339]) );
  CKXOR2D1 C852 ( .A1(t[337]), .A2(n[338]), .Z(t[338]) );
  CKXOR2D1 C851 ( .A1(t[336]), .A2(n[337]), .Z(t[337]) );
  CKXOR2D1 C850 ( .A1(t[335]), .A2(n[336]), .Z(t[336]) );
  CKXOR2D1 C849 ( .A1(t[334]), .A2(n[335]), .Z(t[335]) );
  CKXOR2D1 C848 ( .A1(t[333]), .A2(n[334]), .Z(t[334]) );
  CKXOR2D1 C847 ( .A1(t[332]), .A2(n[333]), .Z(t[333]) );
  CKXOR2D1 C846 ( .A1(t[331]), .A2(n[332]), .Z(t[332]) );
  CKXOR2D1 C845 ( .A1(t[330]), .A2(n[331]), .Z(t[331]) );
  CKXOR2D1 C844 ( .A1(t[329]), .A2(n[330]), .Z(t[330]) );
  CKXOR2D1 C843 ( .A1(t[328]), .A2(n[329]), .Z(t[329]) );
  CKXOR2D1 C842 ( .A1(t[327]), .A2(n[328]), .Z(t[328]) );
  CKXOR2D1 C841 ( .A1(t[326]), .A2(n[327]), .Z(t[327]) );
  CKXOR2D1 C840 ( .A1(t[325]), .A2(n[326]), .Z(t[326]) );
  CKXOR2D1 C839 ( .A1(t[324]), .A2(n[325]), .Z(t[325]) );
  CKXOR2D1 C838 ( .A1(t[323]), .A2(n[324]), .Z(t[324]) );
  CKXOR2D1 C837 ( .A1(t[322]), .A2(n[323]), .Z(t[323]) );
  CKXOR2D1 C836 ( .A1(t[321]), .A2(n[322]), .Z(t[322]) );
  CKXOR2D1 C835 ( .A1(t[320]), .A2(n[321]), .Z(t[321]) );
  CKXOR2D1 C834 ( .A1(t[319]), .A2(n[320]), .Z(t[320]) );
  CKXOR2D1 C833 ( .A1(t[318]), .A2(n[319]), .Z(t[319]) );
  CKXOR2D1 C832 ( .A1(t[317]), .A2(n[318]), .Z(t[318]) );
  CKXOR2D1 C831 ( .A1(t[316]), .A2(n[317]), .Z(t[317]) );
  CKXOR2D1 C830 ( .A1(t[315]), .A2(n[316]), .Z(t[316]) );
  CKXOR2D1 C829 ( .A1(t[314]), .A2(n[315]), .Z(t[315]) );
  CKXOR2D1 C828 ( .A1(t[313]), .A2(n[314]), .Z(t[314]) );
  CKXOR2D1 C827 ( .A1(t[312]), .A2(n[313]), .Z(t[313]) );
  CKXOR2D1 C826 ( .A1(t[311]), .A2(n[312]), .Z(t[312]) );
  CKXOR2D1 C825 ( .A1(t[310]), .A2(n[311]), .Z(t[311]) );
  CKXOR2D1 C824 ( .A1(t[309]), .A2(n[310]), .Z(t[310]) );
  CKXOR2D1 C823 ( .A1(t[308]), .A2(n[309]), .Z(t[309]) );
  CKXOR2D1 C822 ( .A1(t[307]), .A2(n[308]), .Z(t[308]) );
  CKXOR2D1 C821 ( .A1(t[306]), .A2(n[307]), .Z(t[307]) );
  CKXOR2D1 C820 ( .A1(t[305]), .A2(n[306]), .Z(t[306]) );
  CKXOR2D1 C819 ( .A1(t[304]), .A2(n[305]), .Z(t[305]) );
  CKXOR2D1 C818 ( .A1(t[303]), .A2(n[304]), .Z(t[304]) );
  CKXOR2D1 C817 ( .A1(t[302]), .A2(n[303]), .Z(t[303]) );
  CKXOR2D1 C816 ( .A1(t[301]), .A2(n[302]), .Z(t[302]) );
  CKXOR2D1 C815 ( .A1(t[300]), .A2(n[301]), .Z(t[301]) );
  CKXOR2D1 C814 ( .A1(t[299]), .A2(n[300]), .Z(t[300]) );
  CKXOR2D1 C813 ( .A1(t[298]), .A2(n[299]), .Z(t[299]) );
  CKXOR2D1 C812 ( .A1(t[297]), .A2(n[298]), .Z(t[298]) );
  CKXOR2D1 C811 ( .A1(t[296]), .A2(n[297]), .Z(t[297]) );
  CKXOR2D1 C810 ( .A1(t[295]), .A2(n[296]), .Z(t[296]) );
  CKXOR2D1 C809 ( .A1(t[294]), .A2(n[295]), .Z(t[295]) );
  CKXOR2D1 C808 ( .A1(t[293]), .A2(n[294]), .Z(t[294]) );
  CKXOR2D1 C807 ( .A1(t[292]), .A2(n[293]), .Z(t[293]) );
  CKXOR2D1 C806 ( .A1(t[291]), .A2(n[292]), .Z(t[292]) );
  CKXOR2D1 C805 ( .A1(t[290]), .A2(n[291]), .Z(t[291]) );
  CKXOR2D1 C804 ( .A1(t[289]), .A2(n[290]), .Z(t[290]) );
  CKXOR2D1 C803 ( .A1(t[288]), .A2(n[289]), .Z(t[289]) );
  CKXOR2D1 C802 ( .A1(t[287]), .A2(n[288]), .Z(t[288]) );
  CKXOR2D1 C801 ( .A1(t[286]), .A2(n[287]), .Z(t[287]) );
  CKXOR2D1 C800 ( .A1(t[285]), .A2(n[286]), .Z(t[286]) );
  CKXOR2D1 C799 ( .A1(t[284]), .A2(n[285]), .Z(t[285]) );
  CKXOR2D1 C798 ( .A1(t[283]), .A2(n[284]), .Z(t[284]) );
  CKXOR2D1 C797 ( .A1(t[282]), .A2(n[283]), .Z(t[283]) );
  CKXOR2D1 C796 ( .A1(t[281]), .A2(n[282]), .Z(t[282]) );
  CKXOR2D1 C795 ( .A1(t[280]), .A2(n[281]), .Z(t[281]) );
  CKXOR2D1 C794 ( .A1(t[279]), .A2(n[280]), .Z(t[280]) );
  CKXOR2D1 C793 ( .A1(t[278]), .A2(n[279]), .Z(t[279]) );
  CKXOR2D1 C792 ( .A1(t[277]), .A2(n[278]), .Z(t[278]) );
  CKXOR2D1 C791 ( .A1(t[276]), .A2(n[277]), .Z(t[277]) );
  CKXOR2D1 C790 ( .A1(t[275]), .A2(n[276]), .Z(t[276]) );
  CKXOR2D1 C789 ( .A1(t[274]), .A2(n[275]), .Z(t[275]) );
  CKXOR2D1 C788 ( .A1(t[273]), .A2(n[274]), .Z(t[274]) );
  CKXOR2D1 C787 ( .A1(t[272]), .A2(n[273]), .Z(t[273]) );
  CKXOR2D1 C786 ( .A1(t[271]), .A2(n[272]), .Z(t[272]) );
  CKXOR2D1 C785 ( .A1(t[270]), .A2(n[271]), .Z(t[271]) );
  CKXOR2D1 C784 ( .A1(t[269]), .A2(n[270]), .Z(t[270]) );
  CKXOR2D1 C783 ( .A1(t[268]), .A2(n[269]), .Z(t[269]) );
  CKXOR2D1 C782 ( .A1(t[267]), .A2(n[268]), .Z(t[268]) );
  CKXOR2D1 C781 ( .A1(t[266]), .A2(n[267]), .Z(t[267]) );
  CKXOR2D1 C780 ( .A1(t[265]), .A2(n[266]), .Z(t[266]) );
  CKXOR2D1 C779 ( .A1(t[264]), .A2(n[265]), .Z(t[265]) );
  CKXOR2D1 C778 ( .A1(t[263]), .A2(n[264]), .Z(t[264]) );
  CKXOR2D1 C777 ( .A1(t[262]), .A2(n[263]), .Z(t[263]) );
  CKXOR2D1 C776 ( .A1(t[261]), .A2(n[262]), .Z(t[262]) );
  CKXOR2D1 C775 ( .A1(t[260]), .A2(n[261]), .Z(t[261]) );
  CKXOR2D1 C774 ( .A1(t[259]), .A2(n[260]), .Z(t[260]) );
  CKXOR2D1 C773 ( .A1(t[258]), .A2(n[259]), .Z(t[259]) );
  CKXOR2D1 C772 ( .A1(t[257]), .A2(n[258]), .Z(t[258]) );
  CKXOR2D1 C771 ( .A1(t[256]), .A2(n[257]), .Z(t[257]) );
  CKXOR2D1 C770 ( .A1(t[255]), .A2(n[256]), .Z(t[256]) );
  CKXOR2D1 C769 ( .A1(t[254]), .A2(n[255]), .Z(t[255]) );
  CKXOR2D1 C768 ( .A1(t[253]), .A2(n[254]), .Z(t[254]) );
  CKXOR2D1 C767 ( .A1(t[252]), .A2(n[253]), .Z(t[253]) );
  CKXOR2D1 C766 ( .A1(t[251]), .A2(n[252]), .Z(t[252]) );
  CKXOR2D1 C765 ( .A1(t[250]), .A2(n[251]), .Z(t[251]) );
  CKXOR2D1 C764 ( .A1(t[249]), .A2(n[250]), .Z(t[250]) );
  CKXOR2D1 C763 ( .A1(t[248]), .A2(n[249]), .Z(t[249]) );
  CKXOR2D1 C762 ( .A1(t[247]), .A2(n[248]), .Z(t[248]) );
  CKXOR2D1 C761 ( .A1(n[246]), .A2(n[247]), .Z(t[247]) );
  CKXOR2D1 C760 ( .A1(a[6]), .A2(b[6]), .Z(N6) );
  CKXOR2D1 C759 ( .A1(N6), .A2(t_245), .Z(s[6]) );
  CKXOR2D1 C758 ( .A1(t_244), .A2(n[245]), .Z(t_245) );
  CKXOR2D1 C757 ( .A1(t_243), .A2(n[244]), .Z(t_244) );
  CKXOR2D1 C756 ( .A1(t_242), .A2(n[243]), .Z(t_243) );
  CKXOR2D1 C755 ( .A1(t_241), .A2(n[242]), .Z(t_242) );
  CKXOR2D1 C754 ( .A1(t_240), .A2(n[241]), .Z(t_241) );
  CKXOR2D1 C753 ( .A1(t_239), .A2(n[240]), .Z(t_240) );
  CKXOR2D1 C752 ( .A1(t_238), .A2(n[239]), .Z(t_239) );
  CKXOR2D1 C751 ( .A1(t_237), .A2(n[238]), .Z(t_238) );
  CKXOR2D1 C750 ( .A1(t_236), .A2(n[237]), .Z(t_237) );
  CKXOR2D1 C749 ( .A1(t_235), .A2(n[236]), .Z(t_236) );
  CKXOR2D1 C748 ( .A1(t_234), .A2(n[235]), .Z(t_235) );
  CKXOR2D1 C747 ( .A1(t_233), .A2(n[234]), .Z(t_234) );
  CKXOR2D1 C746 ( .A1(t_232), .A2(n[233]), .Z(t_233) );
  CKXOR2D1 C745 ( .A1(t_231), .A2(n[232]), .Z(t_232) );
  CKXOR2D1 C744 ( .A1(t_230), .A2(n[231]), .Z(t_231) );
  CKXOR2D1 C743 ( .A1(t_229), .A2(n[230]), .Z(t_230) );
  CKXOR2D1 C742 ( .A1(t_228), .A2(n[229]), .Z(t_229) );
  CKXOR2D1 C741 ( .A1(t_227), .A2(n[228]), .Z(t_228) );
  CKXOR2D1 C740 ( .A1(t_226), .A2(n[227]), .Z(t_227) );
  CKXOR2D1 C739 ( .A1(t_225), .A2(n[226]), .Z(t_226) );
  CKXOR2D1 C738 ( .A1(t_224), .A2(n[225]), .Z(t_225) );
  CKXOR2D1 C737 ( .A1(t_223), .A2(n[224]), .Z(t_224) );
  CKXOR2D1 C736 ( .A1(t_222), .A2(n[223]), .Z(t_223) );
  CKXOR2D1 C735 ( .A1(t_221), .A2(n[222]), .Z(t_222) );
  CKXOR2D1 C734 ( .A1(t_220), .A2(n[221]), .Z(t_221) );
  CKXOR2D1 C733 ( .A1(t_219), .A2(n[220]), .Z(t_220) );
  CKXOR2D1 C732 ( .A1(t_218), .A2(n[219]), .Z(t_219) );
  CKXOR2D1 C731 ( .A1(t_217), .A2(n[218]), .Z(t_218) );
  CKXOR2D1 C730 ( .A1(t_216), .A2(n[217]), .Z(t_217) );
  CKXOR2D1 C729 ( .A1(t_215), .A2(n[216]), .Z(t_216) );
  CKXOR2D1 C728 ( .A1(t_214), .A2(n[215]), .Z(t_215) );
  CKXOR2D1 C727 ( .A1(t_213), .A2(n[214]), .Z(t_214) );
  CKXOR2D1 C726 ( .A1(t_212), .A2(n[213]), .Z(t_213) );
  CKXOR2D1 C725 ( .A1(t_211), .A2(n[212]), .Z(t_212) );
  CKXOR2D1 C724 ( .A1(t_210), .A2(n[211]), .Z(t_211) );
  CKXOR2D1 C723 ( .A1(t_209), .A2(n[210]), .Z(t_210) );
  CKXOR2D1 C722 ( .A1(t_208), .A2(n[209]), .Z(t_209) );
  CKXOR2D1 C721 ( .A1(t_207), .A2(n[208]), .Z(t_208) );
  CKXOR2D1 C720 ( .A1(t_206), .A2(n[207]), .Z(t_207) );
  CKXOR2D1 C719 ( .A1(t_205), .A2(n[206]), .Z(t_206) );
  CKXOR2D1 C718 ( .A1(t_204), .A2(n[205]), .Z(t_205) );
  CKXOR2D1 C717 ( .A1(t_203), .A2(n[204]), .Z(t_204) );
  CKXOR2D1 C716 ( .A1(t_202), .A2(n[203]), .Z(t_203) );
  CKXOR2D1 C715 ( .A1(t_201), .A2(n[202]), .Z(t_202) );
  CKXOR2D1 C714 ( .A1(t_200), .A2(n[201]), .Z(t_201) );
  CKXOR2D1 C713 ( .A1(t_199), .A2(n[200]), .Z(t_200) );
  CKXOR2D1 C712 ( .A1(t_198), .A2(n[199]), .Z(t_199) );
  CKXOR2D1 C711 ( .A1(t_197), .A2(n[198]), .Z(t_198) );
  CKXOR2D1 C710 ( .A1(t_196), .A2(n[197]), .Z(t_197) );
  CKXOR2D1 C709 ( .A1(t_195), .A2(n[196]), .Z(t_196) );
  CKXOR2D1 C708 ( .A1(t_194), .A2(n[195]), .Z(t_195) );
  CKXOR2D1 C707 ( .A1(t_193), .A2(n[194]), .Z(t_194) );
  CKXOR2D1 C706 ( .A1(t_192), .A2(n[193]), .Z(t_193) );
  CKXOR2D1 C705 ( .A1(t_191), .A2(n[192]), .Z(t_192) );
  CKXOR2D1 C704 ( .A1(t_190), .A2(n[191]), .Z(t_191) );
  CKXOR2D1 C703 ( .A1(t_189), .A2(n[190]), .Z(t_190) );
  CKXOR2D1 C702 ( .A1(t_188), .A2(n[189]), .Z(t_189) );
  CKXOR2D1 C701 ( .A1(t_187), .A2(n[188]), .Z(t_188) );
  CKXOR2D1 C700 ( .A1(t_186), .A2(n[187]), .Z(t_187) );
  CKXOR2D1 C699 ( .A1(t_185), .A2(n[186]), .Z(t_186) );
  CKXOR2D1 C698 ( .A1(t_184), .A2(n[185]), .Z(t_185) );
  CKXOR2D1 C697 ( .A1(t_183), .A2(n[184]), .Z(t_184) );
  CKXOR2D1 C696 ( .A1(t_182), .A2(n[183]), .Z(t_183) );
  CKXOR2D1 C695 ( .A1(t_181), .A2(n[182]), .Z(t_182) );
  CKXOR2D1 C694 ( .A1(t_180), .A2(n[181]), .Z(t_181) );
  CKXOR2D1 C693 ( .A1(t_179), .A2(n[180]), .Z(t_180) );
  CKXOR2D1 C692 ( .A1(t_178), .A2(n[179]), .Z(t_179) );
  CKXOR2D1 C691 ( .A1(t_177), .A2(n[178]), .Z(t_178) );
  CKXOR2D1 C690 ( .A1(t_176), .A2(n[177]), .Z(t_177) );
  CKXOR2D1 C689 ( .A1(t_175), .A2(n[176]), .Z(t_176) );
  CKXOR2D1 C688 ( .A1(t_174), .A2(n[175]), .Z(t_175) );
  CKXOR2D1 C687 ( .A1(t_173), .A2(n[174]), .Z(t_174) );
  CKXOR2D1 C686 ( .A1(t_172), .A2(n[173]), .Z(t_173) );
  CKXOR2D1 C685 ( .A1(t_171), .A2(n[172]), .Z(t_172) );
  CKXOR2D1 C684 ( .A1(t_170), .A2(n[171]), .Z(t_171) );
  CKXOR2D1 C683 ( .A1(t_169), .A2(n[170]), .Z(t_170) );
  CKXOR2D1 C682 ( .A1(t_168), .A2(n[169]), .Z(t_169) );
  CKXOR2D1 C681 ( .A1(t_167), .A2(n[168]), .Z(t_168) );
  CKXOR2D1 C680 ( .A1(t_166), .A2(n[167]), .Z(t_167) );
  CKXOR2D1 C679 ( .A1(t_165), .A2(n[166]), .Z(t_166) );
  CKXOR2D1 C678 ( .A1(t_164), .A2(n[165]), .Z(t_165) );
  CKXOR2D1 C677 ( .A1(t_163), .A2(n[164]), .Z(t_164) );
  CKXOR2D1 C676 ( .A1(t_162), .A2(n[163]), .Z(t_163) );
  CKXOR2D1 C675 ( .A1(t_161), .A2(n[162]), .Z(t_162) );
  CKXOR2D1 C674 ( .A1(t_160), .A2(n[161]), .Z(t_161) );
  CKXOR2D1 C673 ( .A1(t_159), .A2(n[160]), .Z(t_160) );
  CKXOR2D1 C672 ( .A1(t_158), .A2(n[159]), .Z(t_159) );
  CKXOR2D1 C671 ( .A1(t_157), .A2(n[158]), .Z(t_158) );
  CKXOR2D1 C670 ( .A1(t_156), .A2(n[157]), .Z(t_157) );
  CKXOR2D1 C669 ( .A1(t_155), .A2(n[156]), .Z(t_156) );
  CKXOR2D1 C668 ( .A1(t_154), .A2(n[155]), .Z(t_155) );
  CKXOR2D1 C667 ( .A1(t_153), .A2(n[154]), .Z(t_154) );
  CKXOR2D1 C666 ( .A1(t_152), .A2(n[153]), .Z(t_153) );
  CKXOR2D1 C665 ( .A1(t_151), .A2(n[152]), .Z(t_152) );
  CKXOR2D1 C664 ( .A1(t_150), .A2(n[151]), .Z(t_151) );
  CKXOR2D1 C663 ( .A1(t_149), .A2(n[150]), .Z(t_150) );
  CKXOR2D1 C662 ( .A1(t_148), .A2(n[149]), .Z(t_149) );
  CKXOR2D1 C661 ( .A1(t_147), .A2(n[148]), .Z(t_148) );
  CKXOR2D1 C660 ( .A1(t_146), .A2(n[147]), .Z(t_147) );
  CKXOR2D1 C659 ( .A1(t_145), .A2(n[146]), .Z(t_146) );
  CKXOR2D1 C658 ( .A1(t_144), .A2(n[145]), .Z(t_145) );
  CKXOR2D1 C657 ( .A1(t_143), .A2(n[144]), .Z(t_144) );
  CKXOR2D1 C656 ( .A1(t_142), .A2(n[143]), .Z(t_143) );
  CKXOR2D1 C655 ( .A1(t_141), .A2(n[142]), .Z(t_142) );
  CKXOR2D1 C654 ( .A1(t_140), .A2(n[141]), .Z(t_141) );
  CKXOR2D1 C653 ( .A1(t_139), .A2(n[140]), .Z(t_140) );
  CKXOR2D1 C652 ( .A1(t_138), .A2(n[139]), .Z(t_139) );
  CKXOR2D1 C651 ( .A1(t_137), .A2(n[138]), .Z(t_138) );
  CKXOR2D1 C650 ( .A1(t_136), .A2(n[137]), .Z(t_137) );
  CKXOR2D1 C649 ( .A1(t_135), .A2(n[136]), .Z(t_136) );
  CKXOR2D1 C648 ( .A1(t_134), .A2(n[135]), .Z(t_135) );
  CKXOR2D1 C647 ( .A1(t_133), .A2(n[134]), .Z(t_134) );
  CKXOR2D1 C646 ( .A1(t_132), .A2(n[133]), .Z(t_133) );
  CKXOR2D1 C645 ( .A1(t_131), .A2(n[132]), .Z(t_132) );
  CKXOR2D1 C644 ( .A1(t_130), .A2(n[131]), .Z(t_131) );
  CKXOR2D1 C643 ( .A1(t_129), .A2(n[130]), .Z(t_130) );
  CKXOR2D1 C642 ( .A1(t_128), .A2(n[129]), .Z(t_129) );
  CKXOR2D1 C641 ( .A1(t_127), .A2(n[128]), .Z(t_128) );
  CKXOR2D1 C640 ( .A1(t_126), .A2(n[127]), .Z(t_127) );
  CKXOR2D1 C639 ( .A1(t_125), .A2(n[126]), .Z(t_126) );
  CKXOR2D1 C638 ( .A1(t_124), .A2(n[125]), .Z(t_125) );
  CKXOR2D1 C637 ( .A1(t_123), .A2(n[124]), .Z(t_124) );
  CKXOR2D1 C636 ( .A1(t_122), .A2(n[123]), .Z(t_123) );
  CKXOR2D1 C635 ( .A1(t_121), .A2(n[122]), .Z(t_122) );
  CKXOR2D1 C634 ( .A1(t_120), .A2(n[121]), .Z(t_121) );
  CKXOR2D1 C633 ( .A1(n[119]), .A2(n[120]), .Z(t_120) );
  CKXOR2D1 C632 ( .A1(a[5]), .A2(b[5]), .Z(N5) );
  CKXOR2D1 C631 ( .A1(N5), .A2(t_118), .Z(s[5]) );
  CKXOR2D1 C630 ( .A1(t_117), .A2(n[118]), .Z(t_118) );
  CKXOR2D1 C629 ( .A1(t_116), .A2(n[117]), .Z(t_117) );
  CKXOR2D1 C628 ( .A1(t_115), .A2(n[116]), .Z(t_116) );
  CKXOR2D1 C627 ( .A1(t_114), .A2(n[115]), .Z(t_115) );
  CKXOR2D1 C626 ( .A1(t_113), .A2(n[114]), .Z(t_114) );
  CKXOR2D1 C625 ( .A1(t_112), .A2(n[113]), .Z(t_113) );
  CKXOR2D1 C624 ( .A1(t_111), .A2(n[112]), .Z(t_112) );
  CKXOR2D1 C623 ( .A1(t_110), .A2(n[111]), .Z(t_111) );
  CKXOR2D1 C622 ( .A1(t_109), .A2(n[110]), .Z(t_110) );
  CKXOR2D1 C621 ( .A1(t_108), .A2(n[109]), .Z(t_109) );
  CKXOR2D1 C620 ( .A1(t_107), .A2(n[108]), .Z(t_108) );
  CKXOR2D1 C619 ( .A1(t_106), .A2(n[107]), .Z(t_107) );
  CKXOR2D1 C618 ( .A1(t_105), .A2(n[106]), .Z(t_106) );
  CKXOR2D1 C617 ( .A1(t_104), .A2(n[105]), .Z(t_105) );
  CKXOR2D1 C616 ( .A1(t_103), .A2(n[104]), .Z(t_104) );
  CKXOR2D1 C615 ( .A1(t_102), .A2(n[103]), .Z(t_103) );
  CKXOR2D1 C614 ( .A1(t_101), .A2(n[102]), .Z(t_102) );
  CKXOR2D1 C613 ( .A1(t_100), .A2(n[101]), .Z(t_101) );
  CKXOR2D1 C612 ( .A1(t_99), .A2(n[100]), .Z(t_100) );
  CKXOR2D1 C611 ( .A1(t_98), .A2(n[99]), .Z(t_99) );
  CKXOR2D1 C610 ( .A1(t_97), .A2(n[98]), .Z(t_98) );
  CKXOR2D1 C609 ( .A1(t_96), .A2(n[97]), .Z(t_97) );
  CKXOR2D1 C608 ( .A1(t_95), .A2(n[96]), .Z(t_96) );
  CKXOR2D1 C607 ( .A1(t_94), .A2(n[95]), .Z(t_95) );
  CKXOR2D1 C606 ( .A1(t_93), .A2(n[94]), .Z(t_94) );
  CKXOR2D1 C605 ( .A1(t_92), .A2(n[93]), .Z(t_93) );
  CKXOR2D1 C604 ( .A1(t_91), .A2(n[92]), .Z(t_92) );
  CKXOR2D1 C603 ( .A1(t_90), .A2(n[91]), .Z(t_91) );
  CKXOR2D1 C602 ( .A1(t_89), .A2(n[90]), .Z(t_90) );
  CKXOR2D1 C601 ( .A1(t_88), .A2(n[89]), .Z(t_89) );
  CKXOR2D1 C600 ( .A1(t_87), .A2(n[88]), .Z(t_88) );
  CKXOR2D1 C599 ( .A1(t_86), .A2(n[87]), .Z(t_87) );
  CKXOR2D1 C598 ( .A1(t_85), .A2(n[86]), .Z(t_86) );
  CKXOR2D1 C597 ( .A1(t_84), .A2(n[85]), .Z(t_85) );
  CKXOR2D1 C596 ( .A1(t_83), .A2(n[84]), .Z(t_84) );
  CKXOR2D1 C595 ( .A1(t_82), .A2(n[83]), .Z(t_83) );
  CKXOR2D1 C594 ( .A1(t_81), .A2(n[82]), .Z(t_82) );
  CKXOR2D1 C593 ( .A1(t_80), .A2(n[81]), .Z(t_81) );
  CKXOR2D1 C592 ( .A1(t_79), .A2(n[80]), .Z(t_80) );
  CKXOR2D1 C591 ( .A1(t_78), .A2(n[79]), .Z(t_79) );
  CKXOR2D1 C590 ( .A1(t_77), .A2(n[78]), .Z(t_78) );
  CKXOR2D1 C589 ( .A1(t_76), .A2(n[77]), .Z(t_77) );
  CKXOR2D1 C588 ( .A1(t_75), .A2(n[76]), .Z(t_76) );
  CKXOR2D1 C587 ( .A1(t_74), .A2(n[75]), .Z(t_75) );
  CKXOR2D1 C586 ( .A1(t_73), .A2(n[74]), .Z(t_74) );
  CKXOR2D1 C585 ( .A1(t_72), .A2(n[73]), .Z(t_73) );
  CKXOR2D1 C584 ( .A1(t_71), .A2(n[72]), .Z(t_72) );
  CKXOR2D1 C583 ( .A1(t_70), .A2(n[71]), .Z(t_71) );
  CKXOR2D1 C582 ( .A1(t_69), .A2(n[70]), .Z(t_70) );
  CKXOR2D1 C581 ( .A1(t_68), .A2(n[69]), .Z(t_69) );
  CKXOR2D1 C580 ( .A1(t_67), .A2(n[68]), .Z(t_68) );
  CKXOR2D1 C579 ( .A1(t_66), .A2(n[67]), .Z(t_67) );
  CKXOR2D1 C578 ( .A1(t_65), .A2(n[66]), .Z(t_66) );
  CKXOR2D1 C577 ( .A1(t_64), .A2(n[65]), .Z(t_65) );
  CKXOR2D1 C576 ( .A1(t_63), .A2(n[64]), .Z(t_64) );
  CKXOR2D1 C575 ( .A1(t_62), .A2(n[63]), .Z(t_63) );
  CKXOR2D1 C574 ( .A1(t_61), .A2(n[62]), .Z(t_62) );
  CKXOR2D1 C573 ( .A1(t_60), .A2(n[61]), .Z(t_61) );
  CKXOR2D1 C572 ( .A1(t_59), .A2(n[60]), .Z(t_60) );
  CKXOR2D1 C571 ( .A1(t_58), .A2(n[59]), .Z(t_59) );
  CKXOR2D1 C570 ( .A1(t_57), .A2(n[58]), .Z(t_58) );
  CKXOR2D1 C569 ( .A1(n[56]), .A2(n[57]), .Z(t_57) );
  CKXOR2D1 C568 ( .A1(a[4]), .A2(b[4]), .Z(N4) );
  CKXOR2D1 C567 ( .A1(N4), .A2(t_55), .Z(s[4]) );
  CKXOR2D1 C566 ( .A1(t_54), .A2(n[55]), .Z(t_55) );
  CKXOR2D1 C565 ( .A1(t_53), .A2(n[54]), .Z(t_54) );
  CKXOR2D1 C564 ( .A1(t_52), .A2(n[53]), .Z(t_53) );
  CKXOR2D1 C563 ( .A1(t_51), .A2(n[52]), .Z(t_52) );
  CKXOR2D1 C562 ( .A1(t_50), .A2(n[51]), .Z(t_51) );
  CKXOR2D1 C561 ( .A1(t_49), .A2(n[50]), .Z(t_50) );
  CKXOR2D1 C560 ( .A1(t_48), .A2(n[49]), .Z(t_49) );
  CKXOR2D1 C559 ( .A1(t_47), .A2(n[48]), .Z(t_48) );
  CKXOR2D1 C558 ( .A1(t_46), .A2(n[47]), .Z(t_47) );
  CKXOR2D1 C557 ( .A1(t_45), .A2(n[46]), .Z(t_46) );
  CKXOR2D1 C556 ( .A1(t_44), .A2(n[45]), .Z(t_45) );
  CKXOR2D1 C555 ( .A1(t_43), .A2(n[44]), .Z(t_44) );
  CKXOR2D1 C554 ( .A1(t_42), .A2(n[43]), .Z(t_43) );
  CKXOR2D1 C553 ( .A1(t_41), .A2(n[42]), .Z(t_42) );
  CKXOR2D1 C552 ( .A1(t_40), .A2(n[41]), .Z(t_41) );
  CKXOR2D1 C551 ( .A1(t_39), .A2(n[40]), .Z(t_40) );
  CKXOR2D1 C550 ( .A1(t_38), .A2(n[39]), .Z(t_39) );
  CKXOR2D1 C549 ( .A1(t_37), .A2(n[38]), .Z(t_38) );
  CKXOR2D1 C548 ( .A1(t_36), .A2(n[37]), .Z(t_37) );
  CKXOR2D1 C547 ( .A1(t_35), .A2(n[36]), .Z(t_36) );
  CKXOR2D1 C546 ( .A1(t_34), .A2(n[35]), .Z(t_35) );
  CKXOR2D1 C545 ( .A1(t_33), .A2(n[34]), .Z(t_34) );
  CKXOR2D1 C544 ( .A1(t_32), .A2(n[33]), .Z(t_33) );
  CKXOR2D1 C543 ( .A1(t_31), .A2(n[32]), .Z(t_32) );
  CKXOR2D1 C542 ( .A1(t_30), .A2(n[31]), .Z(t_31) );
  CKXOR2D1 C541 ( .A1(t_29), .A2(n[30]), .Z(t_30) );
  CKXOR2D1 C540 ( .A1(t_28), .A2(n[29]), .Z(t_29) );
  CKXOR2D1 C539 ( .A1(t_27), .A2(n[28]), .Z(t_28) );
  CKXOR2D1 C538 ( .A1(t_26), .A2(n[27]), .Z(t_27) );
  CKXOR2D1 C537 ( .A1(n[25]), .A2(n[26]), .Z(t_26) );
  CKXOR2D1 C536 ( .A1(a[3]), .A2(b[3]), .Z(N3) );
  CKXOR2D1 C535 ( .A1(N3), .A2(t_24), .Z(s[3]) );
  CKXOR2D1 C534 ( .A1(t_23), .A2(n[24]), .Z(t_24) );
  CKXOR2D1 C533 ( .A1(t_22), .A2(n[23]), .Z(t_23) );
  CKXOR2D1 C532 ( .A1(t_21), .A2(n[22]), .Z(t_22) );
  CKXOR2D1 C531 ( .A1(t_20), .A2(n[21]), .Z(t_21) );
  CKXOR2D1 C530 ( .A1(t_19), .A2(n[20]), .Z(t_20) );
  CKXOR2D1 C529 ( .A1(t_18), .A2(n[19]), .Z(t_19) );
  CKXOR2D1 C528 ( .A1(t_17), .A2(n[18]), .Z(t_18) );
  CKXOR2D1 C527 ( .A1(t_16), .A2(n[17]), .Z(t_17) );
  CKXOR2D1 C526 ( .A1(t_15), .A2(n[16]), .Z(t_16) );
  CKXOR2D1 C525 ( .A1(t_14), .A2(n[15]), .Z(t_15) );
  CKXOR2D1 C524 ( .A1(t_13), .A2(n[14]), .Z(t_14) );
  CKXOR2D1 C523 ( .A1(t_12), .A2(n[13]), .Z(t_13) );
  CKXOR2D1 C522 ( .A1(t_11), .A2(n[12]), .Z(t_12) );
  CKXOR2D1 C521 ( .A1(n[10]), .A2(n[11]), .Z(t_11) );
  CKXOR2D1 C520 ( .A1(a[2]), .A2(b[2]), .Z(N2) );
  CKXOR2D1 C519 ( .A1(N2), .A2(t_9), .Z(s[2]) );
  CKXOR2D1 C518 ( .A1(t_8), .A2(n[9]), .Z(t_9) );
  CKXOR2D1 C517 ( .A1(t_7), .A2(n[8]), .Z(t_8) );
  CKXOR2D1 C516 ( .A1(t_6), .A2(n[7]), .Z(t_7) );
  CKXOR2D1 C515 ( .A1(t_5), .A2(n[6]), .Z(t_6) );
  CKXOR2D1 C514 ( .A1(t_4), .A2(n[5]), .Z(t_5) );
  CKXOR2D1 C513 ( .A1(n[3]), .A2(n[4]), .Z(t_4) );
  CKXOR2D1 C512 ( .A1(a[1]), .A2(b[1]), .Z(N1) );
  CKXOR2D1 C511 ( .A1(N1), .A2(t_2), .Z(s[1]) );
  CKXOR2D1 C510 ( .A1(t_1), .A2(n[2]), .Z(t_2) );
  CKXOR2D1 C509 ( .A1(n[0]), .A2(n[1]), .Z(t_1) );
  CKXOR2D1 C508 ( .A1(a[0]), .A2(b[0]), .Z(N0) );
  CKXOR2D1 C507 ( .A1(N0), .A2(c_in), .Z(s[0]) );
endmodule

