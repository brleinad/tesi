
module linear ( a, b, n, code );
  input [6:0] a;
  input [6:0] b;
  input [500:0] n;
  output [14:0] code;
  wire   N2, t_118, t_117, t_116, t_115, t_114, t_113, t_112, t_111, t_110,
         t_109, t_108, t_107, t_106, t_105, t_104, t_103, t_102, t_101, t_100,
         t_99, t_98, t_97, t_96, t_95, t_94, t_93, t_92, t_91, t_90, t_89,
         t_88, t_87, t_86, t_85, t_84, t_83, t_82, t_81, t_80, t_79, t_78,
         t_77, t_76, t_75, t_74, t_73, t_72, t_71, t_70, t_69, t_68, t_67,
         t_66, t_65, t_64, t_63, t_62, t_61, t_60, t_59, t_58, t_57, t_55,
         t_54, t_53, t_52, t_51, t_50, t_49, t_48, t_47, t_46, t_45, t_44,
         t_43, t_42, t_41, t_40, t_39, t_38, t_37, t_36, t_35, t_34, t_33,
         t_32, t_31, t_30, t_29, t_28, t_27, t_26, t_24, t_23, t_22, t_21,
         t_20, t_19, t_18, t_17, t_16, t_15, t_14, t_13, t_12, t_11, t_9, t_8,
         t_7, t_6, t_5, t_4, t_2, t_1, N14, N15, N16, N17, N18, N19, n1, n2,
         n3, n4, n5, n6, n7;
  wire   [245:120] t;

  CKXOR2D1HVT C759 ( .A1(a[6]), .A2(b[6]), .Z(N19) );
  CKXOR2D1HVT C758 ( .A1(N19), .A2(t[245]), .Z(code[6]) );
  CKXOR2D1HVT C757 ( .A1(t[244]), .A2(n[245]), .Z(t[245]) );
  CKXOR2D1HVT C756 ( .A1(t[243]), .A2(n[244]), .Z(t[244]) );
  CKXOR2D1HVT C755 ( .A1(t[242]), .A2(n[243]), .Z(t[243]) );
  CKXOR2D1HVT C754 ( .A1(t[241]), .A2(n[242]), .Z(t[242]) );
  CKXOR2D1HVT C753 ( .A1(t[240]), .A2(n[241]), .Z(t[241]) );
  CKXOR2D1HVT C752 ( .A1(t[239]), .A2(n[240]), .Z(t[240]) );
  CKXOR2D1HVT C751 ( .A1(t[238]), .A2(n[239]), .Z(t[239]) );
  CKXOR2D1HVT C750 ( .A1(t[237]), .A2(n[238]), .Z(t[238]) );
  CKXOR2D1HVT C749 ( .A1(t[236]), .A2(n[237]), .Z(t[237]) );
  CKXOR2D1HVT C748 ( .A1(t[235]), .A2(n[236]), .Z(t[236]) );
  CKXOR2D1HVT C747 ( .A1(t[234]), .A2(n[235]), .Z(t[235]) );
  CKXOR2D1HVT C746 ( .A1(t[233]), .A2(n[234]), .Z(t[234]) );
  CKXOR2D1HVT C745 ( .A1(t[232]), .A2(n[233]), .Z(t[233]) );
  CKXOR2D1HVT C744 ( .A1(t[231]), .A2(n[232]), .Z(t[232]) );
  CKXOR2D1HVT C743 ( .A1(t[230]), .A2(n[231]), .Z(t[231]) );
  CKXOR2D1HVT C742 ( .A1(t[229]), .A2(n[230]), .Z(t[230]) );
  CKXOR2D1HVT C741 ( .A1(t[228]), .A2(n[229]), .Z(t[229]) );
  CKXOR2D1HVT C740 ( .A1(t[227]), .A2(n[228]), .Z(t[228]) );
  CKXOR2D1HVT C739 ( .A1(t[226]), .A2(n[227]), .Z(t[227]) );
  CKXOR2D1HVT C738 ( .A1(t[225]), .A2(n[226]), .Z(t[226]) );
  CKXOR2D1HVT C737 ( .A1(t[224]), .A2(n[225]), .Z(t[225]) );
  CKXOR2D1HVT C736 ( .A1(t[223]), .A2(n[224]), .Z(t[224]) );
  CKXOR2D1HVT C735 ( .A1(t[222]), .A2(n[223]), .Z(t[223]) );
  CKXOR2D1HVT C734 ( .A1(t[221]), .A2(n[222]), .Z(t[222]) );
  CKXOR2D1HVT C733 ( .A1(t[220]), .A2(n[221]), .Z(t[221]) );
  CKXOR2D1HVT C732 ( .A1(t[219]), .A2(n[220]), .Z(t[220]) );
  CKXOR2D1HVT C731 ( .A1(t[218]), .A2(n[219]), .Z(t[219]) );
  CKXOR2D1HVT C730 ( .A1(t[217]), .A2(n[218]), .Z(t[218]) );
  CKXOR2D1HVT C729 ( .A1(t[216]), .A2(n[217]), .Z(t[217]) );
  CKXOR2D1HVT C728 ( .A1(t[215]), .A2(n[216]), .Z(t[216]) );
  CKXOR2D1HVT C727 ( .A1(t[214]), .A2(n[215]), .Z(t[215]) );
  CKXOR2D1HVT C726 ( .A1(t[213]), .A2(n[214]), .Z(t[214]) );
  CKXOR2D1HVT C725 ( .A1(t[212]), .A2(n[213]), .Z(t[213]) );
  CKXOR2D1HVT C724 ( .A1(t[211]), .A2(n[212]), .Z(t[212]) );
  CKXOR2D1HVT C723 ( .A1(t[210]), .A2(n[211]), .Z(t[211]) );
  CKXOR2D1HVT C722 ( .A1(t[209]), .A2(n[210]), .Z(t[210]) );
  CKXOR2D1HVT C721 ( .A1(t[208]), .A2(n[209]), .Z(t[209]) );
  CKXOR2D1HVT C720 ( .A1(t[207]), .A2(n[208]), .Z(t[208]) );
  CKXOR2D1HVT C719 ( .A1(t[206]), .A2(n[207]), .Z(t[207]) );
  CKXOR2D1HVT C718 ( .A1(t[205]), .A2(n[206]), .Z(t[206]) );
  CKXOR2D1HVT C717 ( .A1(t[204]), .A2(n[205]), .Z(t[205]) );
  CKXOR2D1HVT C716 ( .A1(t[203]), .A2(n[204]), .Z(t[204]) );
  CKXOR2D1HVT C715 ( .A1(t[202]), .A2(n[203]), .Z(t[203]) );
  CKXOR2D1HVT C714 ( .A1(t[201]), .A2(n[202]), .Z(t[202]) );
  CKXOR2D1HVT C713 ( .A1(t[200]), .A2(n[201]), .Z(t[201]) );
  CKXOR2D1HVT C712 ( .A1(t[199]), .A2(n[200]), .Z(t[200]) );
  CKXOR2D1HVT C711 ( .A1(t[198]), .A2(n[199]), .Z(t[199]) );
  CKXOR2D1HVT C710 ( .A1(t[197]), .A2(n[198]), .Z(t[198]) );
  CKXOR2D1HVT C709 ( .A1(t[196]), .A2(n[197]), .Z(t[197]) );
  CKXOR2D1HVT C708 ( .A1(t[195]), .A2(n[196]), .Z(t[196]) );
  CKXOR2D1HVT C707 ( .A1(t[194]), .A2(n[195]), .Z(t[195]) );
  CKXOR2D1HVT C706 ( .A1(t[193]), .A2(n[194]), .Z(t[194]) );
  CKXOR2D1HVT C705 ( .A1(t[192]), .A2(n[193]), .Z(t[193]) );
  CKXOR2D1HVT C704 ( .A1(t[191]), .A2(n[192]), .Z(t[192]) );
  CKXOR2D1HVT C703 ( .A1(t[190]), .A2(n[191]), .Z(t[191]) );
  CKXOR2D1HVT C702 ( .A1(t[189]), .A2(n[190]), .Z(t[190]) );
  CKXOR2D1HVT C701 ( .A1(t[188]), .A2(n[189]), .Z(t[189]) );
  CKXOR2D1HVT C700 ( .A1(t[187]), .A2(n[188]), .Z(t[188]) );
  CKXOR2D1HVT C699 ( .A1(t[186]), .A2(n[187]), .Z(t[187]) );
  CKXOR2D1HVT C698 ( .A1(t[185]), .A2(n[186]), .Z(t[186]) );
  CKXOR2D1HVT C697 ( .A1(t[184]), .A2(n[185]), .Z(t[185]) );
  CKXOR2D1HVT C696 ( .A1(t[183]), .A2(n[184]), .Z(t[184]) );
  CKXOR2D1HVT C695 ( .A1(t[182]), .A2(n[183]), .Z(t[183]) );
  CKXOR2D1HVT C694 ( .A1(t[181]), .A2(n[182]), .Z(t[182]) );
  CKXOR2D1HVT C693 ( .A1(t[180]), .A2(n[181]), .Z(t[181]) );
  CKXOR2D1HVT C692 ( .A1(t[179]), .A2(n[180]), .Z(t[180]) );
  CKXOR2D1HVT C691 ( .A1(t[178]), .A2(n[179]), .Z(t[179]) );
  CKXOR2D1HVT C690 ( .A1(t[177]), .A2(n[178]), .Z(t[178]) );
  CKXOR2D1HVT C689 ( .A1(t[176]), .A2(n[177]), .Z(t[177]) );
  CKXOR2D1HVT C688 ( .A1(t[175]), .A2(n[176]), .Z(t[176]) );
  CKXOR2D1HVT C687 ( .A1(t[174]), .A2(n[175]), .Z(t[175]) );
  CKXOR2D1HVT C686 ( .A1(t[173]), .A2(n[174]), .Z(t[174]) );
  CKXOR2D1HVT C685 ( .A1(t[172]), .A2(n[173]), .Z(t[173]) );
  CKXOR2D1HVT C684 ( .A1(t[171]), .A2(n[172]), .Z(t[172]) );
  CKXOR2D1HVT C683 ( .A1(t[170]), .A2(n[171]), .Z(t[171]) );
  CKXOR2D1HVT C682 ( .A1(t[169]), .A2(n[170]), .Z(t[170]) );
  CKXOR2D1HVT C681 ( .A1(t[168]), .A2(n[169]), .Z(t[169]) );
  CKXOR2D1HVT C680 ( .A1(t[167]), .A2(n[168]), .Z(t[168]) );
  CKXOR2D1HVT C679 ( .A1(t[166]), .A2(n[167]), .Z(t[167]) );
  CKXOR2D1HVT C678 ( .A1(t[165]), .A2(n[166]), .Z(t[166]) );
  CKXOR2D1HVT C677 ( .A1(t[164]), .A2(n[165]), .Z(t[165]) );
  CKXOR2D1HVT C676 ( .A1(t[163]), .A2(n[164]), .Z(t[164]) );
  CKXOR2D1HVT C675 ( .A1(t[162]), .A2(n[163]), .Z(t[163]) );
  CKXOR2D1HVT C674 ( .A1(t[161]), .A2(n[162]), .Z(t[162]) );
  CKXOR2D1HVT C673 ( .A1(t[160]), .A2(n[161]), .Z(t[161]) );
  CKXOR2D1HVT C672 ( .A1(t[159]), .A2(n[160]), .Z(t[160]) );
  CKXOR2D1HVT C671 ( .A1(t[158]), .A2(n[159]), .Z(t[159]) );
  CKXOR2D1HVT C670 ( .A1(t[157]), .A2(n[158]), .Z(t[158]) );
  CKXOR2D1HVT C669 ( .A1(t[156]), .A2(n[157]), .Z(t[157]) );
  CKXOR2D1HVT C668 ( .A1(t[155]), .A2(n[156]), .Z(t[156]) );
  CKXOR2D1HVT C667 ( .A1(t[154]), .A2(n[155]), .Z(t[155]) );
  CKXOR2D1HVT C666 ( .A1(t[153]), .A2(n[154]), .Z(t[154]) );
  CKXOR2D1HVT C665 ( .A1(t[152]), .A2(n[153]), .Z(t[153]) );
  CKXOR2D1HVT C664 ( .A1(t[151]), .A2(n[152]), .Z(t[152]) );
  CKXOR2D1HVT C663 ( .A1(t[150]), .A2(n[151]), .Z(t[151]) );
  CKXOR2D1HVT C662 ( .A1(t[149]), .A2(n[150]), .Z(t[150]) );
  CKXOR2D1HVT C661 ( .A1(t[148]), .A2(n[149]), .Z(t[149]) );
  CKXOR2D1HVT C660 ( .A1(t[147]), .A2(n[148]), .Z(t[148]) );
  CKXOR2D1HVT C659 ( .A1(t[146]), .A2(n[147]), .Z(t[147]) );
  CKXOR2D1HVT C658 ( .A1(t[145]), .A2(n[146]), .Z(t[146]) );
  CKXOR2D1HVT C657 ( .A1(t[144]), .A2(n[145]), .Z(t[145]) );
  CKXOR2D1HVT C656 ( .A1(t[143]), .A2(n[144]), .Z(t[144]) );
  CKXOR2D1HVT C655 ( .A1(t[142]), .A2(n[143]), .Z(t[143]) );
  CKXOR2D1HVT C654 ( .A1(t[141]), .A2(n[142]), .Z(t[142]) );
  CKXOR2D1HVT C653 ( .A1(t[140]), .A2(n[141]), .Z(t[141]) );
  CKXOR2D1HVT C652 ( .A1(t[139]), .A2(n[140]), .Z(t[140]) );
  CKXOR2D1HVT C651 ( .A1(t[138]), .A2(n[139]), .Z(t[139]) );
  CKXOR2D1HVT C650 ( .A1(t[137]), .A2(n[138]), .Z(t[138]) );
  CKXOR2D1HVT C649 ( .A1(t[136]), .A2(n[137]), .Z(t[137]) );
  CKXOR2D1HVT C648 ( .A1(t[135]), .A2(n[136]), .Z(t[136]) );
  CKXOR2D1HVT C647 ( .A1(t[134]), .A2(n[135]), .Z(t[135]) );
  CKXOR2D1HVT C646 ( .A1(t[133]), .A2(n[134]), .Z(t[134]) );
  CKXOR2D1HVT C645 ( .A1(t[132]), .A2(n[133]), .Z(t[133]) );
  CKXOR2D1HVT C644 ( .A1(t[131]), .A2(n[132]), .Z(t[132]) );
  CKXOR2D1HVT C643 ( .A1(t[130]), .A2(n[131]), .Z(t[131]) );
  CKXOR2D1HVT C642 ( .A1(t[129]), .A2(n[130]), .Z(t[130]) );
  CKXOR2D1HVT C641 ( .A1(t[128]), .A2(n[129]), .Z(t[129]) );
  CKXOR2D1HVT C640 ( .A1(t[127]), .A2(n[128]), .Z(t[128]) );
  CKXOR2D1HVT C639 ( .A1(t[126]), .A2(n[127]), .Z(t[127]) );
  CKXOR2D1HVT C638 ( .A1(t[125]), .A2(n[126]), .Z(t[126]) );
  CKXOR2D1HVT C637 ( .A1(t[124]), .A2(n[125]), .Z(t[125]) );
  CKXOR2D1HVT C636 ( .A1(t[123]), .A2(n[124]), .Z(t[124]) );
  CKXOR2D1HVT C635 ( .A1(t[122]), .A2(n[123]), .Z(t[123]) );
  CKXOR2D1HVT C634 ( .A1(t[121]), .A2(n[122]), .Z(t[122]) );
  CKXOR2D1HVT C633 ( .A1(t[120]), .A2(n[121]), .Z(t[121]) );
  CKXOR2D1HVT C632 ( .A1(n[119]), .A2(n[120]), .Z(t[120]) );
  CKXOR2D1HVT C631 ( .A1(a[5]), .A2(b[5]), .Z(N18) );
  CKXOR2D1HVT C630 ( .A1(N18), .A2(t_118), .Z(code[5]) );
  CKXOR2D1HVT C629 ( .A1(t_117), .A2(n[118]), .Z(t_118) );
  CKXOR2D1HVT C628 ( .A1(t_116), .A2(n[117]), .Z(t_117) );
  CKXOR2D1HVT C627 ( .A1(t_115), .A2(n[116]), .Z(t_116) );
  CKXOR2D1HVT C626 ( .A1(t_114), .A2(n[115]), .Z(t_115) );
  CKXOR2D1HVT C625 ( .A1(t_113), .A2(n[114]), .Z(t_114) );
  CKXOR2D1HVT C624 ( .A1(t_112), .A2(n[113]), .Z(t_113) );
  CKXOR2D1HVT C623 ( .A1(t_111), .A2(n[112]), .Z(t_112) );
  CKXOR2D1HVT C622 ( .A1(t_110), .A2(n[111]), .Z(t_111) );
  CKXOR2D1HVT C621 ( .A1(t_109), .A2(n[110]), .Z(t_110) );
  CKXOR2D1HVT C620 ( .A1(t_108), .A2(n[109]), .Z(t_109) );
  CKXOR2D1HVT C619 ( .A1(t_107), .A2(n[108]), .Z(t_108) );
  CKXOR2D1HVT C618 ( .A1(t_106), .A2(n[107]), .Z(t_107) );
  CKXOR2D1HVT C617 ( .A1(t_105), .A2(n[106]), .Z(t_106) );
  CKXOR2D1HVT C616 ( .A1(t_104), .A2(n[105]), .Z(t_105) );
  CKXOR2D1HVT C615 ( .A1(t_103), .A2(n[104]), .Z(t_104) );
  CKXOR2D1HVT C614 ( .A1(t_102), .A2(n[103]), .Z(t_103) );
  CKXOR2D1HVT C613 ( .A1(t_101), .A2(n[102]), .Z(t_102) );
  CKXOR2D1HVT C612 ( .A1(t_100), .A2(n[101]), .Z(t_101) );
  CKXOR2D1HVT C611 ( .A1(t_99), .A2(n[100]), .Z(t_100) );
  CKXOR2D1HVT C610 ( .A1(t_98), .A2(n[99]), .Z(t_99) );
  CKXOR2D1HVT C609 ( .A1(t_97), .A2(n[98]), .Z(t_98) );
  CKXOR2D1HVT C608 ( .A1(t_96), .A2(n[97]), .Z(t_97) );
  CKXOR2D1HVT C607 ( .A1(t_95), .A2(n[96]), .Z(t_96) );
  CKXOR2D1HVT C606 ( .A1(t_94), .A2(n[95]), .Z(t_95) );
  CKXOR2D1HVT C605 ( .A1(t_93), .A2(n[94]), .Z(t_94) );
  CKXOR2D1HVT C604 ( .A1(t_92), .A2(n[93]), .Z(t_93) );
  CKXOR2D1HVT C603 ( .A1(t_91), .A2(n[92]), .Z(t_92) );
  CKXOR2D1HVT C602 ( .A1(t_90), .A2(n[91]), .Z(t_91) );
  CKXOR2D1HVT C601 ( .A1(t_89), .A2(n[90]), .Z(t_90) );
  CKXOR2D1HVT C600 ( .A1(t_88), .A2(n[89]), .Z(t_89) );
  CKXOR2D1HVT C599 ( .A1(t_87), .A2(n[88]), .Z(t_88) );
  CKXOR2D1HVT C598 ( .A1(t_86), .A2(n[87]), .Z(t_87) );
  CKXOR2D1HVT C597 ( .A1(t_85), .A2(n[86]), .Z(t_86) );
  CKXOR2D1HVT C596 ( .A1(t_84), .A2(n[85]), .Z(t_85) );
  CKXOR2D1HVT C595 ( .A1(t_83), .A2(n[84]), .Z(t_84) );
  CKXOR2D1HVT C594 ( .A1(t_82), .A2(n[83]), .Z(t_83) );
  CKXOR2D1HVT C593 ( .A1(t_81), .A2(n[82]), .Z(t_82) );
  CKXOR2D1HVT C592 ( .A1(t_80), .A2(n[81]), .Z(t_81) );
  CKXOR2D1HVT C591 ( .A1(t_79), .A2(n[80]), .Z(t_80) );
  CKXOR2D1HVT C590 ( .A1(t_78), .A2(n[79]), .Z(t_79) );
  CKXOR2D1HVT C589 ( .A1(t_77), .A2(n[78]), .Z(t_78) );
  CKXOR2D1HVT C588 ( .A1(t_76), .A2(n[77]), .Z(t_77) );
  CKXOR2D1HVT C587 ( .A1(t_75), .A2(n[76]), .Z(t_76) );
  CKXOR2D1HVT C586 ( .A1(t_74), .A2(n[75]), .Z(t_75) );
  CKXOR2D1HVT C585 ( .A1(t_73), .A2(n[74]), .Z(t_74) );
  CKXOR2D1HVT C584 ( .A1(t_72), .A2(n[73]), .Z(t_73) );
  CKXOR2D1HVT C583 ( .A1(t_71), .A2(n[72]), .Z(t_72) );
  CKXOR2D1HVT C582 ( .A1(t_70), .A2(n[71]), .Z(t_71) );
  CKXOR2D1HVT C581 ( .A1(t_69), .A2(n[70]), .Z(t_70) );
  CKXOR2D1HVT C580 ( .A1(t_68), .A2(n[69]), .Z(t_69) );
  CKXOR2D1HVT C579 ( .A1(t_67), .A2(n[68]), .Z(t_68) );
  CKXOR2D1HVT C578 ( .A1(t_66), .A2(n[67]), .Z(t_67) );
  CKXOR2D1HVT C577 ( .A1(t_65), .A2(n[66]), .Z(t_66) );
  CKXOR2D1HVT C576 ( .A1(t_64), .A2(n[65]), .Z(t_65) );
  CKXOR2D1HVT C575 ( .A1(t_63), .A2(n[64]), .Z(t_64) );
  CKXOR2D1HVT C574 ( .A1(t_62), .A2(n[63]), .Z(t_63) );
  CKXOR2D1HVT C573 ( .A1(t_61), .A2(n[62]), .Z(t_62) );
  CKXOR2D1HVT C572 ( .A1(t_60), .A2(n[61]), .Z(t_61) );
  CKXOR2D1HVT C571 ( .A1(t_59), .A2(n[60]), .Z(t_60) );
  CKXOR2D1HVT C570 ( .A1(t_58), .A2(n[59]), .Z(t_59) );
  CKXOR2D1HVT C569 ( .A1(t_57), .A2(n[58]), .Z(t_58) );
  CKXOR2D1HVT C568 ( .A1(n[56]), .A2(n[57]), .Z(t_57) );
  CKXOR2D1HVT C567 ( .A1(a[4]), .A2(b[4]), .Z(N17) );
  CKXOR2D1HVT C566 ( .A1(N17), .A2(t_55), .Z(code[4]) );
  CKXOR2D1HVT C565 ( .A1(t_54), .A2(n[55]), .Z(t_55) );
  CKXOR2D1HVT C564 ( .A1(t_53), .A2(n[54]), .Z(t_54) );
  CKXOR2D1HVT C563 ( .A1(t_52), .A2(n[53]), .Z(t_53) );
  CKXOR2D1HVT C562 ( .A1(t_51), .A2(n[52]), .Z(t_52) );
  CKXOR2D1HVT C561 ( .A1(t_50), .A2(n[51]), .Z(t_51) );
  CKXOR2D1HVT C560 ( .A1(t_49), .A2(n[50]), .Z(t_50) );
  CKXOR2D1HVT C559 ( .A1(t_48), .A2(n[49]), .Z(t_49) );
  CKXOR2D1HVT C558 ( .A1(t_47), .A2(n[48]), .Z(t_48) );
  CKXOR2D1HVT C557 ( .A1(t_46), .A2(n[47]), .Z(t_47) );
  CKXOR2D1HVT C556 ( .A1(t_45), .A2(n[46]), .Z(t_46) );
  CKXOR2D1HVT C555 ( .A1(t_44), .A2(n[45]), .Z(t_45) );
  CKXOR2D1HVT C554 ( .A1(t_43), .A2(n[44]), .Z(t_44) );
  CKXOR2D1HVT C553 ( .A1(t_42), .A2(n[43]), .Z(t_43) );
  CKXOR2D1HVT C552 ( .A1(t_41), .A2(n[42]), .Z(t_42) );
  CKXOR2D1HVT C551 ( .A1(t_40), .A2(n[41]), .Z(t_41) );
  CKXOR2D1HVT C550 ( .A1(t_39), .A2(n[40]), .Z(t_40) );
  CKXOR2D1HVT C549 ( .A1(t_38), .A2(n[39]), .Z(t_39) );
  CKXOR2D1HVT C548 ( .A1(t_37), .A2(n[38]), .Z(t_38) );
  CKXOR2D1HVT C547 ( .A1(t_36), .A2(n[37]), .Z(t_37) );
  CKXOR2D1HVT C546 ( .A1(t_35), .A2(n[36]), .Z(t_36) );
  CKXOR2D1HVT C545 ( .A1(t_34), .A2(n[35]), .Z(t_35) );
  CKXOR2D1HVT C544 ( .A1(t_33), .A2(n[34]), .Z(t_34) );
  CKXOR2D1HVT C543 ( .A1(t_32), .A2(n[33]), .Z(t_33) );
  CKXOR2D1HVT C542 ( .A1(t_31), .A2(n[32]), .Z(t_32) );
  CKXOR2D1HVT C541 ( .A1(t_30), .A2(n[31]), .Z(t_31) );
  CKXOR2D1HVT C540 ( .A1(t_29), .A2(n[30]), .Z(t_30) );
  CKXOR2D1HVT C539 ( .A1(t_28), .A2(n[29]), .Z(t_29) );
  CKXOR2D1HVT C538 ( .A1(t_27), .A2(n[28]), .Z(t_28) );
  CKXOR2D1HVT C537 ( .A1(t_26), .A2(n[27]), .Z(t_27) );
  CKXOR2D1HVT C536 ( .A1(n[25]), .A2(n[26]), .Z(t_26) );
  CKXOR2D1HVT C535 ( .A1(a[3]), .A2(b[3]), .Z(N16) );
  CKXOR2D1HVT C534 ( .A1(N16), .A2(t_24), .Z(code[3]) );
  CKXOR2D1HVT C533 ( .A1(t_23), .A2(n[24]), .Z(t_24) );
  CKXOR2D1HVT C532 ( .A1(t_22), .A2(n[23]), .Z(t_23) );
  CKXOR2D1HVT C531 ( .A1(t_21), .A2(n[22]), .Z(t_22) );
  CKXOR2D1HVT C530 ( .A1(t_20), .A2(n[21]), .Z(t_21) );
  CKXOR2D1HVT C529 ( .A1(t_19), .A2(n[20]), .Z(t_20) );
  CKXOR2D1HVT C528 ( .A1(t_18), .A2(n[19]), .Z(t_19) );
  CKXOR2D1HVT C527 ( .A1(t_17), .A2(n[18]), .Z(t_18) );
  CKXOR2D1HVT C526 ( .A1(t_16), .A2(n[17]), .Z(t_17) );
  CKXOR2D1HVT C525 ( .A1(t_15), .A2(n[16]), .Z(t_16) );
  CKXOR2D1HVT C524 ( .A1(t_14), .A2(n[15]), .Z(t_15) );
  CKXOR2D1HVT C523 ( .A1(t_13), .A2(n[14]), .Z(t_14) );
  CKXOR2D1HVT C522 ( .A1(t_12), .A2(n[13]), .Z(t_13) );
  CKXOR2D1HVT C521 ( .A1(t_11), .A2(n[12]), .Z(t_12) );
  CKXOR2D1HVT C520 ( .A1(n[10]), .A2(n[11]), .Z(t_11) );
  CKXOR2D1HVT C519 ( .A1(a[2]), .A2(b[2]), .Z(N15) );
  CKXOR2D1HVT C518 ( .A1(N15), .A2(t_9), .Z(code[2]) );
  CKXOR2D1HVT C517 ( .A1(t_8), .A2(n[9]), .Z(t_9) );
  CKXOR2D1HVT C516 ( .A1(t_7), .A2(n[8]), .Z(t_8) );
  CKXOR2D1HVT C515 ( .A1(t_6), .A2(n[7]), .Z(t_7) );
  CKXOR2D1HVT C514 ( .A1(t_5), .A2(n[6]), .Z(t_6) );
  CKXOR2D1HVT C513 ( .A1(t_4), .A2(n[5]), .Z(t_5) );
  CKXOR2D1HVT C512 ( .A1(n[3]), .A2(n[4]), .Z(t_4) );
  CKXOR2D1HVT C511 ( .A1(a[1]), .A2(b[1]), .Z(N14) );
  CKXOR2D1HVT C510 ( .A1(N14), .A2(t_2), .Z(code[1]) );
  CKXOR2D1HVT C509 ( .A1(t_1), .A2(n[2]), .Z(t_2) );
  CKXOR2D1HVT C508 ( .A1(n[0]), .A2(n[1]), .Z(t_1) );
  CKXOR2D1HVT C507 ( .A1(a[0]), .A2(b[0]), .Z(code[0]) );
  CKXOR2D1HVT __tmp122_2 ( .A1(N2), .A2(code[5]), .Z(code[9]) );
  CKXOR2D1HVT __tmp122_1 ( .A1(code[2]), .A2(code[3]), .Z(N2) );
  CKXOR2D1HVT U1 ( .A1(code[3]), .A2(code[4]), .Z(n4) );
  CKXOR2D1HVT U2 ( .A1(code[6]), .A2(n4), .Z(code[10]) );
  CKXOR2D1HVT U3 ( .A1(code[1]), .A2(code[4]), .Z(n3) );
  CKXOR2D1HVT U4 ( .A1(code[2]), .A2(n3), .Z(code[8]) );
  CKXOR2D1HVT U5 ( .A1(code[0]), .A2(code[1]), .Z(n2) );
  CKXOR2D1HVT U6 ( .A1(n7), .A2(n4), .Z(code[11]) );
  CKXOR2D1HVT U7 ( .A1(code[5]), .A2(n2), .Z(n7) );
  CKXOR2D1HVT U8 ( .A1(code[3]), .A2(n2), .Z(code[7]) );
  CKXOR2D1HVT U9 ( .A1(code[2]), .A2(code[6]), .Z(n1) );
  CKXOR2D1HVT U10 ( .A1(code[0]), .A2(n1), .Z(code[14]) );
  CKXOR2D1HVT U11 ( .A1(n6), .A2(n2), .Z(code[13]) );
  CKXOR2D1HVT U12 ( .A1(code[5]), .A2(n1), .Z(n6) );
  CKXOR2D1HVT U13 ( .A1(n5), .A2(n3), .Z(code[12]) );
  CKXOR2D1HVT U14 ( .A1(code[5]), .A2(n1), .Z(n5) );
endmodule

