module Encoder_Logic(
in  [13:0] iv_data;
out [13:0] ov_data;
) ;										
	assign ov_data(0) = 	assign ov_data(1) = 	assign ov_data(2) = 	assign ov_data(3) = 	assign ov_data(4) = 	assign ov_data(5) = 	assign ov_data(6) = 	assign ov_data(7) = 	assign ov_data(8) = 	assign ov_data(9) = 	assign ov_data(10) = 	assign ov_data(11) = 	assign ov_data(12) = 	assign ov_data(13) = endmodule;
